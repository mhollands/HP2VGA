-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 14 2018 01:24:42

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    TVP_VIDEO : in std_logic_vector(9 downto 0);
    ADV_B : out std_logic_vector(7 downto 0);
    ADV_G : out std_logic_vector(7 downto 0);
    ADV_R : out std_logic_vector(7 downto 0);
    DEBUG : inout std_logic_vector(7 downto 0);
    TVP_CLK : in std_logic;
    ADV_CLK : out std_logic;
    TVP_HSYNC : in std_logic;
    ADV_HSYNC : out std_logic;
    TVP_VSYNC : in std_logic;
    ADV_VSYNC : out std_logic;
    ADV_BLANK_N : out std_logic;
    LED : out std_logic;
    ADV_SYNC_N : out std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__18943\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \VCCG0\ : std_logic;
signal \TVP_VIDEO_c_4\ : std_logic;
signal \GNDG0\ : std_logic;
signal \TVP_VIDEO_c_5\ : std_logic;
signal \TVP_VIDEO_c_3\ : std_logic;
signal \TVP_VIDEO_c_7\ : std_logic;
signal \TVP_VIDEO_c_6\ : std_logic;
signal \TVP_VIDEO_c_8\ : std_logic;
signal \TVP_VIDEO_c_9\ : std_logic;
signal \TVP_VIDEO_c_2\ : std_logic;
signal \line_buffer.n730\ : std_logic;
signal \line_buffer.n632\ : std_logic;
signal \line_buffer.n762\ : std_logic;
signal \line_buffer.n759\ : std_logic;
signal \line_buffer.n751\ : std_logic;
signal \receive_module.rx_counter.n2975_cascade_\ : std_logic;
signal \line_buffer.n698\ : std_logic;
signal \receive_module.rx_counter.n2900\ : std_logic;
signal \receive_module.rx_counter.n2900_cascade_\ : std_logic;
signal \receive_module.rx_counter.n2943\ : std_logic;
signal \receive_module.rx_counter.n10\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \receive_module.rx_counter.n9\ : std_logic;
signal \receive_module.rx_counter.n2782\ : std_logic;
signal \receive_module.rx_counter.n8\ : std_logic;
signal \receive_module.rx_counter.n2783\ : std_logic;
signal \receive_module.rx_counter.X_3\ : std_logic;
signal \receive_module.rx_counter.n2784\ : std_logic;
signal \receive_module.rx_counter.X_4\ : std_logic;
signal \receive_module.rx_counter.n2785\ : std_logic;
signal \receive_module.rx_counter.X_5\ : std_logic;
signal \receive_module.rx_counter.n2786\ : std_logic;
signal \receive_module.rx_counter.X_6\ : std_logic;
signal \receive_module.rx_counter.n2787\ : std_logic;
signal \receive_module.rx_counter.X_7\ : std_logic;
signal \receive_module.rx_counter.n2788\ : std_logic;
signal \receive_module.rx_counter.n2789\ : std_logic;
signal \receive_module.rx_counter.X_8\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \receive_module.rx_counter.n2790\ : std_logic;
signal \receive_module.rx_counter.X_9\ : std_logic;
signal n3184 : std_logic;
signal \receive_module.rx_counter.n4_cascade_\ : std_logic;
signal \receive_module.rx_counter.n2986_cascade_\ : std_logic;
signal \receive_module.rx_counter.n2989_cascade_\ : std_logic;
signal \receive_module.rx_counter.n31_adj_572\ : std_logic;
signal \receive_module.rx_counter.n7\ : std_logic;
signal \receive_module.rx_counter.n3166\ : std_logic;
signal \receive_module.rx_counter.n2978_cascade_\ : std_logic;
signal \receive_module.rx_counter.n4_adj_571\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \receive_module.rx_counter.n2758\ : std_logic;
signal \receive_module.rx_counter.n2759\ : std_logic;
signal \receive_module.rx_counter.n2760\ : std_logic;
signal \receive_module.rx_counter.n2761\ : std_logic;
signal \receive_module.rx_counter.n2762\ : std_logic;
signal \receive_module.rx_counter.n2763\ : std_logic;
signal \receive_module.rx_counter.n2764\ : std_logic;
signal \receive_module.rx_counter.n2765\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \receive_module.rx_counter.Y_7\ : std_logic;
signal \receive_module.rx_counter.Y_4\ : std_logic;
signal \receive_module.rx_counter.Y_2\ : std_logic;
signal \receive_module.rx_counter.Y_8\ : std_logic;
signal \receive_module.rx_counter.n6_cascade_\ : std_logic;
signal \receive_module.rx_counter.Y_3\ : std_logic;
signal \line_buffer.n723\ : std_logic;
signal \line_buffer.n715\ : std_logic;
signal \transmit_module.video_signal_controller.n2972\ : std_logic;
signal \transmit_module.video_signal_controller.n3014\ : std_logic;
signal \transmit_module.video_signal_controller.n3186_cascade_\ : std_logic;
signal \ADV_HSYNC_c\ : std_logic;
signal \transmit_module.video_signal_controller.n12\ : std_logic;
signal \transmit_module.video_signal_controller.n3182_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n8\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_8\ : std_logic;
signal \line_buffer.n758\ : std_logic;
signal \line_buffer.n750\ : std_logic;
signal \receive_module.n2152\ : std_logic;
signal \TVP_HSYNC_c\ : std_logic;
signal \receive_module.old_HS\ : std_logic;
signal \transmit_module.video_signal_controller.n2484\ : std_logic;
signal \receive_module.rx_counter.Y_5\ : std_logic;
signal \n2147_cascade_\ : std_logic;
signal \receive_module.rx_counter.Y_6\ : std_logic;
signal \Y_0\ : std_logic;
signal \Y_1\ : std_logic;
signal \n5_cascade_\ : std_logic;
signal n3009 : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_0\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_1\ : std_logic;
signal \transmit_module.video_signal_controller.n2766\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_2\ : std_logic;
signal \transmit_module.video_signal_controller.n2767\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_3\ : std_logic;
signal \transmit_module.video_signal_controller.n2768\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_4\ : std_logic;
signal \transmit_module.video_signal_controller.n2769\ : std_logic;
signal \transmit_module.video_signal_controller.n2770\ : std_logic;
signal \transmit_module.video_signal_controller.n2771\ : std_logic;
signal \transmit_module.video_signal_controller.n2772\ : std_logic;
signal \transmit_module.video_signal_controller.n2773\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n2774\ : std_logic;
signal \transmit_module.video_signal_controller.n2775\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_14\ : std_logic;
signal \line_buffer.n754\ : std_logic;
signal \line_buffer.n746\ : std_logic;
signal \line_buffer.n682\ : std_logic;
signal \line_buffer.n3143_cascade_\ : std_logic;
signal \line_buffer.n690\ : std_logic;
signal \line_buffer.n694\ : std_logic;
signal \line_buffer.n686\ : std_logic;
signal \line_buffer.n3101\ : std_logic;
signal \line_buffer.n691\ : std_logic;
signal \line_buffer.n683\ : std_logic;
signal \line_buffer.n722\ : std_logic;
signal \line_buffer.n714\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n2776\ : std_logic;
signal \transmit_module.video_signal_controller.n2777\ : std_logic;
signal \transmit_module.video_signal_controller.n2778\ : std_logic;
signal \transmit_module.video_signal_controller.n2779\ : std_logic;
signal \transmit_module.video_signal_controller.n2780\ : std_logic;
signal \transmit_module.video_signal_controller.n2781\ : std_logic;
signal n2147 : std_logic;
signal \transmit_module.video_signal_controller.n2262\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_0\ : std_logic;
signal \transmit_module.video_signal_controller.n3022_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_8\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_6\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_5\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_7\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_1\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_2\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_5\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_6\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_3\ : std_logic;
signal \line_buffer.n755\ : std_logic;
signal \line_buffer.n747\ : std_logic;
signal \line_buffer.n3031_cascade_\ : std_logic;
signal \line_buffer.n3030\ : std_logic;
signal \line_buffer.n3095_cascade_\ : std_logic;
signal \line_buffer.n3040\ : std_logic;
signal \line_buffer.n625\ : std_logic;
signal \line_buffer.n617\ : std_logic;
signal \line_buffer.n3089\ : std_logic;
signal \line_buffer.n3092_cascade_\ : std_logic;
signal \line_buffer.n3146\ : std_logic;
signal \line_buffer.n626\ : std_logic;
signal \line_buffer.n618\ : std_logic;
signal \line_buffer.n3039\ : std_logic;
signal \receive_module.rx_counter.n10_adj_570_cascade_\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_1\ : std_logic;
signal \receive_module.rx_counter.n2753\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_2\ : std_logic;
signal \receive_module.rx_counter.n2754\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_3\ : std_logic;
signal \receive_module.rx_counter.n2755\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_4\ : std_logic;
signal \receive_module.rx_counter.n2756\ : std_logic;
signal \receive_module.rx_counter.n2757\ : std_logic;
signal \receive_module.rx_counter.n2227\ : std_logic;
signal n1955 : std_logic;
signal \INVADV_R__i1C_net\ : std_logic;
signal \TX_DATA_2\ : std_logic;
signal n1953 : std_logic;
signal \INVADV_R__i3C_net\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_4\ : std_logic;
signal \transmit_module.video_signal_controller.n3183\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_3\ : std_logic;
signal \transmit_module.video_signal_controller.n6\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_9\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_10\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_VISIBLE_N_558_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n18\ : std_logic;
signal \VGA_VISIBLE_cascade_\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_0\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \transmit_module.n2740\ : std_logic;
signal \transmit_module.n2741\ : std_logic;
signal \transmit_module.n2742\ : std_logic;
signal \transmit_module.n2743\ : std_logic;
signal \transmit_module.n2744\ : std_logic;
signal \transmit_module.n2745\ : std_logic;
signal \transmit_module.n2746\ : std_logic;
signal \transmit_module.n2747\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \transmit_module.n2748\ : std_logic;
signal \transmit_module.n2749\ : std_logic;
signal \transmit_module.n2750\ : std_logic;
signal \transmit_module.n2751\ : std_logic;
signal \transmit_module.n2752\ : std_logic;
signal \transmit_module.n2200\ : std_logic;
signal \DEBUG_c_6\ : std_logic;
signal \transmit_module.n382\ : std_logic;
signal n22 : std_logic;
signal \transmit_module.n383\ : std_logic;
signal \DEBUG_c_5\ : std_logic;
signal n23 : std_logic;
signal \transmit_module.n384\ : std_logic;
signal \DEBUG_c_4\ : std_logic;
signal n24 : std_logic;
signal \transmit_module.n386\ : std_logic;
signal \DEBUG_c_2\ : std_logic;
signal n26 : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_5\ : std_logic;
signal \receive_module.rx_counter.n10_adj_570\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_0\ : std_logic;
signal \LED_c\ : std_logic;
signal \receive_module.old_VS\ : std_logic;
signal \receive_module.n252\ : std_logic;
signal n1950 : std_logic;
signal \INVADV_R__i6C_net\ : std_logic;
signal n1954 : std_logic;
signal \TX_DATA_3\ : std_logic;
signal n1952 : std_logic;
signal n1951 : std_logic;
signal n1949 : std_logic;
signal \ADV_B_c\ : std_logic;
signal \INVADV_R__i2C_net\ : std_logic;
signal n19 : std_logic;
signal \transmit_module.n379\ : std_logic;
signal \transmit_module.TX_ADDR_9\ : std_logic;
signal \transmit_module.TX_ADDR_8\ : std_logic;
signal \transmit_module.n380\ : std_logic;
signal n20 : std_logic;
signal \transmit_module.TX_ADDR_10\ : std_logic;
signal \transmit_module.n378\ : std_logic;
signal n18 : std_logic;
signal \line_buffer.n3104\ : std_logic;
signal \TX_DATA_6\ : std_logic;
signal \GB_BUFFER_TVP_CLK_c_THRU_CO\ : std_logic;
signal \line_buffer.n689\ : std_logic;
signal \line_buffer.n681\ : std_logic;
signal \line_buffer.n3140_cascade_\ : std_logic;
signal \TX_DATA_1\ : std_logic;
signal \line_buffer.n713\ : std_logic;
signal \line_buffer.n721\ : std_logic;
signal \line_buffer.n624\ : std_logic;
signal \line_buffer.n616\ : std_logic;
signal \line_buffer.n3107_cascade_\ : std_logic;
signal \line_buffer.n3110\ : std_logic;
signal \line_buffer.n745\ : std_logic;
signal \line_buffer.n753\ : std_logic;
signal \line_buffer.n3137\ : std_logic;
signal \line_buffer.n761\ : std_logic;
signal \transmit_module.n387\ : std_logic;
signal \DEBUG_c_1\ : std_logic;
signal n27 : std_logic;
signal \DEBUG_c_7\ : std_logic;
signal \transmit_module.n381\ : std_logic;
signal n21 : std_logic;
signal \transmit_module.n385\ : std_logic;
signal \DEBUG_c_3\ : std_logic;
signal n25_adj_573 : std_logic;
signal \line_buffer.n3028\ : std_logic;
signal \line_buffer.n3125_cascade_\ : std_logic;
signal \TX_DATA_7\ : std_logic;
signal \line_buffer.n727\ : std_logic;
signal \line_buffer.n719\ : std_logic;
signal \line_buffer.n3043\ : std_logic;
signal \line_buffer.n726\ : std_logic;
signal \line_buffer.n718\ : std_logic;
signal \line_buffer.n629\ : std_logic;
signal \line_buffer.n621\ : std_logic;
signal \line_buffer.n3161_cascade_\ : std_logic;
signal \line_buffer.n3164\ : std_logic;
signal \line_buffer.n630\ : std_logic;
signal \line_buffer.n622\ : std_logic;
signal \line_buffer.n3042\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \line_buffer.n623\ : std_logic;
signal \line_buffer.n615\ : std_logic;
signal \line_buffer.n720\ : std_logic;
signal \line_buffer.n712\ : std_logic;
signal \line_buffer.n3113\ : std_logic;
signal \line_buffer.n688\ : std_logic;
signal \line_buffer.n680\ : std_logic;
signal \line_buffer.n3122_cascade_\ : std_logic;
signal \line_buffer.n3116\ : std_logic;
signal \TX_DATA_0\ : std_logic;
signal \RX_ADDR_0\ : std_logic;
signal \receive_module.n136\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \receive_module.n2727\ : std_logic;
signal \receive_module.n2728\ : std_logic;
signal \receive_module.n2729\ : std_logic;
signal \receive_module.n2730\ : std_logic;
signal \RX_ADDR_5\ : std_logic;
signal \receive_module.n131\ : std_logic;
signal \receive_module.n2731\ : std_logic;
signal \receive_module.n2732\ : std_logic;
signal \RX_ADDR_7\ : std_logic;
signal \receive_module.n129\ : std_logic;
signal \receive_module.n2733\ : std_logic;
signal \receive_module.n2734\ : std_logic;
signal \RX_ADDR_8\ : std_logic;
signal \receive_module.n128\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \RX_ADDR_9\ : std_logic;
signal \receive_module.n127\ : std_logic;
signal \receive_module.n2735\ : std_logic;
signal \receive_module.n2736\ : std_logic;
signal \receive_module.n2737\ : std_logic;
signal \receive_module.n2738\ : std_logic;
signal \receive_module.n2739\ : std_logic;
signal \receive_module.n3181\ : std_logic;
signal \transmit_module.n388\ : std_logic;
signal \ADV_VSYNC_c\ : std_logic;
signal \DEBUG_c_0\ : std_logic;
signal \VGA_VISIBLE\ : std_logic;
signal n28 : std_logic;
signal \line_buffer.n744\ : std_logic;
signal \line_buffer.n752\ : std_logic;
signal \line_buffer.n3119\ : std_logic;
signal \line_buffer.n695\ : std_logic;
signal \line_buffer.n687\ : std_logic;
signal \line_buffer.n3027\ : std_logic;
signal \line_buffer.n725\ : std_logic;
signal \line_buffer.n717\ : std_logic;
signal \receive_module.n133\ : std_logic;
signal \RX_ADDR_3\ : std_logic;
signal \receive_module.n134\ : std_logic;
signal \RX_ADDR_2\ : std_logic;
signal \receive_module.n135\ : std_logic;
signal \RX_ADDR_1\ : std_logic;
signal \line_buffer.n628\ : std_logic;
signal \line_buffer.n620\ : std_logic;
signal \line_buffer.n3149\ : std_logic;
signal \line_buffer.n3152_cascade_\ : std_logic;
signal \TX_DATA_5\ : std_logic;
signal \line_buffer.n692\ : std_logic;
signal \line_buffer.n684\ : std_logic;
signal \line_buffer.n3024\ : std_logic;
signal \line_buffer.n3131_cascade_\ : std_logic;
signal \TX_ADDR_13\ : std_logic;
signal \TX_DATA_4\ : std_logic;
signal \ADV_CLK_c\ : std_logic;
signal \line_buffer.n716\ : std_logic;
signal \line_buffer.n724\ : std_logic;
signal \line_buffer.n3046\ : std_logic;
signal \receive_module.n132\ : std_logic;
signal \RX_ADDR_4\ : std_logic;
signal \receive_module.n130\ : std_logic;
signal \RX_ADDR_6\ : std_logic;
signal \receive_module.n126\ : std_logic;
signal \TVP_VSYNC_c\ : std_logic;
signal \RX_ADDR_10\ : std_logic;
signal \TVP_CLK_c\ : std_logic;
signal \receive_module.n3185\ : std_logic;
signal \line_buffer.n757\ : std_logic;
signal \line_buffer.n749\ : std_logic;
signal \line_buffer.n685\ : std_logic;
signal \line_buffer.n693\ : std_logic;
signal \line_buffer.n3155_cascade_\ : std_logic;
signal \TX_ADDR_12\ : std_logic;
signal \line_buffer.n3158\ : std_logic;
signal \line_buffer.n627\ : std_logic;
signal \line_buffer.n619\ : std_logic;
signal \line_buffer.n3045\ : std_logic;
signal \TX_ADDR_11\ : std_logic;
signal \line_buffer.n756\ : std_logic;
signal \line_buffer.n748\ : std_logic;
signal \line_buffer.n3025\ : std_logic;
signal \line_buffer.n729\ : std_logic;
signal \line_buffer.n697\ : std_logic;
signal \RX_ADDR_12\ : std_logic;
signal \RX_ADDR_11\ : std_logic;
signal \RX_ADDR_13\ : std_logic;
signal n25 : std_logic;
signal \line_buffer.n633\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \TVP_CLK_wire\ : std_logic;
signal \ADV_CLK_wire\ : std_logic;
signal \TVP_VIDEO_wire\ : std_logic_vector(9 downto 0);
signal \ADV_G_wire\ : std_logic_vector(7 downto 0);
signal \ADV_B_wire\ : std_logic_vector(7 downto 0);
signal \ADV_R_wire\ : std_logic_vector(7 downto 0);
signal \ADV_VSYNC_wire\ : std_logic;
signal \ADV_HSYNC_wire\ : std_logic;
signal \ADV_SYNC_N_wire\ : std_logic;
signal \TVP_HSYNC_wire\ : std_logic;
signal \TVP_VSYNC_wire\ : std_logic;
signal \ADV_BLANK_N_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \line_buffer.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \TVP_CLK_wire\ <= TVP_CLK;
    ADV_CLK <= \ADV_CLK_wire\;
    \TVP_VIDEO_wire\ <= TVP_VIDEO;
    ADV_G <= \ADV_G_wire\;
    ADV_B <= \ADV_B_wire\;
    ADV_R <= \ADV_R_wire\;
    ADV_VSYNC <= \ADV_VSYNC_wire\;
    ADV_HSYNC <= \ADV_HSYNC_wire\;
    ADV_SYNC_N <= \ADV_SYNC_N_wire\;
    \TVP_HSYNC_wire\ <= TVP_HSYNC;
    \TVP_VSYNC_wire\ <= TVP_VSYNC;
    ADV_BLANK_N <= \ADV_BLANK_N_wire\;
    LED <= \LED_wire\;
    \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.n630\ <= \line_buffer.mem2_physical_RDATA_wire\(11);
    \line_buffer.n629\ <= \line_buffer.mem2_physical_RDATA_wire\(3);
    \line_buffer.mem2_physical_RADDR_wire\ <= \N__10449\&\N__10983\&\N__10710\&\N__11640\&\N__9738\&\N__9459\&\N__9195\&\N__11364\&\N__8931\&\N__11919\&\N__13905\;
    \line_buffer.mem2_physical_WADDR_wire\ <= \N__16212\&\N__14607\&\N__12846\&\N__13098\&\N__16575\&\N__13341\&\N__16827\&\N__15426\&\N__15177\&\N__14943\&\N__13602\;
    \line_buffer.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6514\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6634\&'0'&'0'&'0';
    \line_buffer.n717\ <= \line_buffer.mem14_physical_RDATA_wire\(11);
    \line_buffer.n716\ <= \line_buffer.mem14_physical_RDATA_wire\(3);
    \line_buffer.mem14_physical_RADDR_wire\ <= \N__10521\&\N__11055\&\N__10782\&\N__11712\&\N__9810\&\N__9531\&\N__9267\&\N__11436\&\N__9003\&\N__11991\&\N__13977\;
    \line_buffer.mem14_physical_WADDR_wire\ <= \N__16284\&\N__14679\&\N__12918\&\N__13170\&\N__16647\&\N__13413\&\N__16899\&\N__15498\&\N__15249\&\N__15015\&\N__13674\;
    \line_buffer.mem14_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem14_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6432\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6304\&'0'&'0'&'0';
    \line_buffer.n620\ <= \line_buffer.mem8_physical_RDATA_wire\(11);
    \line_buffer.n619\ <= \line_buffer.mem8_physical_RDATA_wire\(3);
    \line_buffer.mem8_physical_RADDR_wire\ <= \N__10434\&\N__10962\&\N__10677\&\N__11631\&\N__9717\&\N__9432\&\N__9168\&\N__11343\&\N__8892\&\N__11898\&\N__13884\;
    \line_buffer.mem8_physical_WADDR_wire\ <= \N__16185\&\N__14580\&\N__12819\&\N__13059\&\N__16548\&\N__13320\&\N__16794\&\N__15399\&\N__15162\&\N__14916\&\N__13581\;
    \line_buffer.mem8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem8_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6442\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6324\&'0'&'0'&'0';
    \line_buffer.n721\ <= \line_buffer.mem28_physical_RDATA_wire\(11);
    \line_buffer.n720\ <= \line_buffer.mem28_physical_RDATA_wire\(3);
    \line_buffer.mem28_physical_RADDR_wire\ <= \N__10542\&\N__11070\&\N__10785\&\N__11739\&\N__9825\&\N__9540\&\N__9276\&\N__11451\&\N__9000\&\N__12006\&\N__13992\;
    \line_buffer.mem28_physical_WADDR_wire\ <= \N__16293\&\N__14688\&\N__12927\&\N__13167\&\N__16656\&\N__13428\&\N__16902\&\N__15507\&\N__15270\&\N__15024\&\N__13689\;
    \line_buffer.mem28_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem28_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6171\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6848\&'0'&'0'&'0';
    \line_buffer.n727\ <= \line_buffer.mem5_physical_RDATA_wire\(11);
    \line_buffer.n726\ <= \line_buffer.mem5_physical_RDATA_wire\(3);
    \line_buffer.mem5_physical_RADDR_wire\ <= \N__10470\&\N__10998\&\N__10713\&\N__11667\&\N__9753\&\N__9468\&\N__9204\&\N__11379\&\N__8928\&\N__11934\&\N__13920\;
    \line_buffer.mem5_physical_WADDR_wire\ <= \N__16221\&\N__14616\&\N__12855\&\N__13095\&\N__16584\&\N__13356\&\N__16830\&\N__15435\&\N__15198\&\N__14952\&\N__13617\;
    \line_buffer.mem5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6536\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6647\&'0'&'0'&'0';
    \line_buffer.n685\ <= \line_buffer.mem11_physical_RDATA_wire\(11);
    \line_buffer.n684\ <= \line_buffer.mem11_physical_RDATA_wire\(3);
    \line_buffer.mem11_physical_RADDR_wire\ <= \N__10557\&\N__11091\&\N__10818\&\N__11748\&\N__9846\&\N__9567\&\N__9303\&\N__11472\&\N__9039\&\N__12027\&\N__14013\;
    \line_buffer.mem11_physical_WADDR_wire\ <= \N__16320\&\N__14715\&\N__12954\&\N__13206\&\N__16683\&\N__13449\&\N__16935\&\N__15534\&\N__15285\&\N__15051\&\N__13710\;
    \line_buffer.mem11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem11_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6389\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6283\&'0'&'0'&'0';
    \line_buffer.n747\ <= \line_buffer.mem21_physical_RDATA_wire\(11);
    \line_buffer.n746\ <= \line_buffer.mem21_physical_RDATA_wire\(3);
    \line_buffer.mem21_physical_RADDR_wire\ <= \N__10425\&\N__10959\&\N__10686\&\N__11616\&\N__9714\&\N__9435\&\N__9171\&\N__11340\&\N__8907\&\N__11895\&\N__13881\;
    \line_buffer.mem21_physical_WADDR_wire\ <= \N__16188\&\N__14583\&\N__12822\&\N__13074\&\N__16551\&\N__13317\&\N__16803\&\N__15402\&\N__15153\&\N__14919\&\N__13578\;
    \line_buffer.mem21_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem21_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6112\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6010\&'0'&'0'&'0';
    \line_buffer.n683\ <= \line_buffer.mem12_physical_RDATA_wire\(11);
    \line_buffer.n682\ <= \line_buffer.mem12_physical_RDATA_wire\(3);
    \line_buffer.mem12_physical_RADDR_wire\ <= \N__10545\&\N__11079\&\N__10806\&\N__11736\&\N__9834\&\N__9555\&\N__9291\&\N__11460\&\N__9027\&\N__12015\&\N__14001\;
    \line_buffer.mem12_physical_WADDR_wire\ <= \N__16308\&\N__14703\&\N__12942\&\N__13194\&\N__16671\&\N__13437\&\N__16923\&\N__15522\&\N__15273\&\N__15039\&\N__13698\;
    \line_buffer.mem12_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem12_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6069\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6002\&'0'&'0'&'0';
    \line_buffer.n626\ <= \line_buffer.mem18_physical_RDATA_wire\(11);
    \line_buffer.n625\ <= \line_buffer.mem18_physical_RDATA_wire\(3);
    \line_buffer.mem18_physical_RADDR_wire\ <= \N__10473\&\N__11007\&\N__10734\&\N__11664\&\N__9762\&\N__9483\&\N__9219\&\N__11388\&\N__8955\&\N__11943\&\N__13929\;
    \line_buffer.mem18_physical_WADDR_wire\ <= \N__16236\&\N__14631\&\N__12870\&\N__13122\&\N__16599\&\N__13365\&\N__16851\&\N__15450\&\N__15201\&\N__14967\&\N__13626\;
    \line_buffer.mem18_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem18_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6101\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6003\&'0'&'0'&'0';
    \line_buffer.n691\ <= \line_buffer.mem24_physical_RDATA_wire\(11);
    \line_buffer.n690\ <= \line_buffer.mem24_physical_RDATA_wire\(3);
    \line_buffer.mem24_physical_RADDR_wire\ <= \N__10590\&\N__11118\&\N__10833\&\N__11785\&\N__9873\&\N__9588\&\N__9324\&\N__11499\&\N__9048\&\N__12054\&\N__14040\;
    \line_buffer.mem24_physical_WADDR_wire\ <= \N__16341\&\N__14736\&\N__12975\&\N__13215\&\N__16704\&\N__13476\&\N__16950\&\N__15555\&\N__15318\&\N__15072\&\N__13737\;
    \line_buffer.mem24_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem24_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6038\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5927\&'0'&'0'&'0';
    \line_buffer.n719\ <= \line_buffer.mem1_physical_RDATA_wire\(11);
    \line_buffer.n718\ <= \line_buffer.mem1_physical_RDATA_wire\(3);
    \line_buffer.mem1_physical_RADDR_wire\ <= \N__10581\&\N__11115\&\N__10842\&\N__11772\&\N__9870\&\N__9591\&\N__9327\&\N__11496\&\N__9061\&\N__12051\&\N__14037\;
    \line_buffer.mem1_physical_WADDR_wire\ <= \N__16344\&\N__14739\&\N__12978\&\N__13228\&\N__16707\&\N__13473\&\N__16959\&\N__15558\&\N__15309\&\N__15075\&\N__13734\;
    \line_buffer.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6493\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6608\&'0'&'0'&'0';
    \line_buffer.n715\ <= \line_buffer.mem15_physical_RDATA_wire\(11);
    \line_buffer.n714\ <= \line_buffer.mem15_physical_RDATA_wire\(3);
    \line_buffer.mem15_physical_RADDR_wire\ <= \N__10509\&\N__11043\&\N__10770\&\N__11700\&\N__9798\&\N__9519\&\N__9255\&\N__11424\&\N__8991\&\N__11979\&\N__13965\;
    \line_buffer.mem15_physical_WADDR_wire\ <= \N__16272\&\N__14667\&\N__12906\&\N__13158\&\N__16635\&\N__13401\&\N__16887\&\N__15486\&\N__15237\&\N__15003\&\N__13662\;
    \line_buffer.mem15_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem15_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6082\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5994\&'0'&'0'&'0';
    \line_buffer.n723\ <= \line_buffer.mem27_physical_RDATA_wire\(11);
    \line_buffer.n722\ <= \line_buffer.mem27_physical_RDATA_wire\(3);
    \line_buffer.mem27_physical_RADDR_wire\ <= \N__10554\&\N__11082\&\N__10797\&\N__11751\&\N__9837\&\N__9552\&\N__9288\&\N__11463\&\N__9012\&\N__12018\&\N__14004\;
    \line_buffer.mem27_physical_WADDR_wire\ <= \N__16305\&\N__14700\&\N__12939\&\N__13179\&\N__16668\&\N__13440\&\N__16914\&\N__15519\&\N__15282\&\N__15036\&\N__13701\;
    \line_buffer.mem27_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem27_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6063\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5958\&'0'&'0'&'0';
    \line_buffer.n745\ <= \line_buffer.mem22_physical_RDATA_wire\(11);
    \line_buffer.n744\ <= \line_buffer.mem22_physical_RDATA_wire\(3);
    \line_buffer.mem22_physical_RADDR_wire\ <= \N__10413\&\N__10947\&\N__10674\&\N__11604\&\N__9702\&\N__9423\&\N__9159\&\N__11328\&\N__8895\&\N__11883\&\N__13869\;
    \line_buffer.mem22_physical_WADDR_wire\ <= \N__16176\&\N__14571\&\N__12810\&\N__13062\&\N__16539\&\N__13305\&\N__16791\&\N__15390\&\N__15141\&\N__14907\&\N__13566\;
    \line_buffer.mem22_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem22_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6223\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6907\&'0'&'0'&'0';
    \line_buffer.n695\ <= \line_buffer.mem4_physical_RDATA_wire\(11);
    \line_buffer.n694\ <= \line_buffer.mem4_physical_RDATA_wire\(3);
    \line_buffer.mem4_physical_RADDR_wire\ <= \N__10482\&\N__11010\&\N__10725\&\N__11679\&\N__9765\&\N__9480\&\N__9216\&\N__11391\&\N__8940\&\N__11946\&\N__13932\;
    \line_buffer.mem4_physical_WADDR_wire\ <= \N__16233\&\N__14628\&\N__12867\&\N__13107\&\N__16596\&\N__13368\&\N__16842\&\N__15447\&\N__15210\&\N__14964\&\N__13629\;
    \line_buffer.mem4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6521\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6646\&'0'&'0'&'0';
    \line_buffer.n713\ <= \line_buffer.mem16_physical_RDATA_wire\(11);
    \line_buffer.n712\ <= \line_buffer.mem16_physical_RDATA_wire\(3);
    \line_buffer.mem16_physical_RADDR_wire\ <= \N__10497\&\N__11031\&\N__10758\&\N__11688\&\N__9786\&\N__9507\&\N__9243\&\N__11412\&\N__8979\&\N__11967\&\N__13953\;
    \line_buffer.mem16_physical_WADDR_wire\ <= \N__16260\&\N__14655\&\N__12894\&\N__13146\&\N__16623\&\N__13389\&\N__16875\&\N__15474\&\N__15225\&\N__14991\&\N__13650\;
    \line_buffer.mem16_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem16_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6222\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6888\&'0'&'0'&'0';
    \line_buffer.n755\ <= \line_buffer.mem30_physical_RDATA_wire\(11);
    \line_buffer.n754\ <= \line_buffer.mem30_physical_RDATA_wire\(3);
    \line_buffer.mem30_physical_RADDR_wire\ <= \N__10506\&\N__11034\&\N__10749\&\N__11703\&\N__9789\&\N__9504\&\N__9240\&\N__11415\&\N__8964\&\N__11970\&\N__13956\;
    \line_buffer.mem30_physical_WADDR_wire\ <= \N__16257\&\N__14652\&\N__12891\&\N__13131\&\N__16620\&\N__13392\&\N__16866\&\N__15471\&\N__15234\&\N__14988\&\N__13653\;
    \line_buffer.mem30_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem30_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6088\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5990\&'0'&'0'&'0';
    \line_buffer.n689\ <= \line_buffer.mem25_physical_RDATA_wire\(11);
    \line_buffer.n688\ <= \line_buffer.mem25_physical_RDATA_wire\(3);
    \line_buffer.mem25_physical_RADDR_wire\ <= \N__10578\&\N__11106\&\N__10821\&\N__11775\&\N__9861\&\N__9576\&\N__9312\&\N__11487\&\N__9036\&\N__12042\&\N__14028\;
    \line_buffer.mem25_physical_WADDR_wire\ <= \N__16329\&\N__14724\&\N__12963\&\N__13203\&\N__16692\&\N__13464\&\N__16938\&\N__15543\&\N__15306\&\N__15060\&\N__13725\;
    \line_buffer.mem25_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem25_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6190\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6835\&'0'&'0'&'0';
    \line_buffer.n622\ <= \line_buffer.mem7_physical_RDATA_wire\(11);
    \line_buffer.n621\ <= \line_buffer.mem7_physical_RDATA_wire\(3);
    \line_buffer.mem7_physical_RADDR_wire\ <= \N__10446\&\N__10974\&\N__10689\&\N__11643\&\N__9729\&\N__9444\&\N__9180\&\N__11355\&\N__8904\&\N__11910\&\N__13896\;
    \line_buffer.mem7_physical_WADDR_wire\ <= \N__16197\&\N__14592\&\N__12831\&\N__13071\&\N__16560\&\N__13332\&\N__16806\&\N__15411\&\N__15174\&\N__14928\&\N__13593\;
    \line_buffer.mem7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem7_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6544\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6655\&'0'&'0'&'0';
    \line_buffer.n749\ <= \line_buffer.mem20_physical_RDATA_wire\(11);
    \line_buffer.n748\ <= \line_buffer.mem20_physical_RDATA_wire\(3);
    \line_buffer.mem20_physical_RADDR_wire\ <= \N__10437\&\N__10971\&\N__10698\&\N__11628\&\N__9726\&\N__9447\&\N__9183\&\N__11352\&\N__8919\&\N__11907\&\N__13893\;
    \line_buffer.mem20_physical_WADDR_wire\ <= \N__16200\&\N__14595\&\N__12834\&\N__13086\&\N__16563\&\N__13329\&\N__16815\&\N__15414\&\N__15165\&\N__14931\&\N__13590\;
    \line_buffer.mem20_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem20_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6440\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6325\&'0'&'0'&'0';
    \line_buffer.n681\ <= \line_buffer.mem13_physical_RDATA_wire\(11);
    \line_buffer.n680\ <= \line_buffer.mem13_physical_RDATA_wire\(3);
    \line_buffer.mem13_physical_RADDR_wire\ <= \N__10533\&\N__11067\&\N__10794\&\N__11724\&\N__9822\&\N__9543\&\N__9279\&\N__11448\&\N__9015\&\N__12003\&\N__13989\;
    \line_buffer.mem13_physical_WADDR_wire\ <= \N__16296\&\N__14691\&\N__12930\&\N__13182\&\N__16659\&\N__13425\&\N__16911\&\N__15510\&\N__15261\&\N__15027\&\N__13686\;
    \line_buffer.mem13_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem13_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6191\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6881\&'0'&'0'&'0';
    \line_buffer.n624\ <= \line_buffer.mem19_physical_RDATA_wire\(11);
    \line_buffer.n623\ <= \line_buffer.mem19_physical_RDATA_wire\(3);
    \line_buffer.mem19_physical_RADDR_wire\ <= \N__10461\&\N__10995\&\N__10722\&\N__11652\&\N__9750\&\N__9471\&\N__9207\&\N__11376\&\N__8943\&\N__11931\&\N__13917\;
    \line_buffer.mem19_physical_WADDR_wire\ <= \N__16224\&\N__14619\&\N__12858\&\N__13110\&\N__16587\&\N__13353\&\N__16839\&\N__15438\&\N__15189\&\N__14955\&\N__13614\;
    \line_buffer.mem19_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem19_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6205\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6900\&'0'&'0'&'0';
    \line_buffer.n693\ <= \line_buffer.mem23_physical_RDATA_wire\(11);
    \line_buffer.n692\ <= \line_buffer.mem23_physical_RDATA_wire\(3);
    \line_buffer.mem23_physical_RADDR_wire\ <= \N__10597\&\N__11128\&\N__10845\&\N__11791\&\N__9883\&\N__9600\&\N__9336\&\N__11509\&\N__9060\&\N__12064\&\N__14050\;
    \line_buffer.mem23_physical_WADDR_wire\ <= \N__16353\&\N__14748\&\N__12987\&\N__13227\&\N__16716\&\N__13486\&\N__16962\&\N__15567\&\N__15325\&\N__15084\&\N__13747\;
    \line_buffer.mem23_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem23_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6402\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6251\&'0'&'0'&'0';
    \line_buffer.n687\ <= \line_buffer.mem0_physical_RDATA_wire\(11);
    \line_buffer.n686\ <= \line_buffer.mem0_physical_RDATA_wire\(3);
    \line_buffer.mem0_physical_RADDR_wire\ <= \N__10593\&\N__11127\&\N__10849\&\N__11784\&\N__9882\&\N__9601\&\N__9337\&\N__11508\&\N__9067\&\N__12063\&\N__14049\;
    \line_buffer.mem0_physical_WADDR_wire\ <= \N__16354\&\N__14749\&\N__12988\&\N__13234\&\N__16717\&\N__13485\&\N__16966\&\N__15568\&\N__15321\&\N__15085\&\N__13746\;
    \line_buffer.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6468\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6607\&'0'&'0'&'0';
    \line_buffer.n725\ <= \line_buffer.mem26_physical_RDATA_wire\(11);
    \line_buffer.n724\ <= \line_buffer.mem26_physical_RDATA_wire\(3);
    \line_buffer.mem26_physical_RADDR_wire\ <= \N__10566\&\N__11094\&\N__10809\&\N__11763\&\N__9849\&\N__9564\&\N__9300\&\N__11475\&\N__9024\&\N__12030\&\N__14016\;
    \line_buffer.mem26_physical_WADDR_wire\ <= \N__16317\&\N__14712\&\N__12951\&\N__13191\&\N__16680\&\N__13452\&\N__16926\&\N__15531\&\N__15294\&\N__15048\&\N__13713\;
    \line_buffer.mem26_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem26_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6388\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6276\&'0'&'0'&'0';
    \line_buffer.n751\ <= \line_buffer.mem3_physical_RDATA_wire\(11);
    \line_buffer.n750\ <= \line_buffer.mem3_physical_RDATA_wire\(3);
    \line_buffer.mem3_physical_RADDR_wire\ <= \N__10518\&\N__11046\&\N__10761\&\N__11715\&\N__9801\&\N__9516\&\N__9252\&\N__11427\&\N__8976\&\N__11982\&\N__13968\;
    \line_buffer.mem3_physical_WADDR_wire\ <= \N__16269\&\N__14664\&\N__12903\&\N__13143\&\N__16632\&\N__13404\&\N__16878\&\N__15483\&\N__15246\&\N__15000\&\N__13665\;
    \line_buffer.mem3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6522\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6626\&'0'&'0'&'0';
    \line_buffer.n628\ <= \line_buffer.mem17_physical_RDATA_wire\(11);
    \line_buffer.n627\ <= \line_buffer.mem17_physical_RDATA_wire\(3);
    \line_buffer.mem17_physical_RADDR_wire\ <= \N__10485\&\N__11019\&\N__10746\&\N__11676\&\N__9774\&\N__9495\&\N__9231\&\N__11400\&\N__8967\&\N__11955\&\N__13941\;
    \line_buffer.mem17_physical_WADDR_wire\ <= \N__16248\&\N__14643\&\N__12882\&\N__13134\&\N__16611\&\N__13377\&\N__16863\&\N__15462\&\N__15213\&\N__14979\&\N__13638\;
    \line_buffer.mem17_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem17_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6441\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6314\&'0'&'0'&'0';
    \line_buffer.n753\ <= \line_buffer.mem31_physical_RDATA_wire\(11);
    \line_buffer.n752\ <= \line_buffer.mem31_physical_RDATA_wire\(3);
    \line_buffer.mem31_physical_RADDR_wire\ <= \N__10494\&\N__11022\&\N__10737\&\N__11691\&\N__9777\&\N__9492\&\N__9228\&\N__11403\&\N__8952\&\N__11958\&\N__13944\;
    \line_buffer.mem31_physical_WADDR_wire\ <= \N__16245\&\N__14640\&\N__12879\&\N__13119\&\N__16608\&\N__13380\&\N__16854\&\N__15459\&\N__15222\&\N__14976\&\N__13641\;
    \line_buffer.mem31_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem31_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6195\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6866\&'0'&'0'&'0';
    \line_buffer.n618\ <= \line_buffer.mem9_physical_RDATA_wire\(11);
    \line_buffer.n617\ <= \line_buffer.mem9_physical_RDATA_wire\(3);
    \line_buffer.mem9_physical_RADDR_wire\ <= \N__10422\&\N__10950\&\N__10665\&\N__11619\&\N__9705\&\N__9420\&\N__9156\&\N__11331\&\N__8880\&\N__11886\&\N__13872\;
    \line_buffer.mem9_physical_WADDR_wire\ <= \N__16173\&\N__14568\&\N__12807\&\N__13047\&\N__16536\&\N__13308\&\N__16782\&\N__15387\&\N__15150\&\N__14904\&\N__13569\;
    \line_buffer.mem9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem9_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6111\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6001\&'0'&'0'&'0';
    \line_buffer.n757\ <= \line_buffer.mem29_physical_RDATA_wire\(11);
    \line_buffer.n756\ <= \line_buffer.mem29_physical_RDATA_wire\(3);
    \line_buffer.mem29_physical_RADDR_wire\ <= \N__10530\&\N__11058\&\N__10773\&\N__11727\&\N__9813\&\N__9528\&\N__9264\&\N__11439\&\N__8988\&\N__11994\&\N__13980\;
    \line_buffer.mem29_physical_WADDR_wire\ <= \N__16281\&\N__14676\&\N__12915\&\N__13155\&\N__16644\&\N__13416\&\N__16890\&\N__15495\&\N__15258\&\N__15012\&\N__13677\;
    \line_buffer.mem29_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem29_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6436\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6289\&'0'&'0'&'0';
    \line_buffer.n759\ <= \line_buffer.mem6_physical_RDATA_wire\(11);
    \line_buffer.n758\ <= \line_buffer.mem6_physical_RDATA_wire\(3);
    \line_buffer.mem6_physical_RADDR_wire\ <= \N__10458\&\N__10986\&\N__10701\&\N__11655\&\N__9741\&\N__9456\&\N__9192\&\N__11367\&\N__8916\&\N__11922\&\N__13908\;
    \line_buffer.mem6_physical_WADDR_wire\ <= \N__16209\&\N__14604\&\N__12843\&\N__13083\&\N__16572\&\N__13344\&\N__16818\&\N__15423\&\N__15186\&\N__14940\&\N__13605\;
    \line_buffer.mem6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6543\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6654\&'0'&'0'&'0';
    \line_buffer.n616\ <= \line_buffer.mem10_physical_RDATA_wire\(11);
    \line_buffer.n615\ <= \line_buffer.mem10_physical_RDATA_wire\(3);
    \line_buffer.mem10_physical_RADDR_wire\ <= \N__10569\&\N__11103\&\N__10830\&\N__11760\&\N__9858\&\N__9579\&\N__9315\&\N__11484\&\N__9051\&\N__12039\&\N__14025\;
    \line_buffer.mem10_physical_WADDR_wire\ <= \N__16332\&\N__14727\&\N__12966\&\N__13218\&\N__16695\&\N__13461\&\N__16947\&\N__15546\&\N__15297\&\N__15063\&\N__13722\;
    \line_buffer.mem10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem10_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__6215\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__6867\&'0'&'0'&'0';

    \tx_pll.TX_PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0100110",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \ADV_CLK_c\,
            REFERENCECLK => \N__10366\,
            RESETB => \N__12536\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \line_buffer.mem2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem2_physical_RDATA_wire\,
            RADDR => \line_buffer.mem2_physical_RADDR_wire\,
            WADDR => \line_buffer.mem2_physical_WADDR_wire\,
            MASK => \line_buffer.mem2_physical_MASK_wire\,
            WDATA => \line_buffer.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17397\,
            RE => \N__12569\,
            WCLKE => 'H',
            WCLK => \N__16118\,
            WE => \N__17737\
        );

    \line_buffer.mem14_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem14_physical_RDATA_wire\,
            RADDR => \line_buffer.mem14_physical_RADDR_wire\,
            WADDR => \line_buffer.mem14_physical_WADDR_wire\,
            MASK => \line_buffer.mem14_physical_MASK_wire\,
            WDATA => \line_buffer.mem14_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17531\,
            RE => \N__12471\,
            WCLKE => 'H',
            WCLK => \N__16102\,
            WE => \N__18235\
        );

    \line_buffer.mem8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem8_physical_RDATA_wire\,
            RADDR => \line_buffer.mem8_physical_RADDR_wire\,
            WADDR => \line_buffer.mem8_physical_WADDR_wire\,
            MASK => \line_buffer.mem8_physical_MASK_wire\,
            WDATA => \line_buffer.mem8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17245\,
            RE => \N__12627\,
            WCLKE => 'H',
            WCLK => \N__16123\,
            WE => \N__6746\
        );

    \line_buffer.mem28_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem28_physical_RDATA_wire\,
            RADDR => \line_buffer.mem28_physical_RADDR_wire\,
            WADDR => \line_buffer.mem28_physical_WADDR_wire\,
            MASK => \line_buffer.mem28_physical_MASK_wire\,
            WDATA => \line_buffer.mem28_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17268\,
            RE => \N__12553\,
            WCLKE => 'H',
            WCLK => \N__16100\,
            WE => \N__6764\
        );

    \line_buffer.mem5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem5_physical_RDATA_wire\,
            RADDR => \line_buffer.mem5_physical_RADDR_wire\,
            WADDR => \line_buffer.mem5_physical_WADDR_wire\,
            MASK => \line_buffer.mem5_physical_MASK_wire\,
            WDATA => \line_buffer.mem5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17213\,
            RE => \N__12615\,
            WCLKE => 'H',
            WCLK => \N__16114\,
            WE => \N__6796\
        );

    \line_buffer.mem11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem11_physical_RDATA_wire\,
            RADDR => \line_buffer.mem11_physical_RADDR_wire\,
            WADDR => \line_buffer.mem11_physical_WADDR_wire\,
            MASK => \line_buffer.mem11_physical_MASK_wire\,
            WDATA => \line_buffer.mem11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17579\,
            RE => \N__12436\,
            WCLKE => 'H',
            WCLK => \N__16088\,
            WE => \N__18192\
        );

    \line_buffer.mem21_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem21_physical_RDATA_wire\,
            RADDR => \line_buffer.mem21_physical_RADDR_wire\,
            WADDR => \line_buffer.mem21_physical_WADDR_wire\,
            MASK => \line_buffer.mem21_physical_MASK_wire\,
            WDATA => \line_buffer.mem21_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17313\,
            RE => \N__12595\,
            WCLKE => 'H',
            WCLK => \N__16122\,
            WE => \N__12161\
        );

    \line_buffer.mem12_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem12_physical_RDATA_wire\,
            RADDR => \line_buffer.mem12_physical_RADDR_wire\,
            WADDR => \line_buffer.mem12_physical_WADDR_wire\,
            MASK => \line_buffer.mem12_physical_MASK_wire\,
            WDATA => \line_buffer.mem12_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17559\,
            RE => \N__12437\,
            WCLKE => 'H',
            WCLK => \N__16095\,
            WE => \N__18191\
        );

    \line_buffer.mem18_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem18_physical_RDATA_wire\,
            RADDR => \line_buffer.mem18_physical_RADDR_wire\,
            WADDR => \line_buffer.mem18_physical_WADDR_wire\,
            MASK => \line_buffer.mem18_physical_MASK_wire\,
            WDATA => \line_buffer.mem18_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17457\,
            RE => \N__12539\,
            WCLKE => 'H',
            WCLK => \N__16111\,
            WE => \N__17729\
        );

    \line_buffer.mem24_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem24_physical_RDATA_wire\,
            RADDR => \line_buffer.mem24_physical_RADDR_wire\,
            WADDR => \line_buffer.mem24_physical_WADDR_wire\,
            MASK => \line_buffer.mem24_physical_MASK_wire\,
            WDATA => \line_buffer.mem24_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17587\,
            RE => \N__12485\,
            WCLKE => 'H',
            WCLK => \N__16083\,
            WE => \N__6993\
        );

    \line_buffer.mem1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem1_physical_RDATA_wire\,
            RADDR => \line_buffer.mem1_physical_RADDR_wire\,
            WADDR => \line_buffer.mem1_physical_WADDR_wire\,
            MASK => \line_buffer.mem1_physical_MASK_wire\,
            WDATA => \line_buffer.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17589\,
            RE => \N__12408\,
            WCLKE => 'H',
            WCLK => \N__16081\,
            WE => \N__18244\
        );

    \line_buffer.mem15_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem15_physical_RDATA_wire\,
            RADDR => \line_buffer.mem15_physical_RADDR_wire\,
            WADDR => \line_buffer.mem15_physical_WADDR_wire\,
            MASK => \line_buffer.mem15_physical_MASK_wire\,
            WDATA => \line_buffer.mem15_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17530\,
            RE => \N__12506\,
            WCLKE => 'H',
            WCLK => \N__16105\,
            WE => \N__18236\
        );

    \line_buffer.mem27_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem27_physical_RDATA_wire\,
            RADDR => \line_buffer.mem27_physical_RADDR_wire\,
            WADDR => \line_buffer.mem27_physical_WADDR_wire\,
            MASK => \line_buffer.mem27_physical_MASK_wire\,
            WDATA => \line_buffer.mem27_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17548\,
            RE => \N__12522\,
            WCLKE => 'H',
            WCLK => \N__16098\,
            WE => \N__6788\
        );

    \line_buffer.mem22_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem22_physical_RDATA_wire\,
            RADDR => \line_buffer.mem22_physical_RADDR_wire\,
            WADDR => \line_buffer.mem22_physical_WADDR_wire\,
            MASK => \line_buffer.mem22_physical_MASK_wire\,
            WDATA => \line_buffer.mem22_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17226\,
            RE => \N__12614\,
            WCLKE => 'H',
            WCLK => \N__16124\,
            WE => \N__12166\
        );

    \line_buffer.mem4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem4_physical_RDATA_wire\,
            RADDR => \line_buffer.mem4_physical_RADDR_wire\,
            WADDR => \line_buffer.mem4_physical_WADDR_wire\,
            MASK => \line_buffer.mem4_physical_MASK_wire\,
            WDATA => \line_buffer.mem4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17425\,
            RE => \N__12600\,
            WCLKE => 'H',
            WCLK => \N__16112\,
            WE => \N__6992\
        );

    \line_buffer.mem16_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem16_physical_RDATA_wire\,
            RADDR => \line_buffer.mem16_physical_RADDR_wire\,
            WADDR => \line_buffer.mem16_physical_WADDR_wire\,
            MASK => \line_buffer.mem16_physical_MASK_wire\,
            WDATA => \line_buffer.mem16_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17499\,
            RE => \N__12507\,
            WCLKE => 'H',
            WCLK => \N__16107\,
            WE => \N__18243\
        );

    \line_buffer.mem30_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem30_physical_RDATA_wire\,
            RADDR => \line_buffer.mem30_physical_RADDR_wire\,
            WADDR => \line_buffer.mem30_physical_WADDR_wire\,
            MASK => \line_buffer.mem30_physical_MASK_wire\,
            WDATA => \line_buffer.mem30_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17481\,
            RE => \N__12580\,
            WCLKE => 'H',
            WCLK => \N__16108\,
            WE => \N__6691\
        );

    \line_buffer.mem25_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem25_physical_RDATA_wire\,
            RADDR => \line_buffer.mem25_physical_RADDR_wire\,
            WADDR => \line_buffer.mem25_physical_WADDR_wire\,
            MASK => \line_buffer.mem25_physical_MASK_wire\,
            WDATA => \line_buffer.mem25_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17572\,
            RE => \N__12486\,
            WCLKE => 'H',
            WCLK => \N__16086\,
            WE => \N__6985\
        );

    \line_buffer.mem7_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem7_physical_RDATA_wire\,
            RADDR => \line_buffer.mem7_physical_RADDR_wire\,
            WADDR => \line_buffer.mem7_physical_WADDR_wire\,
            MASK => \line_buffer.mem7_physical_MASK_wire\,
            WDATA => \line_buffer.mem7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17225\,
            RE => \N__12626\,
            WCLKE => 'H',
            WCLK => \N__16121\,
            WE => \N__6736\
        );

    \line_buffer.mem20_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem20_physical_RDATA_wire\,
            RADDR => \line_buffer.mem20_physical_RADDR_wire\,
            WADDR => \line_buffer.mem20_physical_WADDR_wire\,
            MASK => \line_buffer.mem20_physical_MASK_wire\,
            WDATA => \line_buffer.mem20_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17396\,
            RE => \N__12594\,
            WCLKE => 'H',
            WCLK => \N__16120\,
            WE => \N__12160\
        );

    \line_buffer.mem13_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem13_physical_RDATA_wire\,
            RADDR => \line_buffer.mem13_physical_RADDR_wire\,
            WADDR => \line_buffer.mem13_physical_WADDR_wire\,
            MASK => \line_buffer.mem13_physical_MASK_wire\,
            WDATA => \line_buffer.mem13_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17558\,
            RE => \N__12470\,
            WCLKE => 'H',
            WCLK => \N__16099\,
            WE => \N__18184\
        );

    \line_buffer.mem19_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem19_physical_RDATA_wire\,
            RADDR => \line_buffer.mem19_physical_RADDR_wire\,
            WADDR => \line_buffer.mem19_physical_WADDR_wire\,
            MASK => \line_buffer.mem19_physical_MASK_wire\,
            WDATA => \line_buffer.mem19_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17311\,
            RE => \N__12568\,
            WCLKE => 'H',
            WCLK => \N__16113\,
            WE => \N__17736\
        );

    \line_buffer.mem23_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem23_physical_RDATA_wire\,
            RADDR => \line_buffer.mem23_physical_RADDR_wire\,
            WADDR => \line_buffer.mem23_physical_WADDR_wire\,
            MASK => \line_buffer.mem23_physical_MASK_wire\,
            WDATA => \line_buffer.mem23_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17588\,
            RE => \N__12451\,
            WCLKE => 'H',
            WCLK => \N__16079\,
            WE => \N__6994\
        );

    \line_buffer.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem0_physical_RDATA_wire\,
            RADDR => \line_buffer.mem0_physical_RADDR_wire\,
            WADDR => \line_buffer.mem0_physical_WADDR_wire\,
            MASK => \line_buffer.mem0_physical_MASK_wire\,
            WDATA => \line_buffer.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17590\,
            RE => \N__12407\,
            WCLKE => 'H',
            WCLK => \N__16078\,
            WE => \N__18199\
        );

    \line_buffer.mem26_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem26_physical_RDATA_wire\,
            RADDR => \line_buffer.mem26_physical_RADDR_wire\,
            WADDR => \line_buffer.mem26_physical_WADDR_wire\,
            MASK => \line_buffer.mem26_physical_MASK_wire\,
            WDATA => \line_buffer.mem26_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17327\,
            RE => \N__12521\,
            WCLKE => 'H',
            WCLK => \N__16091\,
            WE => \N__6795\
        );

    \line_buffer.mem3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem3_physical_RDATA_wire\,
            RADDR => \line_buffer.mem3_physical_RADDR_wire\,
            WADDR => \line_buffer.mem3_physical_WADDR_wire\,
            MASK => \line_buffer.mem3_physical_MASK_wire\,
            WDATA => \line_buffer.mem3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17529\,
            RE => \N__12579\,
            WCLKE => 'H',
            WCLK => \N__16106\,
            WE => \N__12165\
        );

    \line_buffer.mem17_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem17_physical_RDATA_wire\,
            RADDR => \line_buffer.mem17_physical_RADDR_wire\,
            WADDR => \line_buffer.mem17_physical_WADDR_wire\,
            MASK => \line_buffer.mem17_physical_MASK_wire\,
            WDATA => \line_buffer.mem17_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17498\,
            RE => \N__12538\,
            WCLKE => 'H',
            WCLK => \N__16109\,
            WE => \N__17712\
        );

    \line_buffer.mem31_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem31_physical_RDATA_wire\,
            RADDR => \line_buffer.mem31_physical_RADDR_wire\,
            WADDR => \line_buffer.mem31_physical_WADDR_wire\,
            MASK => \line_buffer.mem31_physical_MASK_wire\,
            WDATA => \line_buffer.mem31_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17241\,
            RE => \N__12599\,
            WCLKE => 'H',
            WCLK => \N__16110\,
            WE => \N__6692\
        );

    \line_buffer.mem9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem9_physical_RDATA_wire\,
            RADDR => \line_buffer.mem9_physical_RADDR_wire\,
            WADDR => \line_buffer.mem9_physical_WADDR_wire\,
            MASK => \line_buffer.mem9_physical_MASK_wire\,
            WDATA => \line_buffer.mem9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17151\,
            RE => \N__12631\,
            WCLKE => 'H',
            WCLK => \N__16125\,
            WE => \N__6747\
        );

    \line_buffer.mem29_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem29_physical_RDATA_wire\,
            RADDR => \line_buffer.mem29_physical_RADDR_wire\,
            WADDR => \line_buffer.mem29_physical_WADDR_wire\,
            MASK => \line_buffer.mem29_physical_MASK_wire\,
            WDATA => \line_buffer.mem29_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17518\,
            RE => \N__12554\,
            WCLKE => 'H',
            WCLK => \N__16104\,
            WE => \N__6696\
        );

    \line_buffer.mem6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem6_physical_RDATA_wire\,
            RADDR => \line_buffer.mem6_physical_RADDR_wire\,
            WADDR => \line_buffer.mem6_physical_WADDR_wire\,
            MASK => \line_buffer.mem6_physical_MASK_wire\,
            WDATA => \line_buffer.mem6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17328\,
            RE => \N__12616\,
            WCLKE => 'H',
            WCLK => \N__16119\,
            WE => \N__6700\
        );

    \line_buffer.mem10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem10_physical_RDATA_wire\,
            RADDR => \line_buffer.mem10_physical_RADDR_wire\,
            WADDR => \line_buffer.mem10_physical_WADDR_wire\,
            MASK => \line_buffer.mem10_physical_MASK_wire\,
            WDATA => \line_buffer.mem10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17580\,
            RE => \N__12409\,
            WCLKE => 'H',
            WCLK => \N__16085\,
            WE => \N__6751\
        );

    \TVP_CLK_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__18941\,
            GLOBALBUFFEROUTPUT => \TVP_CLK_c\
        );

    \TVP_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18943\,
            DIN => \N__18942\,
            DOUT => \N__18941\,
            PACKAGEPIN => \TVP_CLK_wire\
        );

    \TVP_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18943\,
            PADOUT => \N__18942\,
            PADIN => \N__18941\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18932\,
            DIN => \N__18931\,
            DOUT => \N__18930\,
            PACKAGEPIN => \ADV_CLK_wire\
        );

    \ADV_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18932\,
            PADOUT => \N__18931\,
            PADIN => \N__18930\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17312\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18923\,
            DIN => \N__18922\,
            DOUT => \N__18921\,
            PACKAGEPIN => DEBUG(3)
        );

    \DEBUG_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18923\,
            PADOUT => \N__18922\,
            PADIN => \N__18921\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11557\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18914\,
            DIN => \N__18913\,
            DOUT => \N__18912\,
            PACKAGEPIN => \TVP_VIDEO_wire\(2)
        );

    \TVP_VIDEO_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18914\,
            PADOUT => \N__18913\,
            PADIN => \N__18912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18905\,
            DIN => \N__18904\,
            DOUT => \N__18903\,
            PACKAGEPIN => \ADV_G_wire\(5)
        );

    \ADV_G_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18905\,
            PADOUT => \N__18904\,
            PADIN => \N__18903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10311\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18896\,
            DIN => \N__18895\,
            DOUT => \N__18894\,
            PACKAGEPIN => \ADV_B_wire\(3)
        );

    \ADV_B_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18896\,
            PADOUT => \N__18895\,
            PADIN => \N__18894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10197\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18887\,
            DIN => \N__18886\,
            DOUT => \N__18885\,
            PACKAGEPIN => \ADV_R_wire\(4)
        );

    \ADV_R_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18887\,
            PADOUT => \N__18886\,
            PADIN => \N__18885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10127\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18878\,
            DIN => \N__18877\,
            DOUT => \N__18876\,
            PACKAGEPIN => \TVP_VIDEO_wire\(8)
        );

    \TVP_VIDEO_pad_8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18878\,
            PADOUT => \N__18877\,
            PADIN => \N__18876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18869\,
            DIN => \N__18868\,
            DOUT => \N__18867\,
            PACKAGEPIN => \ADV_B_wire\(0)
        );

    \ADV_B_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18869\,
            PADOUT => \N__18868\,
            PADIN => \N__18867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8502\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18860\,
            DIN => \N__18859\,
            DOUT => \N__18858\,
            PACKAGEPIN => \TVP_VIDEO_wire\(5)
        );

    \TVP_VIDEO_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18860\,
            PADOUT => \N__18859\,
            PADIN => \N__18858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18851\,
            DIN => \N__18850\,
            DOUT => \N__18849\,
            PACKAGEPIN => \ADV_G_wire\(2)
        );

    \ADV_G_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18851\,
            PADOUT => \N__18850\,
            PADIN => \N__18849\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8433\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18842\,
            DIN => \N__18841\,
            DOUT => \N__18840\,
            PACKAGEPIN => \ADV_VSYNC_wire\
        );

    \ADV_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18842\,
            PADOUT => \N__18841\,
            PADIN => \N__18840\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14452\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18833\,
            DIN => \N__18832\,
            DOUT => \N__18831\,
            PACKAGEPIN => \ADV_R_wire\(3)
        );

    \ADV_R_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18833\,
            PADOUT => \N__18832\,
            PADIN => \N__18831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10196\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18824\,
            DIN => \N__18823\,
            DOUT => \N__18822\,
            PACKAGEPIN => \ADV_B_wire\(5)
        );

    \ADV_B_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18824\,
            PADOUT => \N__18823\,
            PADIN => \N__18822\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10310\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18815\,
            DIN => \N__18814\,
            DOUT => \N__18813\,
            PACKAGEPIN => DEBUG(7)
        );

    \DEBUG_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18815\,
            PADOUT => \N__18814\,
            PADIN => \N__18813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11851\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18806\,
            DIN => \N__18805\,
            DOUT => \N__18804\,
            PACKAGEPIN => \TVP_VIDEO_wire\(6)
        );

    \TVP_VIDEO_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18806\,
            PADOUT => \N__18805\,
            PADIN => \N__18804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18797\,
            DIN => \N__18796\,
            DOUT => \N__18795\,
            PACKAGEPIN => \ADV_G_wire\(1)
        );

    \ADV_G_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18797\,
            PADOUT => \N__18796\,
            PADIN => \N__18795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10264\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18788\,
            DIN => \N__18787\,
            DOUT => \N__18786\,
            PACKAGEPIN => \ADV_R_wire\(0)
        );

    \ADV_R_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18788\,
            PADOUT => \N__18787\,
            PADIN => \N__18786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8498\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18779\,
            DIN => \N__18778\,
            DOUT => \N__18777\,
            PACKAGEPIN => DEBUG(2)
        );

    \DEBUG_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18779\,
            PADOUT => \N__18778\,
            PADIN => \N__18777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9112\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18770\,
            DIN => \N__18769\,
            DOUT => \N__18768\,
            PACKAGEPIN => \TVP_VIDEO_wire\(3)
        );

    \TVP_VIDEO_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18770\,
            PADOUT => \N__18769\,
            PADIN => \N__18768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18761\,
            DIN => \N__18760\,
            DOUT => \N__18759\,
            PACKAGEPIN => \ADV_G_wire\(4)
        );

    \ADV_G_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18761\,
            PADOUT => \N__18760\,
            PADIN => \N__18759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10138\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18752\,
            DIN => \N__18751\,
            DOUT => \N__18750\,
            PACKAGEPIN => \ADV_R_wire\(5)
        );

    \ADV_R_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18752\,
            PADOUT => \N__18751\,
            PADIN => \N__18750\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10318\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18743\,
            DIN => \N__18742\,
            DOUT => \N__18741\,
            PACKAGEPIN => \TVP_VIDEO_wire\(9)
        );

    \TVP_VIDEO_pad_9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18743\,
            PADOUT => \N__18742\,
            PADIN => \N__18741\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18734\,
            DIN => \N__18733\,
            DOUT => \N__18732\,
            PACKAGEPIN => \ADV_G_wire\(3)
        );

    \ADV_G_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18734\,
            PADOUT => \N__18733\,
            PADIN => \N__18732\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10198\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18725\,
            DIN => \N__18724\,
            DOUT => \N__18723\,
            PACKAGEPIN => \ADV_HSYNC_wire\
        );

    \ADV_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18725\,
            PADOUT => \N__18724\,
            PADIN => \N__18723\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7309\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18716\,
            DIN => \N__18715\,
            DOUT => \N__18714\,
            PACKAGEPIN => \ADV_R_wire\(2)
        );

    \ADV_R_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18716\,
            PADOUT => \N__18715\,
            PADIN => \N__18714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8429\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18707\,
            DIN => \N__18706\,
            DOUT => \N__18705\,
            PACKAGEPIN => DEBUG(1)
        );

    \DEBUG_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18707\,
            PADOUT => \N__18706\,
            PADIN => \N__18705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12100\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18698\,
            DIN => \N__18697\,
            DOUT => \N__18696\,
            PACKAGEPIN => \ADV_B_wire\(4)
        );

    \ADV_B_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18698\,
            PADOUT => \N__18697\,
            PADIN => \N__18696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10137\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18689\,
            DIN => \N__18688\,
            DOUT => \N__18687\,
            PACKAGEPIN => DEBUG(4)
        );

    \DEBUG_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18689\,
            PADOUT => \N__18688\,
            PADIN => \N__18687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9370\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18680\,
            DIN => \N__18679\,
            DOUT => \N__18678\,
            PACKAGEPIN => \ADV_B_wire\(1)
        );

    \ADV_B_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18680\,
            PADOUT => \N__18679\,
            PADIN => \N__18678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10256\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18671\,
            DIN => \N__18670\,
            DOUT => \N__18669\,
            PACKAGEPIN => \ADV_G_wire\(6)
        );

    \ADV_G_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18671\,
            PADOUT => \N__18670\,
            PADIN => \N__18669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10077\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_SYNC_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18662\,
            DIN => \N__18661\,
            DOUT => \N__18660\,
            PACKAGEPIN => \ADV_SYNC_N_wire\
        );

    \ADV_SYNC_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18662\,
            PADOUT => \N__18661\,
            PADIN => \N__18660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18653\,
            DIN => \N__18652\,
            DOUT => \N__18651\,
            PACKAGEPIN => \ADV_R_wire\(7)
        );

    \ADV_R_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18653\,
            PADOUT => \N__18652\,
            PADIN => \N__18651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10020\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18644\,
            DIN => \N__18643\,
            DOUT => \N__18642\,
            PACKAGEPIN => \ADV_B_wire\(6)
        );

    \ADV_B_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18644\,
            PADOUT => \N__18643\,
            PADIN => \N__18642\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18635\,
            DIN => \N__18634\,
            DOUT => \N__18633\,
            PACKAGEPIN => DEBUG(6)
        );

    \DEBUG_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18635\,
            PADOUT => \N__18634\,
            PADIN => \N__18633\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9934\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18626\,
            DIN => \N__18625\,
            DOUT => \N__18624\,
            PACKAGEPIN => \TVP_VIDEO_wire\(7)
        );

    \TVP_VIDEO_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18626\,
            PADOUT => \N__18625\,
            PADIN => \N__18624\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18617\,
            DIN => \N__18616\,
            DOUT => \N__18615\,
            PACKAGEPIN => \ADV_G_wire\(0)
        );

    \ADV_G_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18617\,
            PADOUT => \N__18616\,
            PADIN => \N__18615\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8509\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18608\,
            DIN => \N__18607\,
            DOUT => \N__18606\,
            PACKAGEPIN => \ADV_R_wire\(1)
        );

    \ADV_R_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18608\,
            PADOUT => \N__18607\,
            PADIN => \N__18606\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10257\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18599\,
            DIN => \N__18598\,
            DOUT => \N__18597\,
            PACKAGEPIN => DEBUG(5)
        );

    \DEBUG_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18599\,
            PADOUT => \N__18598\,
            PADIN => \N__18597\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9643\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18590\,
            DIN => \N__18589\,
            DOUT => \N__18588\,
            PACKAGEPIN => \TVP_HSYNC_wire\
        );

    \TVP_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18590\,
            PADOUT => \N__18589\,
            PADIN => \N__18588\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_HSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18581\,
            DIN => \N__18580\,
            DOUT => \N__18579\,
            PACKAGEPIN => \ADV_G_wire\(7)
        );

    \ADV_G_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18581\,
            PADOUT => \N__18580\,
            PADIN => \N__18579\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10019\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18572\,
            DIN => \N__18571\,
            DOUT => \N__18570\,
            PACKAGEPIN => \ADV_R_wire\(6)
        );

    \ADV_R_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18572\,
            PADOUT => \N__18571\,
            PADIN => \N__18570\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10081\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18563\,
            DIN => \N__18562\,
            DOUT => \N__18561\,
            PACKAGEPIN => \TVP_VSYNC_wire\
        );

    \TVP_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18563\,
            PADOUT => \N__18562\,
            PADIN => \N__18561\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_BLANK_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18554\,
            DIN => \N__18553\,
            DOUT => \N__18552\,
            PACKAGEPIN => \ADV_BLANK_N_wire\
        );

    \ADV_BLANK_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18554\,
            PADOUT => \N__18553\,
            PADIN => \N__18552\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12537\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18545\,
            DIN => \N__18544\,
            DOUT => \N__18543\,
            PACKAGEPIN => DEBUG(0)
        );

    \DEBUG_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18545\,
            PADOUT => \N__18544\,
            PADIN => \N__18543\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18536\,
            DIN => \N__18535\,
            DOUT => \N__18534\,
            PACKAGEPIN => \ADV_B_wire\(2)
        );

    \ADV_B_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18536\,
            PADOUT => \N__18535\,
            PADIN => \N__18534\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8440\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18527\,
            DIN => \N__18526\,
            DOUT => \N__18525\,
            PACKAGEPIN => \ADV_B_wire\(7)
        );

    \ADV_B_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18527\,
            PADOUT => \N__18526\,
            PADIN => \N__18525\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10021\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18518\,
            DIN => \N__18517\,
            DOUT => \N__18516\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18518\,
            PADOUT => \N__18517\,
            PADIN => \N__18516\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8803\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__18509\,
            DIN => \N__18508\,
            DOUT => \N__18507\,
            PACKAGEPIN => \TVP_VIDEO_wire\(4)
        );

    \TVP_VIDEO_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18509\,
            PADOUT => \N__18508\,
            PADIN => \N__18507\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__4528\ : InMux
    port map (
            O => \N__18490\,
            I => \N__18484\
        );

    \I__4527\ : InMux
    port map (
            O => \N__18489\,
            I => \N__18481\
        );

    \I__4526\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18478\
        );

    \I__4525\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18466\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__18484\,
            I => \N__18461\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__18481\,
            I => \N__18461\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__18478\,
            I => \N__18458\
        );

    \I__4521\ : InMux
    port map (
            O => \N__18477\,
            I => \N__18455\
        );

    \I__4520\ : InMux
    port map (
            O => \N__18476\,
            I => \N__18452\
        );

    \I__4519\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18445\
        );

    \I__4518\ : InMux
    port map (
            O => \N__18474\,
            I => \N__18442\
        );

    \I__4517\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18436\
        );

    \I__4516\ : InMux
    port map (
            O => \N__18472\,
            I => \N__18433\
        );

    \I__4515\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18430\
        );

    \I__4514\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18427\
        );

    \I__4513\ : InMux
    port map (
            O => \N__18469\,
            I => \N__18424\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__18466\,
            I => \N__18421\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__18461\,
            I => \N__18412\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__18458\,
            I => \N__18412\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__18455\,
            I => \N__18412\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__18452\,
            I => \N__18412\
        );

    \I__4507\ : InMux
    port map (
            O => \N__18451\,
            I => \N__18409\
        );

    \I__4506\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18406\
        );

    \I__4505\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18403\
        );

    \I__4504\ : InMux
    port map (
            O => \N__18448\,
            I => \N__18400\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__18445\,
            I => \N__18397\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__18442\,
            I => \N__18394\
        );

    \I__4501\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18390\
        );

    \I__4500\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18387\
        );

    \I__4499\ : InMux
    port map (
            O => \N__18439\,
            I => \N__18382\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__18436\,
            I => \N__18379\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__18433\,
            I => \N__18376\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__18430\,
            I => \N__18373\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__18427\,
            I => \N__18368\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18368\
        );

    \I__4493\ : Span4Mux_h
    port map (
            O => \N__18421\,
            I => \N__18363\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__18412\,
            I => \N__18363\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__18409\,
            I => \N__18360\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__18406\,
            I => \N__18351\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__18403\,
            I => \N__18351\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__18400\,
            I => \N__18351\
        );

    \I__4487\ : Span4Mux_v
    port map (
            O => \N__18397\,
            I => \N__18351\
        );

    \I__4486\ : Span4Mux_v
    port map (
            O => \N__18394\,
            I => \N__18348\
        );

    \I__4485\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18345\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__18390\,
            I => \N__18342\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__18387\,
            I => \N__18339\
        );

    \I__4482\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18336\
        );

    \I__4481\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18333\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__18382\,
            I => \N__18330\
        );

    \I__4479\ : Span12Mux_v
    port map (
            O => \N__18379\,
            I => \N__18327\
        );

    \I__4478\ : Span12Mux_h
    port map (
            O => \N__18376\,
            I => \N__18322\
        );

    \I__4477\ : Span12Mux_h
    port map (
            O => \N__18373\,
            I => \N__18322\
        );

    \I__4476\ : Span4Mux_h
    port map (
            O => \N__18368\,
            I => \N__18317\
        );

    \I__4475\ : Span4Mux_v
    port map (
            O => \N__18363\,
            I => \N__18317\
        );

    \I__4474\ : Span4Mux_v
    port map (
            O => \N__18360\,
            I => \N__18310\
        );

    \I__4473\ : Span4Mux_v
    port map (
            O => \N__18351\,
            I => \N__18310\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__18348\,
            I => \N__18310\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__18345\,
            I => \N__18303\
        );

    \I__4470\ : Span4Mux_v
    port map (
            O => \N__18342\,
            I => \N__18303\
        );

    \I__4469\ : Span4Mux_v
    port map (
            O => \N__18339\,
            I => \N__18303\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__18336\,
            I => \TX_ADDR_11\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__18333\,
            I => \TX_ADDR_11\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__18330\,
            I => \TX_ADDR_11\
        );

    \I__4465\ : Odrv12
    port map (
            O => \N__18327\,
            I => \TX_ADDR_11\
        );

    \I__4464\ : Odrv12
    port map (
            O => \N__18322\,
            I => \TX_ADDR_11\
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__18317\,
            I => \TX_ADDR_11\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__18310\,
            I => \TX_ADDR_11\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__18303\,
            I => \TX_ADDR_11\
        );

    \I__4460\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18283\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__18283\,
            I => \N__18280\
        );

    \I__4458\ : Span4Mux_v
    port map (
            O => \N__18280\,
            I => \N__18277\
        );

    \I__4457\ : Sp12to4
    port map (
            O => \N__18277\,
            I => \N__18274\
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__18274\,
            I => \line_buffer.n756\
        );

    \I__4455\ : InMux
    port map (
            O => \N__18271\,
            I => \N__18268\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__18268\,
            I => \N__18265\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__18265\,
            I => \N__18262\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__18262\,
            I => \N__18259\
        );

    \I__4451\ : Span4Mux_v
    port map (
            O => \N__18259\,
            I => \N__18256\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__18256\,
            I => \N__18253\
        );

    \I__4449\ : Odrv4
    port map (
            O => \N__18253\,
            I => \line_buffer.n748\
        );

    \I__4448\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18247\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__18247\,
            I => \line_buffer.n3025\
        );

    \I__4446\ : SRMux
    port map (
            O => \N__18244\,
            I => \N__18240\
        );

    \I__4445\ : SRMux
    port map (
            O => \N__18243\,
            I => \N__18237\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__18240\,
            I => \N__18232\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__18237\,
            I => \N__18229\
        );

    \I__4442\ : SRMux
    port map (
            O => \N__18236\,
            I => \N__18226\
        );

    \I__4441\ : SRMux
    port map (
            O => \N__18235\,
            I => \N__18223\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__18232\,
            I => \N__18220\
        );

    \I__4439\ : Span4Mux_v
    port map (
            O => \N__18229\,
            I => \N__18213\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__18226\,
            I => \N__18213\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__18223\,
            I => \N__18213\
        );

    \I__4436\ : Span4Mux_v
    port map (
            O => \N__18220\,
            I => \N__18210\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__18213\,
            I => \N__18207\
        );

    \I__4434\ : Span4Mux_v
    port map (
            O => \N__18210\,
            I => \N__18202\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__18207\,
            I => \N__18202\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__18202\,
            I => \line_buffer.n729\
        );

    \I__4431\ : SRMux
    port map (
            O => \N__18199\,
            I => \N__18196\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__18196\,
            I => \N__18193\
        );

    \I__4429\ : Span4Mux_s3_v
    port map (
            O => \N__18193\,
            I => \N__18188\
        );

    \I__4428\ : SRMux
    port map (
            O => \N__18192\,
            I => \N__18185\
        );

    \I__4427\ : SRMux
    port map (
            O => \N__18191\,
            I => \N__18181\
        );

    \I__4426\ : Span4Mux_v
    port map (
            O => \N__18188\,
            I => \N__18176\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__18185\,
            I => \N__18176\
        );

    \I__4424\ : SRMux
    port map (
            O => \N__18184\,
            I => \N__18173\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__18181\,
            I => \N__18170\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__18176\,
            I => \N__18167\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__18173\,
            I => \N__18164\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__18170\,
            I => \N__18161\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__18167\,
            I => \N__18156\
        );

    \I__4418\ : Span4Mux_h
    port map (
            O => \N__18164\,
            I => \N__18156\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__18161\,
            I => \line_buffer.n697\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__18156\,
            I => \line_buffer.n697\
        );

    \I__4415\ : InMux
    port map (
            O => \N__18151\,
            I => \N__18146\
        );

    \I__4414\ : InMux
    port map (
            O => \N__18150\,
            I => \N__18143\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__18149\,
            I => \N__18140\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__18146\,
            I => \N__18130\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__18143\,
            I => \N__18130\
        );

    \I__4410\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18125\
        );

    \I__4409\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18125\
        );

    \I__4408\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18122\
        );

    \I__4407\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18119\
        );

    \I__4406\ : InMux
    port map (
            O => \N__18136\,
            I => \N__18116\
        );

    \I__4405\ : InMux
    port map (
            O => \N__18135\,
            I => \N__18113\
        );

    \I__4404\ : Span4Mux_v
    port map (
            O => \N__18130\,
            I => \N__18108\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__18125\,
            I => \N__18108\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__18122\,
            I => \N__18104\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__18119\,
            I => \N__18101\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__18116\,
            I => \N__18098\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__18113\,
            I => \N__18095\
        );

    \I__4398\ : Sp12to4
    port map (
            O => \N__18108\,
            I => \N__18092\
        );

    \I__4397\ : InMux
    port map (
            O => \N__18107\,
            I => \N__18089\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__18104\,
            I => \N__18084\
        );

    \I__4395\ : Span4Mux_v
    port map (
            O => \N__18101\,
            I => \N__18084\
        );

    \I__4394\ : Span12Mux_v
    port map (
            O => \N__18098\,
            I => \N__18077\
        );

    \I__4393\ : Span12Mux_v
    port map (
            O => \N__18095\,
            I => \N__18077\
        );

    \I__4392\ : Span12Mux_v
    port map (
            O => \N__18092\,
            I => \N__18077\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__18089\,
            I => \RX_ADDR_12\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__18084\,
            I => \RX_ADDR_12\
        );

    \I__4389\ : Odrv12
    port map (
            O => \N__18077\,
            I => \RX_ADDR_12\
        );

    \I__4388\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18064\
        );

    \I__4387\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18059\
        );

    \I__4386\ : InMux
    port map (
            O => \N__18068\,
            I => \N__18059\
        );

    \I__4385\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18056\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__18064\,
            I => \N__18051\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__18059\,
            I => \N__18048\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__18056\,
            I => \N__18043\
        );

    \I__4381\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18040\
        );

    \I__4380\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18037\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__18051\,
            I => \N__18032\
        );

    \I__4378\ : Span4Mux_v
    port map (
            O => \N__18048\,
            I => \N__18032\
        );

    \I__4377\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18029\
        );

    \I__4376\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18026\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__18043\,
            I => \N__18023\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__18040\,
            I => \N__18020\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__18037\,
            I => \N__18017\
        );

    \I__4372\ : Span4Mux_h
    port map (
            O => \N__18032\,
            I => \N__18014\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__18029\,
            I => \N__18011\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__18026\,
            I => \N__18008\
        );

    \I__4369\ : Span4Mux_h
    port map (
            O => \N__18023\,
            I => \N__18004\
        );

    \I__4368\ : Span4Mux_v
    port map (
            O => \N__18020\,
            I => \N__17999\
        );

    \I__4367\ : Span4Mux_v
    port map (
            O => \N__18017\,
            I => \N__17999\
        );

    \I__4366\ : Span4Mux_h
    port map (
            O => \N__18014\,
            I => \N__17992\
        );

    \I__4365\ : Span4Mux_v
    port map (
            O => \N__18011\,
            I => \N__17992\
        );

    \I__4364\ : Span4Mux_v
    port map (
            O => \N__18008\,
            I => \N__17992\
        );

    \I__4363\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17989\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__18004\,
            I => \RX_ADDR_11\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__17999\,
            I => \RX_ADDR_11\
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__17992\,
            I => \RX_ADDR_11\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__17989\,
            I => \RX_ADDR_11\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__17980\,
            I => \N__17976\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__17979\,
            I => \N__17968\
        );

    \I__4356\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17965\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__17975\,
            I => \N__17962\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__17974\,
            I => \N__17959\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__17973\,
            I => \N__17956\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__17972\,
            I => \N__17953\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__17971\,
            I => \N__17949\
        );

    \I__4350\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17946\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__17965\,
            I => \N__17943\
        );

    \I__4348\ : InMux
    port map (
            O => \N__17962\,
            I => \N__17940\
        );

    \I__4347\ : InMux
    port map (
            O => \N__17959\,
            I => \N__17937\
        );

    \I__4346\ : InMux
    port map (
            O => \N__17956\,
            I => \N__17934\
        );

    \I__4345\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17931\
        );

    \I__4344\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17926\
        );

    \I__4343\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17926\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__17946\,
            I => \N__17922\
        );

    \I__4341\ : Span4Mux_h
    port map (
            O => \N__17943\,
            I => \N__17919\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__17940\,
            I => \N__17916\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__17937\,
            I => \N__17911\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__17934\,
            I => \N__17911\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__17931\,
            I => \N__17908\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__17926\,
            I => \N__17905\
        );

    \I__4335\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17902\
        );

    \I__4334\ : Span4Mux_v
    port map (
            O => \N__17922\,
            I => \N__17897\
        );

    \I__4333\ : Span4Mux_h
    port map (
            O => \N__17919\,
            I => \N__17897\
        );

    \I__4332\ : Span4Mux_h
    port map (
            O => \N__17916\,
            I => \N__17892\
        );

    \I__4331\ : Span4Mux_h
    port map (
            O => \N__17911\,
            I => \N__17892\
        );

    \I__4330\ : Span12Mux_v
    port map (
            O => \N__17908\,
            I => \N__17887\
        );

    \I__4329\ : Span12Mux_v
    port map (
            O => \N__17905\,
            I => \N__17887\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__17902\,
            I => \RX_ADDR_13\
        );

    \I__4327\ : Odrv4
    port map (
            O => \N__17897\,
            I => \RX_ADDR_13\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__17892\,
            I => \RX_ADDR_13\
        );

    \I__4325\ : Odrv12
    port map (
            O => \N__17887\,
            I => \RX_ADDR_13\
        );

    \I__4324\ : InMux
    port map (
            O => \N__17878\,
            I => \N__17862\
        );

    \I__4323\ : InMux
    port map (
            O => \N__17877\,
            I => \N__17858\
        );

    \I__4322\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17854\
        );

    \I__4321\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17851\
        );

    \I__4320\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17846\
        );

    \I__4319\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17846\
        );

    \I__4318\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17839\
        );

    \I__4317\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17839\
        );

    \I__4316\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17839\
        );

    \I__4315\ : InMux
    port map (
            O => \N__17869\,
            I => \N__17828\
        );

    \I__4314\ : InMux
    port map (
            O => \N__17868\,
            I => \N__17828\
        );

    \I__4313\ : InMux
    port map (
            O => \N__17867\,
            I => \N__17828\
        );

    \I__4312\ : InMux
    port map (
            O => \N__17866\,
            I => \N__17828\
        );

    \I__4311\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17828\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__17862\,
            I => \N__17825\
        );

    \I__4309\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17822\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__17858\,
            I => \N__17819\
        );

    \I__4307\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17816\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__17854\,
            I => \N__17813\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__17851\,
            I => \N__17806\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__17846\,
            I => \N__17806\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__17839\,
            I => \N__17803\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17796\
        );

    \I__4301\ : Span4Mux_v
    port map (
            O => \N__17825\,
            I => \N__17796\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17796\
        );

    \I__4299\ : Span4Mux_h
    port map (
            O => \N__17819\,
            I => \N__17789\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17789\
        );

    \I__4297\ : Span4Mux_v
    port map (
            O => \N__17813\,
            I => \N__17789\
        );

    \I__4296\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17784\
        );

    \I__4295\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17784\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__17806\,
            I => \N__17781\
        );

    \I__4293\ : Span4Mux_v
    port map (
            O => \N__17803\,
            I => \N__17777\
        );

    \I__4292\ : Span4Mux_v
    port map (
            O => \N__17796\,
            I => \N__17772\
        );

    \I__4291\ : Span4Mux_h
    port map (
            O => \N__17789\,
            I => \N__17772\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__17784\,
            I => \N__17769\
        );

    \I__4289\ : Span4Mux_h
    port map (
            O => \N__17781\,
            I => \N__17766\
        );

    \I__4288\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17763\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__17777\,
            I => \N__17759\
        );

    \I__4286\ : Span4Mux_h
    port map (
            O => \N__17772\,
            I => \N__17754\
        );

    \I__4285\ : Span4Mux_v
    port map (
            O => \N__17769\,
            I => \N__17754\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__17766\,
            I => \N__17749\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__17763\,
            I => \N__17749\
        );

    \I__4282\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17746\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__17759\,
            I => n25
        );

    \I__4280\ : Odrv4
    port map (
            O => \N__17754\,
            I => n25
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__17749\,
            I => n25
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__17746\,
            I => n25
        );

    \I__4277\ : SRMux
    port map (
            O => \N__17737\,
            I => \N__17733\
        );

    \I__4276\ : SRMux
    port map (
            O => \N__17736\,
            I => \N__17730\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__17733\,
            I => \N__17726\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__17730\,
            I => \N__17723\
        );

    \I__4273\ : SRMux
    port map (
            O => \N__17729\,
            I => \N__17720\
        );

    \I__4272\ : Span4Mux_v
    port map (
            O => \N__17726\,
            I => \N__17713\
        );

    \I__4271\ : Span4Mux_h
    port map (
            O => \N__17723\,
            I => \N__17713\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__17720\,
            I => \N__17713\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__17713\,
            I => \N__17709\
        );

    \I__4268\ : SRMux
    port map (
            O => \N__17712\,
            I => \N__17706\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__17709\,
            I => \N__17701\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__17706\,
            I => \N__17701\
        );

    \I__4265\ : Span4Mux_h
    port map (
            O => \N__17701\,
            I => \N__17698\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__17698\,
            I => \line_buffer.n633\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__17695\,
            I => \N__17690\
        );

    \I__4262\ : InMux
    port map (
            O => \N__17694\,
            I => \N__17687\
        );

    \I__4261\ : InMux
    port map (
            O => \N__17693\,
            I => \N__17679\
        );

    \I__4260\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17679\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17676\
        );

    \I__4258\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17673\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__17685\,
            I => \N__17669\
        );

    \I__4256\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17665\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__17679\,
            I => \N__17662\
        );

    \I__4254\ : Span4Mux_v
    port map (
            O => \N__17676\,
            I => \N__17657\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__17673\,
            I => \N__17657\
        );

    \I__4252\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17652\
        );

    \I__4251\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17652\
        );

    \I__4250\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17646\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__17665\,
            I => \N__17641\
        );

    \I__4248\ : Span4Mux_v
    port map (
            O => \N__17662\,
            I => \N__17641\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__17657\,
            I => \N__17636\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__17652\,
            I => \N__17636\
        );

    \I__4245\ : InMux
    port map (
            O => \N__17651\,
            I => \N__17632\
        );

    \I__4244\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17629\
        );

    \I__4243\ : InMux
    port map (
            O => \N__17649\,
            I => \N__17626\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__17646\,
            I => \N__17621\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__17641\,
            I => \N__17621\
        );

    \I__4240\ : Span4Mux_h
    port map (
            O => \N__17636\,
            I => \N__17618\
        );

    \I__4239\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17615\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__17632\,
            I => \TX_ADDR_13\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__17629\,
            I => \TX_ADDR_13\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__17626\,
            I => \TX_ADDR_13\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__17621\,
            I => \TX_ADDR_13\
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__17618\,
            I => \TX_ADDR_13\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__17615\,
            I => \TX_ADDR_13\
        );

    \I__4232\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17599\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__17599\,
            I => \N__17596\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__17596\,
            I => \N__17593\
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__17593\,
            I => \TX_DATA_4\
        );

    \I__4228\ : ClkMux
    port map (
            O => \N__17590\,
            I => \N__17584\
        );

    \I__4227\ : ClkMux
    port map (
            O => \N__17589\,
            I => \N__17581\
        );

    \I__4226\ : ClkMux
    port map (
            O => \N__17588\,
            I => \N__17576\
        );

    \I__4225\ : ClkMux
    port map (
            O => \N__17587\,
            I => \N__17573\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__17584\,
            I => \N__17569\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__17581\,
            I => \N__17566\
        );

    \I__4222\ : ClkMux
    port map (
            O => \N__17580\,
            I => \N__17563\
        );

    \I__4221\ : ClkMux
    port map (
            O => \N__17579\,
            I => \N__17560\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__17576\,
            I => \N__17555\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__17573\,
            I => \N__17552\
        );

    \I__4218\ : ClkMux
    port map (
            O => \N__17572\,
            I => \N__17549\
        );

    \I__4217\ : Span4Mux_s2_v
    port map (
            O => \N__17569\,
            I => \N__17541\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__17566\,
            I => \N__17541\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__17563\,
            I => \N__17541\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__17560\,
            I => \N__17538\
        );

    \I__4213\ : ClkMux
    port map (
            O => \N__17559\,
            I => \N__17535\
        );

    \I__4212\ : ClkMux
    port map (
            O => \N__17558\,
            I => \N__17532\
        );

    \I__4211\ : Span4Mux_s2_v
    port map (
            O => \N__17555\,
            I => \N__17522\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__17552\,
            I => \N__17522\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17522\
        );

    \I__4208\ : ClkMux
    port map (
            O => \N__17548\,
            I => \N__17519\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__17541\,
            I => \N__17509\
        );

    \I__4206\ : Span4Mux_h
    port map (
            O => \N__17538\,
            I => \N__17509\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__17535\,
            I => \N__17509\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__17532\,
            I => \N__17506\
        );

    \I__4203\ : ClkMux
    port map (
            O => \N__17531\,
            I => \N__17503\
        );

    \I__4202\ : ClkMux
    port map (
            O => \N__17530\,
            I => \N__17500\
        );

    \I__4201\ : ClkMux
    port map (
            O => \N__17529\,
            I => \N__17492\
        );

    \I__4200\ : Span4Mux_v
    port map (
            O => \N__17522\,
            I => \N__17485\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__17519\,
            I => \N__17485\
        );

    \I__4198\ : ClkMux
    port map (
            O => \N__17518\,
            I => \N__17482\
        );

    \I__4197\ : ClkMux
    port map (
            O => \N__17517\,
            I => \N__17478\
        );

    \I__4196\ : ClkMux
    port map (
            O => \N__17516\,
            I => \N__17475\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__17509\,
            I => \N__17467\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__17506\,
            I => \N__17467\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__17503\,
            I => \N__17467\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__17500\,
            I => \N__17464\
        );

    \I__4191\ : ClkMux
    port map (
            O => \N__17499\,
            I => \N__17461\
        );

    \I__4190\ : ClkMux
    port map (
            O => \N__17498\,
            I => \N__17458\
        );

    \I__4189\ : ClkMux
    port map (
            O => \N__17497\,
            I => \N__17454\
        );

    \I__4188\ : ClkMux
    port map (
            O => \N__17496\,
            I => \N__17450\
        );

    \I__4187\ : ClkMux
    port map (
            O => \N__17495\,
            I => \N__17447\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__17492\,
            I => \N__17443\
        );

    \I__4185\ : ClkMux
    port map (
            O => \N__17491\,
            I => \N__17440\
        );

    \I__4184\ : ClkMux
    port map (
            O => \N__17490\,
            I => \N__17437\
        );

    \I__4183\ : Span4Mux_v
    port map (
            O => \N__17485\,
            I => \N__17429\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__17482\,
            I => \N__17429\
        );

    \I__4181\ : ClkMux
    port map (
            O => \N__17481\,
            I => \N__17426\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__17478\,
            I => \N__17420\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__17475\,
            I => \N__17416\
        );

    \I__4178\ : ClkMux
    port map (
            O => \N__17474\,
            I => \N__17413\
        );

    \I__4177\ : Span4Mux_v
    port map (
            O => \N__17467\,
            I => \N__17404\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__17464\,
            I => \N__17404\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__17461\,
            I => \N__17404\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__17458\,
            I => \N__17401\
        );

    \I__4173\ : ClkMux
    port map (
            O => \N__17457\,
            I => \N__17398\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__17454\,
            I => \N__17393\
        );

    \I__4171\ : ClkMux
    port map (
            O => \N__17453\,
            I => \N__17390\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__17450\,
            I => \N__17385\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17385\
        );

    \I__4168\ : ClkMux
    port map (
            O => \N__17446\,
            I => \N__17382\
        );

    \I__4167\ : Span4Mux_h
    port map (
            O => \N__17443\,
            I => \N__17375\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__17440\,
            I => \N__17375\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__17437\,
            I => \N__17375\
        );

    \I__4164\ : ClkMux
    port map (
            O => \N__17436\,
            I => \N__17372\
        );

    \I__4163\ : ClkMux
    port map (
            O => \N__17435\,
            I => \N__17369\
        );

    \I__4162\ : ClkMux
    port map (
            O => \N__17434\,
            I => \N__17366\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__17429\,
            I => \N__17361\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__17426\,
            I => \N__17361\
        );

    \I__4159\ : ClkMux
    port map (
            O => \N__17425\,
            I => \N__17358\
        );

    \I__4158\ : ClkMux
    port map (
            O => \N__17424\,
            I => \N__17355\
        );

    \I__4157\ : ClkMux
    port map (
            O => \N__17423\,
            I => \N__17352\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__17420\,
            I => \N__17349\
        );

    \I__4155\ : ClkMux
    port map (
            O => \N__17419\,
            I => \N__17346\
        );

    \I__4154\ : Span4Mux_v
    port map (
            O => \N__17416\,
            I => \N__17341\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__17413\,
            I => \N__17341\
        );

    \I__4152\ : ClkMux
    port map (
            O => \N__17412\,
            I => \N__17338\
        );

    \I__4151\ : ClkMux
    port map (
            O => \N__17411\,
            I => \N__17334\
        );

    \I__4150\ : Span4Mux_v
    port map (
            O => \N__17404\,
            I => \N__17320\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__17401\,
            I => \N__17320\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__17398\,
            I => \N__17320\
        );

    \I__4147\ : ClkMux
    port map (
            O => \N__17397\,
            I => \N__17317\
        );

    \I__4146\ : ClkMux
    port map (
            O => \N__17396\,
            I => \N__17314\
        );

    \I__4145\ : Span4Mux_v
    port map (
            O => \N__17393\,
            I => \N__17306\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__17390\,
            I => \N__17306\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__17385\,
            I => \N__17301\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__17382\,
            I => \N__17301\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__17375\,
            I => \N__17292\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__17372\,
            I => \N__17292\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__17369\,
            I => \N__17292\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__17366\,
            I => \N__17292\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__17361\,
            I => \N__17287\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__17358\,
            I => \N__17287\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__17355\,
            I => \N__17282\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__17352\,
            I => \N__17282\
        );

    \I__4133\ : Span4Mux_h
    port map (
            O => \N__17349\,
            I => \N__17277\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__17346\,
            I => \N__17277\
        );

    \I__4131\ : Span4Mux_v
    port map (
            O => \N__17341\,
            I => \N__17272\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__17338\,
            I => \N__17272\
        );

    \I__4129\ : ClkMux
    port map (
            O => \N__17337\,
            I => \N__17269\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__17334\,
            I => \N__17265\
        );

    \I__4127\ : ClkMux
    port map (
            O => \N__17333\,
            I => \N__17262\
        );

    \I__4126\ : ClkMux
    port map (
            O => \N__17332\,
            I => \N__17259\
        );

    \I__4125\ : ClkMux
    port map (
            O => \N__17331\,
            I => \N__17256\
        );

    \I__4124\ : ClkMux
    port map (
            O => \N__17330\,
            I => \N__17253\
        );

    \I__4123\ : ClkMux
    port map (
            O => \N__17329\,
            I => \N__17250\
        );

    \I__4122\ : ClkMux
    port map (
            O => \N__17328\,
            I => \N__17246\
        );

    \I__4121\ : ClkMux
    port map (
            O => \N__17327\,
            I => \N__17242\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__17320\,
            I => \N__17236\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__17317\,
            I => \N__17236\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__17314\,
            I => \N__17233\
        );

    \I__4117\ : ClkMux
    port map (
            O => \N__17313\,
            I => \N__17230\
        );

    \I__4116\ : IoInMux
    port map (
            O => \N__17312\,
            I => \N__17227\
        );

    \I__4115\ : ClkMux
    port map (
            O => \N__17311\,
            I => \N__17222\
        );

    \I__4114\ : Span4Mux_v
    port map (
            O => \N__17306\,
            I => \N__17219\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__17301\,
            I => \N__17214\
        );

    \I__4112\ : Span4Mux_v
    port map (
            O => \N__17292\,
            I => \N__17214\
        );

    \I__4111\ : Span4Mux_v
    port map (
            O => \N__17287\,
            I => \N__17210\
        );

    \I__4110\ : Span4Mux_v
    port map (
            O => \N__17282\,
            I => \N__17207\
        );

    \I__4109\ : Span4Mux_v
    port map (
            O => \N__17277\,
            I => \N__17200\
        );

    \I__4108\ : Span4Mux_h
    port map (
            O => \N__17272\,
            I => \N__17200\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__17269\,
            I => \N__17200\
        );

    \I__4106\ : ClkMux
    port map (
            O => \N__17268\,
            I => \N__17197\
        );

    \I__4105\ : Span4Mux_v
    port map (
            O => \N__17265\,
            I => \N__17190\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__17262\,
            I => \N__17190\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__17259\,
            I => \N__17187\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__17256\,
            I => \N__17180\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__17253\,
            I => \N__17180\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__17250\,
            I => \N__17180\
        );

    \I__4099\ : ClkMux
    port map (
            O => \N__17249\,
            I => \N__17177\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__17246\,
            I => \N__17174\
        );

    \I__4097\ : ClkMux
    port map (
            O => \N__17245\,
            I => \N__17171\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__17242\,
            I => \N__17168\
        );

    \I__4095\ : ClkMux
    port map (
            O => \N__17241\,
            I => \N__17165\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__17236\,
            I => \N__17158\
        );

    \I__4093\ : Span4Mux_h
    port map (
            O => \N__17233\,
            I => \N__17158\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__17230\,
            I => \N__17158\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__17227\,
            I => \N__17155\
        );

    \I__4090\ : ClkMux
    port map (
            O => \N__17226\,
            I => \N__17152\
        );

    \I__4089\ : ClkMux
    port map (
            O => \N__17225\,
            I => \N__17148\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__17222\,
            I => \N__17145\
        );

    \I__4087\ : Span4Mux_v
    port map (
            O => \N__17219\,
            I => \N__17140\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__17214\,
            I => \N__17140\
        );

    \I__4085\ : ClkMux
    port map (
            O => \N__17213\,
            I => \N__17137\
        );

    \I__4084\ : Span4Mux_h
    port map (
            O => \N__17210\,
            I => \N__17130\
        );

    \I__4083\ : Span4Mux_v
    port map (
            O => \N__17207\,
            I => \N__17130\
        );

    \I__4082\ : Span4Mux_v
    port map (
            O => \N__17200\,
            I => \N__17130\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__17197\,
            I => \N__17127\
        );

    \I__4080\ : ClkMux
    port map (
            O => \N__17196\,
            I => \N__17124\
        );

    \I__4079\ : ClkMux
    port map (
            O => \N__17195\,
            I => \N__17121\
        );

    \I__4078\ : Span4Mux_v
    port map (
            O => \N__17190\,
            I => \N__17112\
        );

    \I__4077\ : Span4Mux_h
    port map (
            O => \N__17187\,
            I => \N__17112\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__17180\,
            I => \N__17112\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__17177\,
            I => \N__17112\
        );

    \I__4074\ : Span4Mux_h
    port map (
            O => \N__17174\,
            I => \N__17109\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__17171\,
            I => \N__17106\
        );

    \I__4072\ : Span12Mux_h
    port map (
            O => \N__17168\,
            I => \N__17103\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__17165\,
            I => \N__17100\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__17158\,
            I => \N__17097\
        );

    \I__4069\ : Span4Mux_s1_v
    port map (
            O => \N__17155\,
            I => \N__17094\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__17152\,
            I => \N__17091\
        );

    \I__4067\ : ClkMux
    port map (
            O => \N__17151\,
            I => \N__17088\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__17148\,
            I => \N__17085\
        );

    \I__4065\ : Sp12to4
    port map (
            O => \N__17145\,
            I => \N__17080\
        );

    \I__4064\ : Sp12to4
    port map (
            O => \N__17140\,
            I => \N__17080\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__17137\,
            I => \N__17075\
        );

    \I__4062\ : Sp12to4
    port map (
            O => \N__17130\,
            I => \N__17075\
        );

    \I__4061\ : Span12Mux_h
    port map (
            O => \N__17127\,
            I => \N__17068\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__17124\,
            I => \N__17068\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__17121\,
            I => \N__17068\
        );

    \I__4058\ : Span4Mux_v
    port map (
            O => \N__17112\,
            I => \N__17065\
        );

    \I__4057\ : Span4Mux_v
    port map (
            O => \N__17109\,
            I => \N__17060\
        );

    \I__4056\ : Span4Mux_h
    port map (
            O => \N__17106\,
            I => \N__17060\
        );

    \I__4055\ : Span12Mux_v
    port map (
            O => \N__17103\,
            I => \N__17055\
        );

    \I__4054\ : Span12Mux_h
    port map (
            O => \N__17100\,
            I => \N__17055\
        );

    \I__4053\ : Sp12to4
    port map (
            O => \N__17097\,
            I => \N__17048\
        );

    \I__4052\ : Sp12to4
    port map (
            O => \N__17094\,
            I => \N__17048\
        );

    \I__4051\ : Sp12to4
    port map (
            O => \N__17091\,
            I => \N__17048\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__17088\,
            I => \N__17045\
        );

    \I__4049\ : Span12Mux_h
    port map (
            O => \N__17085\,
            I => \N__17042\
        );

    \I__4048\ : Span12Mux_h
    port map (
            O => \N__17080\,
            I => \N__17033\
        );

    \I__4047\ : Span12Mux_h
    port map (
            O => \N__17075\,
            I => \N__17033\
        );

    \I__4046\ : Span12Mux_v
    port map (
            O => \N__17068\,
            I => \N__17033\
        );

    \I__4045\ : Sp12to4
    port map (
            O => \N__17065\,
            I => \N__17033\
        );

    \I__4044\ : Span4Mux_h
    port map (
            O => \N__17060\,
            I => \N__17030\
        );

    \I__4043\ : Span12Mux_v
    port map (
            O => \N__17055\,
            I => \N__17023\
        );

    \I__4042\ : Span12Mux_h
    port map (
            O => \N__17048\,
            I => \N__17023\
        );

    \I__4041\ : Span12Mux_h
    port map (
            O => \N__17045\,
            I => \N__17023\
        );

    \I__4040\ : Odrv12
    port map (
            O => \N__17042\,
            I => \ADV_CLK_c\
        );

    \I__4039\ : Odrv12
    port map (
            O => \N__17033\,
            I => \ADV_CLK_c\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__17030\,
            I => \ADV_CLK_c\
        );

    \I__4037\ : Odrv12
    port map (
            O => \N__17023\,
            I => \ADV_CLK_c\
        );

    \I__4036\ : InMux
    port map (
            O => \N__17014\,
            I => \N__17011\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__17011\,
            I => \N__17008\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__17008\,
            I => \N__17005\
        );

    \I__4033\ : Span4Mux_h
    port map (
            O => \N__17005\,
            I => \N__17002\
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__17002\,
            I => \line_buffer.n716\
        );

    \I__4031\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16996\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__16996\,
            I => \N__16993\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__16993\,
            I => \N__16990\
        );

    \I__4028\ : Span4Mux_v
    port map (
            O => \N__16990\,
            I => \N__16987\
        );

    \I__4027\ : Sp12to4
    port map (
            O => \N__16987\,
            I => \N__16984\
        );

    \I__4026\ : Odrv12
    port map (
            O => \N__16984\,
            I => \line_buffer.n724\
        );

    \I__4025\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16978\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__16978\,
            I => \line_buffer.n3046\
        );

    \I__4023\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16972\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__16972\,
            I => \N__16969\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__16969\,
            I => \receive_module.n132\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__16966\,
            I => \N__16963\
        );

    \I__4019\ : CascadeBuf
    port map (
            O => \N__16963\,
            I => \N__16959\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__16962\,
            I => \N__16956\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__16959\,
            I => \N__16953\
        );

    \I__4016\ : CascadeBuf
    port map (
            O => \N__16956\,
            I => \N__16950\
        );

    \I__4015\ : CascadeBuf
    port map (
            O => \N__16953\,
            I => \N__16947\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__16950\,
            I => \N__16944\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__16947\,
            I => \N__16941\
        );

    \I__4012\ : CascadeBuf
    port map (
            O => \N__16944\,
            I => \N__16938\
        );

    \I__4011\ : CascadeBuf
    port map (
            O => \N__16941\,
            I => \N__16935\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__16938\,
            I => \N__16932\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__16935\,
            I => \N__16929\
        );

    \I__4008\ : CascadeBuf
    port map (
            O => \N__16932\,
            I => \N__16926\
        );

    \I__4007\ : CascadeBuf
    port map (
            O => \N__16929\,
            I => \N__16923\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__16926\,
            I => \N__16920\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__16923\,
            I => \N__16917\
        );

    \I__4004\ : CascadeBuf
    port map (
            O => \N__16920\,
            I => \N__16914\
        );

    \I__4003\ : CascadeBuf
    port map (
            O => \N__16917\,
            I => \N__16911\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__16914\,
            I => \N__16908\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__16911\,
            I => \N__16905\
        );

    \I__4000\ : CascadeBuf
    port map (
            O => \N__16908\,
            I => \N__16902\
        );

    \I__3999\ : CascadeBuf
    port map (
            O => \N__16905\,
            I => \N__16899\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__16902\,
            I => \N__16896\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__16899\,
            I => \N__16893\
        );

    \I__3996\ : CascadeBuf
    port map (
            O => \N__16896\,
            I => \N__16890\
        );

    \I__3995\ : CascadeBuf
    port map (
            O => \N__16893\,
            I => \N__16887\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__16890\,
            I => \N__16884\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__16887\,
            I => \N__16881\
        );

    \I__3992\ : CascadeBuf
    port map (
            O => \N__16884\,
            I => \N__16878\
        );

    \I__3991\ : CascadeBuf
    port map (
            O => \N__16881\,
            I => \N__16875\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__16878\,
            I => \N__16872\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__16875\,
            I => \N__16869\
        );

    \I__3988\ : CascadeBuf
    port map (
            O => \N__16872\,
            I => \N__16866\
        );

    \I__3987\ : CascadeBuf
    port map (
            O => \N__16869\,
            I => \N__16863\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__16866\,
            I => \N__16860\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__16863\,
            I => \N__16857\
        );

    \I__3984\ : CascadeBuf
    port map (
            O => \N__16860\,
            I => \N__16854\
        );

    \I__3983\ : CascadeBuf
    port map (
            O => \N__16857\,
            I => \N__16851\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__16854\,
            I => \N__16848\
        );

    \I__3981\ : CascadeMux
    port map (
            O => \N__16851\,
            I => \N__16845\
        );

    \I__3980\ : CascadeBuf
    port map (
            O => \N__16848\,
            I => \N__16842\
        );

    \I__3979\ : CascadeBuf
    port map (
            O => \N__16845\,
            I => \N__16839\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__16842\,
            I => \N__16836\
        );

    \I__3977\ : CascadeMux
    port map (
            O => \N__16839\,
            I => \N__16833\
        );

    \I__3976\ : CascadeBuf
    port map (
            O => \N__16836\,
            I => \N__16830\
        );

    \I__3975\ : CascadeBuf
    port map (
            O => \N__16833\,
            I => \N__16827\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__16830\,
            I => \N__16824\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__16827\,
            I => \N__16821\
        );

    \I__3972\ : CascadeBuf
    port map (
            O => \N__16824\,
            I => \N__16818\
        );

    \I__3971\ : CascadeBuf
    port map (
            O => \N__16821\,
            I => \N__16815\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__16818\,
            I => \N__16812\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__16815\,
            I => \N__16809\
        );

    \I__3968\ : CascadeBuf
    port map (
            O => \N__16812\,
            I => \N__16806\
        );

    \I__3967\ : CascadeBuf
    port map (
            O => \N__16809\,
            I => \N__16803\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__16806\,
            I => \N__16800\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__16803\,
            I => \N__16797\
        );

    \I__3964\ : CascadeBuf
    port map (
            O => \N__16800\,
            I => \N__16794\
        );

    \I__3963\ : CascadeBuf
    port map (
            O => \N__16797\,
            I => \N__16791\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__16794\,
            I => \N__16788\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__16791\,
            I => \N__16785\
        );

    \I__3960\ : CascadeBuf
    port map (
            O => \N__16788\,
            I => \N__16782\
        );

    \I__3959\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16779\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__16782\,
            I => \N__16776\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__16779\,
            I => \N__16773\
        );

    \I__3956\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16770\
        );

    \I__3955\ : Span4Mux_h
    port map (
            O => \N__16773\,
            I => \N__16767\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__16770\,
            I => \N__16764\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__16767\,
            I => \N__16760\
        );

    \I__3952\ : Span12Mux_s1_v
    port map (
            O => \N__16764\,
            I => \N__16757\
        );

    \I__3951\ : InMux
    port map (
            O => \N__16763\,
            I => \N__16754\
        );

    \I__3950\ : Sp12to4
    port map (
            O => \N__16760\,
            I => \N__16750\
        );

    \I__3949\ : Span12Mux_v
    port map (
            O => \N__16757\,
            I => \N__16747\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__16754\,
            I => \N__16744\
        );

    \I__3947\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16741\
        );

    \I__3946\ : Span12Mux_v
    port map (
            O => \N__16750\,
            I => \N__16736\
        );

    \I__3945\ : Span12Mux_h
    port map (
            O => \N__16747\,
            I => \N__16736\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__16744\,
            I => \RX_ADDR_4\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__16741\,
            I => \RX_ADDR_4\
        );

    \I__3942\ : Odrv12
    port map (
            O => \N__16736\,
            I => \RX_ADDR_4\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__16729\,
            I => \N__16726\
        );

    \I__3940\ : InMux
    port map (
            O => \N__16726\,
            I => \N__16723\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__16723\,
            I => \N__16720\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__16720\,
            I => \receive_module.n130\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__16717\,
            I => \N__16713\
        );

    \I__3936\ : CascadeMux
    port map (
            O => \N__16716\,
            I => \N__16710\
        );

    \I__3935\ : CascadeBuf
    port map (
            O => \N__16713\,
            I => \N__16707\
        );

    \I__3934\ : CascadeBuf
    port map (
            O => \N__16710\,
            I => \N__16704\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__16707\,
            I => \N__16701\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__16704\,
            I => \N__16698\
        );

    \I__3931\ : CascadeBuf
    port map (
            O => \N__16701\,
            I => \N__16695\
        );

    \I__3930\ : CascadeBuf
    port map (
            O => \N__16698\,
            I => \N__16692\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__16695\,
            I => \N__16689\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__16692\,
            I => \N__16686\
        );

    \I__3927\ : CascadeBuf
    port map (
            O => \N__16689\,
            I => \N__16683\
        );

    \I__3926\ : CascadeBuf
    port map (
            O => \N__16686\,
            I => \N__16680\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__16683\,
            I => \N__16677\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__16680\,
            I => \N__16674\
        );

    \I__3923\ : CascadeBuf
    port map (
            O => \N__16677\,
            I => \N__16671\
        );

    \I__3922\ : CascadeBuf
    port map (
            O => \N__16674\,
            I => \N__16668\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__16671\,
            I => \N__16665\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__16668\,
            I => \N__16662\
        );

    \I__3919\ : CascadeBuf
    port map (
            O => \N__16665\,
            I => \N__16659\
        );

    \I__3918\ : CascadeBuf
    port map (
            O => \N__16662\,
            I => \N__16656\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__16659\,
            I => \N__16653\
        );

    \I__3916\ : CascadeMux
    port map (
            O => \N__16656\,
            I => \N__16650\
        );

    \I__3915\ : CascadeBuf
    port map (
            O => \N__16653\,
            I => \N__16647\
        );

    \I__3914\ : CascadeBuf
    port map (
            O => \N__16650\,
            I => \N__16644\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__16647\,
            I => \N__16641\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__16644\,
            I => \N__16638\
        );

    \I__3911\ : CascadeBuf
    port map (
            O => \N__16641\,
            I => \N__16635\
        );

    \I__3910\ : CascadeBuf
    port map (
            O => \N__16638\,
            I => \N__16632\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__16635\,
            I => \N__16629\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__16632\,
            I => \N__16626\
        );

    \I__3907\ : CascadeBuf
    port map (
            O => \N__16629\,
            I => \N__16623\
        );

    \I__3906\ : CascadeBuf
    port map (
            O => \N__16626\,
            I => \N__16620\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__16623\,
            I => \N__16617\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__16620\,
            I => \N__16614\
        );

    \I__3903\ : CascadeBuf
    port map (
            O => \N__16617\,
            I => \N__16611\
        );

    \I__3902\ : CascadeBuf
    port map (
            O => \N__16614\,
            I => \N__16608\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__16611\,
            I => \N__16605\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__16608\,
            I => \N__16602\
        );

    \I__3899\ : CascadeBuf
    port map (
            O => \N__16605\,
            I => \N__16599\
        );

    \I__3898\ : CascadeBuf
    port map (
            O => \N__16602\,
            I => \N__16596\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__16599\,
            I => \N__16593\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__16596\,
            I => \N__16590\
        );

    \I__3895\ : CascadeBuf
    port map (
            O => \N__16593\,
            I => \N__16587\
        );

    \I__3894\ : CascadeBuf
    port map (
            O => \N__16590\,
            I => \N__16584\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__16587\,
            I => \N__16581\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__16584\,
            I => \N__16578\
        );

    \I__3891\ : CascadeBuf
    port map (
            O => \N__16581\,
            I => \N__16575\
        );

    \I__3890\ : CascadeBuf
    port map (
            O => \N__16578\,
            I => \N__16572\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__16575\,
            I => \N__16569\
        );

    \I__3888\ : CascadeMux
    port map (
            O => \N__16572\,
            I => \N__16566\
        );

    \I__3887\ : CascadeBuf
    port map (
            O => \N__16569\,
            I => \N__16563\
        );

    \I__3886\ : CascadeBuf
    port map (
            O => \N__16566\,
            I => \N__16560\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__16563\,
            I => \N__16557\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__16560\,
            I => \N__16554\
        );

    \I__3883\ : CascadeBuf
    port map (
            O => \N__16557\,
            I => \N__16551\
        );

    \I__3882\ : CascadeBuf
    port map (
            O => \N__16554\,
            I => \N__16548\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__16551\,
            I => \N__16545\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__16548\,
            I => \N__16542\
        );

    \I__3879\ : CascadeBuf
    port map (
            O => \N__16545\,
            I => \N__16539\
        );

    \I__3878\ : CascadeBuf
    port map (
            O => \N__16542\,
            I => \N__16536\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__16539\,
            I => \N__16533\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__16536\,
            I => \N__16530\
        );

    \I__3875\ : InMux
    port map (
            O => \N__16533\,
            I => \N__16527\
        );

    \I__3874\ : InMux
    port map (
            O => \N__16530\,
            I => \N__16524\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__16527\,
            I => \N__16520\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__16524\,
            I => \N__16517\
        );

    \I__3871\ : InMux
    port map (
            O => \N__16523\,
            I => \N__16514\
        );

    \I__3870\ : Span12Mux_h
    port map (
            O => \N__16520\,
            I => \N__16508\
        );

    \I__3869\ : Span12Mux_h
    port map (
            O => \N__16517\,
            I => \N__16508\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__16514\,
            I => \N__16505\
        );

    \I__3867\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16502\
        );

    \I__3866\ : Span12Mux_v
    port map (
            O => \N__16508\,
            I => \N__16499\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__16505\,
            I => \RX_ADDR_6\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__16502\,
            I => \RX_ADDR_6\
        );

    \I__3863\ : Odrv12
    port map (
            O => \N__16499\,
            I => \RX_ADDR_6\
        );

    \I__3862\ : InMux
    port map (
            O => \N__16492\,
            I => \N__16489\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__16489\,
            I => \N__16486\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__16486\,
            I => \receive_module.n126\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__16483\,
            I => \N__16476\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__16482\,
            I => \N__16472\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__16481\,
            I => \N__16467\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__16480\,
            I => \N__16463\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__16479\,
            I => \N__16460\
        );

    \I__3854\ : InMux
    port map (
            O => \N__16476\,
            I => \N__16457\
        );

    \I__3853\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16452\
        );

    \I__3852\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16452\
        );

    \I__3851\ : InMux
    port map (
            O => \N__16471\,
            I => \N__16449\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__16470\,
            I => \N__16446\
        );

    \I__3849\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16440\
        );

    \I__3848\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16433\
        );

    \I__3847\ : InMux
    port map (
            O => \N__16463\,
            I => \N__16433\
        );

    \I__3846\ : InMux
    port map (
            O => \N__16460\,
            I => \N__16433\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__16457\,
            I => \N__16427\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__16452\,
            I => \N__16427\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__16449\,
            I => \N__16424\
        );

    \I__3842\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16415\
        );

    \I__3841\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16415\
        );

    \I__3840\ : InMux
    port map (
            O => \N__16444\,
            I => \N__16415\
        );

    \I__3839\ : InMux
    port map (
            O => \N__16443\,
            I => \N__16415\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__16440\,
            I => \N__16410\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__16433\,
            I => \N__16410\
        );

    \I__3836\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16407\
        );

    \I__3835\ : Span4Mux_v
    port map (
            O => \N__16427\,
            I => \N__16402\
        );

    \I__3834\ : Span4Mux_v
    port map (
            O => \N__16424\,
            I => \N__16399\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__16415\,
            I => \N__16392\
        );

    \I__3832\ : Span4Mux_h
    port map (
            O => \N__16410\,
            I => \N__16392\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__16407\,
            I => \N__16392\
        );

    \I__3830\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16387\
        );

    \I__3829\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16387\
        );

    \I__3828\ : Span4Mux_h
    port map (
            O => \N__16402\,
            I => \N__16377\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__16399\,
            I => \N__16377\
        );

    \I__3826\ : Span4Mux_v
    port map (
            O => \N__16392\,
            I => \N__16377\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__16387\,
            I => \N__16377\
        );

    \I__3824\ : InMux
    port map (
            O => \N__16386\,
            I => \N__16374\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__16377\,
            I => \N__16371\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__16374\,
            I => \N__16368\
        );

    \I__3821\ : Span4Mux_v
    port map (
            O => \N__16371\,
            I => \N__16365\
        );

    \I__3820\ : Span12Mux_v
    port map (
            O => \N__16368\,
            I => \N__16362\
        );

    \I__3819\ : IoSpan4Mux
    port map (
            O => \N__16365\,
            I => \N__16359\
        );

    \I__3818\ : Odrv12
    port map (
            O => \N__16362\,
            I => \TVP_VSYNC_c\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__16359\,
            I => \TVP_VSYNC_c\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__16354\,
            I => \N__16350\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__16353\,
            I => \N__16347\
        );

    \I__3814\ : CascadeBuf
    port map (
            O => \N__16350\,
            I => \N__16344\
        );

    \I__3813\ : CascadeBuf
    port map (
            O => \N__16347\,
            I => \N__16341\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__16344\,
            I => \N__16338\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__16341\,
            I => \N__16335\
        );

    \I__3810\ : CascadeBuf
    port map (
            O => \N__16338\,
            I => \N__16332\
        );

    \I__3809\ : CascadeBuf
    port map (
            O => \N__16335\,
            I => \N__16329\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__16332\,
            I => \N__16326\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__16329\,
            I => \N__16323\
        );

    \I__3806\ : CascadeBuf
    port map (
            O => \N__16326\,
            I => \N__16320\
        );

    \I__3805\ : CascadeBuf
    port map (
            O => \N__16323\,
            I => \N__16317\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__16320\,
            I => \N__16314\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__16317\,
            I => \N__16311\
        );

    \I__3802\ : CascadeBuf
    port map (
            O => \N__16314\,
            I => \N__16308\
        );

    \I__3801\ : CascadeBuf
    port map (
            O => \N__16311\,
            I => \N__16305\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__16308\,
            I => \N__16302\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__16305\,
            I => \N__16299\
        );

    \I__3798\ : CascadeBuf
    port map (
            O => \N__16302\,
            I => \N__16296\
        );

    \I__3797\ : CascadeBuf
    port map (
            O => \N__16299\,
            I => \N__16293\
        );

    \I__3796\ : CascadeMux
    port map (
            O => \N__16296\,
            I => \N__16290\
        );

    \I__3795\ : CascadeMux
    port map (
            O => \N__16293\,
            I => \N__16287\
        );

    \I__3794\ : CascadeBuf
    port map (
            O => \N__16290\,
            I => \N__16284\
        );

    \I__3793\ : CascadeBuf
    port map (
            O => \N__16287\,
            I => \N__16281\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__16284\,
            I => \N__16278\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__16281\,
            I => \N__16275\
        );

    \I__3790\ : CascadeBuf
    port map (
            O => \N__16278\,
            I => \N__16272\
        );

    \I__3789\ : CascadeBuf
    port map (
            O => \N__16275\,
            I => \N__16269\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__16272\,
            I => \N__16266\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__16269\,
            I => \N__16263\
        );

    \I__3786\ : CascadeBuf
    port map (
            O => \N__16266\,
            I => \N__16260\
        );

    \I__3785\ : CascadeBuf
    port map (
            O => \N__16263\,
            I => \N__16257\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__16260\,
            I => \N__16254\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__16257\,
            I => \N__16251\
        );

    \I__3782\ : CascadeBuf
    port map (
            O => \N__16254\,
            I => \N__16248\
        );

    \I__3781\ : CascadeBuf
    port map (
            O => \N__16251\,
            I => \N__16245\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__16248\,
            I => \N__16242\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__16245\,
            I => \N__16239\
        );

    \I__3778\ : CascadeBuf
    port map (
            O => \N__16242\,
            I => \N__16236\
        );

    \I__3777\ : CascadeBuf
    port map (
            O => \N__16239\,
            I => \N__16233\
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__16236\,
            I => \N__16230\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__16233\,
            I => \N__16227\
        );

    \I__3774\ : CascadeBuf
    port map (
            O => \N__16230\,
            I => \N__16224\
        );

    \I__3773\ : CascadeBuf
    port map (
            O => \N__16227\,
            I => \N__16221\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__16224\,
            I => \N__16218\
        );

    \I__3771\ : CascadeMux
    port map (
            O => \N__16221\,
            I => \N__16215\
        );

    \I__3770\ : CascadeBuf
    port map (
            O => \N__16218\,
            I => \N__16212\
        );

    \I__3769\ : CascadeBuf
    port map (
            O => \N__16215\,
            I => \N__16209\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__16212\,
            I => \N__16206\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__16209\,
            I => \N__16203\
        );

    \I__3766\ : CascadeBuf
    port map (
            O => \N__16206\,
            I => \N__16200\
        );

    \I__3765\ : CascadeBuf
    port map (
            O => \N__16203\,
            I => \N__16197\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__16200\,
            I => \N__16194\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__16197\,
            I => \N__16191\
        );

    \I__3762\ : CascadeBuf
    port map (
            O => \N__16194\,
            I => \N__16188\
        );

    \I__3761\ : CascadeBuf
    port map (
            O => \N__16191\,
            I => \N__16185\
        );

    \I__3760\ : CascadeMux
    port map (
            O => \N__16188\,
            I => \N__16182\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__16185\,
            I => \N__16179\
        );

    \I__3758\ : CascadeBuf
    port map (
            O => \N__16182\,
            I => \N__16176\
        );

    \I__3757\ : CascadeBuf
    port map (
            O => \N__16179\,
            I => \N__16173\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__16176\,
            I => \N__16170\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__16173\,
            I => \N__16167\
        );

    \I__3754\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16164\
        );

    \I__3753\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16161\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__16164\,
            I => \N__16157\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__16161\,
            I => \N__16154\
        );

    \I__3750\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16151\
        );

    \I__3749\ : Span12Mux_h
    port map (
            O => \N__16157\,
            I => \N__16145\
        );

    \I__3748\ : Span12Mux_h
    port map (
            O => \N__16154\,
            I => \N__16145\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__16151\,
            I => \N__16142\
        );

    \I__3746\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16139\
        );

    \I__3745\ : Span12Mux_v
    port map (
            O => \N__16145\,
            I => \N__16136\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__16142\,
            I => \RX_ADDR_10\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__16139\,
            I => \RX_ADDR_10\
        );

    \I__3742\ : Odrv12
    port map (
            O => \N__16136\,
            I => \RX_ADDR_10\
        );

    \I__3741\ : InMux
    port map (
            O => \N__16129\,
            I => \N__16126\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__16126\,
            I => \N__16115\
        );

    \I__3739\ : ClkMux
    port map (
            O => \N__16125\,
            I => \N__15985\
        );

    \I__3738\ : ClkMux
    port map (
            O => \N__16124\,
            I => \N__15985\
        );

    \I__3737\ : ClkMux
    port map (
            O => \N__16123\,
            I => \N__15985\
        );

    \I__3736\ : ClkMux
    port map (
            O => \N__16122\,
            I => \N__15985\
        );

    \I__3735\ : ClkMux
    port map (
            O => \N__16121\,
            I => \N__15985\
        );

    \I__3734\ : ClkMux
    port map (
            O => \N__16120\,
            I => \N__15985\
        );

    \I__3733\ : ClkMux
    port map (
            O => \N__16119\,
            I => \N__15985\
        );

    \I__3732\ : ClkMux
    port map (
            O => \N__16118\,
            I => \N__15985\
        );

    \I__3731\ : Glb2LocalMux
    port map (
            O => \N__16115\,
            I => \N__15985\
        );

    \I__3730\ : ClkMux
    port map (
            O => \N__16114\,
            I => \N__15985\
        );

    \I__3729\ : ClkMux
    port map (
            O => \N__16113\,
            I => \N__15985\
        );

    \I__3728\ : ClkMux
    port map (
            O => \N__16112\,
            I => \N__15985\
        );

    \I__3727\ : ClkMux
    port map (
            O => \N__16111\,
            I => \N__15985\
        );

    \I__3726\ : ClkMux
    port map (
            O => \N__16110\,
            I => \N__15985\
        );

    \I__3725\ : ClkMux
    port map (
            O => \N__16109\,
            I => \N__15985\
        );

    \I__3724\ : ClkMux
    port map (
            O => \N__16108\,
            I => \N__15985\
        );

    \I__3723\ : ClkMux
    port map (
            O => \N__16107\,
            I => \N__15985\
        );

    \I__3722\ : ClkMux
    port map (
            O => \N__16106\,
            I => \N__15985\
        );

    \I__3721\ : ClkMux
    port map (
            O => \N__16105\,
            I => \N__15985\
        );

    \I__3720\ : ClkMux
    port map (
            O => \N__16104\,
            I => \N__15985\
        );

    \I__3719\ : ClkMux
    port map (
            O => \N__16103\,
            I => \N__15985\
        );

    \I__3718\ : ClkMux
    port map (
            O => \N__16102\,
            I => \N__15985\
        );

    \I__3717\ : ClkMux
    port map (
            O => \N__16101\,
            I => \N__15985\
        );

    \I__3716\ : ClkMux
    port map (
            O => \N__16100\,
            I => \N__15985\
        );

    \I__3715\ : ClkMux
    port map (
            O => \N__16099\,
            I => \N__15985\
        );

    \I__3714\ : ClkMux
    port map (
            O => \N__16098\,
            I => \N__15985\
        );

    \I__3713\ : ClkMux
    port map (
            O => \N__16097\,
            I => \N__15985\
        );

    \I__3712\ : ClkMux
    port map (
            O => \N__16096\,
            I => \N__15985\
        );

    \I__3711\ : ClkMux
    port map (
            O => \N__16095\,
            I => \N__15985\
        );

    \I__3710\ : ClkMux
    port map (
            O => \N__16094\,
            I => \N__15985\
        );

    \I__3709\ : ClkMux
    port map (
            O => \N__16093\,
            I => \N__15985\
        );

    \I__3708\ : ClkMux
    port map (
            O => \N__16092\,
            I => \N__15985\
        );

    \I__3707\ : ClkMux
    port map (
            O => \N__16091\,
            I => \N__15985\
        );

    \I__3706\ : ClkMux
    port map (
            O => \N__16090\,
            I => \N__15985\
        );

    \I__3705\ : ClkMux
    port map (
            O => \N__16089\,
            I => \N__15985\
        );

    \I__3704\ : ClkMux
    port map (
            O => \N__16088\,
            I => \N__15985\
        );

    \I__3703\ : ClkMux
    port map (
            O => \N__16087\,
            I => \N__15985\
        );

    \I__3702\ : ClkMux
    port map (
            O => \N__16086\,
            I => \N__15985\
        );

    \I__3701\ : ClkMux
    port map (
            O => \N__16085\,
            I => \N__15985\
        );

    \I__3700\ : ClkMux
    port map (
            O => \N__16084\,
            I => \N__15985\
        );

    \I__3699\ : ClkMux
    port map (
            O => \N__16083\,
            I => \N__15985\
        );

    \I__3698\ : ClkMux
    port map (
            O => \N__16082\,
            I => \N__15985\
        );

    \I__3697\ : ClkMux
    port map (
            O => \N__16081\,
            I => \N__15985\
        );

    \I__3696\ : ClkMux
    port map (
            O => \N__16080\,
            I => \N__15985\
        );

    \I__3695\ : ClkMux
    port map (
            O => \N__16079\,
            I => \N__15985\
        );

    \I__3694\ : ClkMux
    port map (
            O => \N__16078\,
            I => \N__15985\
        );

    \I__3693\ : GlobalMux
    port map (
            O => \N__15985\,
            I => \N__15982\
        );

    \I__3692\ : gio2CtrlBuf
    port map (
            O => \N__15982\,
            I => \TVP_CLK_c\
        );

    \I__3691\ : SRMux
    port map (
            O => \N__15979\,
            I => \N__15975\
        );

    \I__3690\ : SRMux
    port map (
            O => \N__15978\,
            I => \N__15972\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__15975\,
            I => \N__15969\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__15972\,
            I => \N__15961\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__15969\,
            I => \N__15958\
        );

    \I__3686\ : SRMux
    port map (
            O => \N__15968\,
            I => \N__15955\
        );

    \I__3685\ : SRMux
    port map (
            O => \N__15967\,
            I => \N__15952\
        );

    \I__3684\ : SRMux
    port map (
            O => \N__15966\,
            I => \N__15949\
        );

    \I__3683\ : SRMux
    port map (
            O => \N__15965\,
            I => \N__15946\
        );

    \I__3682\ : SRMux
    port map (
            O => \N__15964\,
            I => \N__15943\
        );

    \I__3681\ : Span4Mux_v
    port map (
            O => \N__15961\,
            I => \N__15940\
        );

    \I__3680\ : Span4Mux_h
    port map (
            O => \N__15958\,
            I => \N__15933\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__15955\,
            I => \N__15933\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__15952\,
            I => \N__15933\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__15949\,
            I => \N__15928\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__15946\,
            I => \N__15928\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__15943\,
            I => \N__15925\
        );

    \I__3674\ : Span4Mux_h
    port map (
            O => \N__15940\,
            I => \N__15920\
        );

    \I__3673\ : Span4Mux_v
    port map (
            O => \N__15933\,
            I => \N__15920\
        );

    \I__3672\ : Span4Mux_v
    port map (
            O => \N__15928\,
            I => \N__15917\
        );

    \I__3671\ : Sp12to4
    port map (
            O => \N__15925\,
            I => \N__15914\
        );

    \I__3670\ : Span4Mux_h
    port map (
            O => \N__15920\,
            I => \N__15911\
        );

    \I__3669\ : Odrv4
    port map (
            O => \N__15917\,
            I => \receive_module.n3185\
        );

    \I__3668\ : Odrv12
    port map (
            O => \N__15914\,
            I => \receive_module.n3185\
        );

    \I__3667\ : Odrv4
    port map (
            O => \N__15911\,
            I => \receive_module.n3185\
        );

    \I__3666\ : InMux
    port map (
            O => \N__15904\,
            I => \N__15901\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__15901\,
            I => \N__15898\
        );

    \I__3664\ : Span12Mux_v
    port map (
            O => \N__15898\,
            I => \N__15895\
        );

    \I__3663\ : Odrv12
    port map (
            O => \N__15895\,
            I => \line_buffer.n757\
        );

    \I__3662\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15889\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__15889\,
            I => \N__15886\
        );

    \I__3660\ : Span4Mux_v
    port map (
            O => \N__15886\,
            I => \N__15883\
        );

    \I__3659\ : Span4Mux_v
    port map (
            O => \N__15883\,
            I => \N__15880\
        );

    \I__3658\ : Span4Mux_h
    port map (
            O => \N__15880\,
            I => \N__15877\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__15877\,
            I => \line_buffer.n749\
        );

    \I__3656\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15871\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__15871\,
            I => \N__15868\
        );

    \I__3654\ : Span4Mux_v
    port map (
            O => \N__15868\,
            I => \N__15865\
        );

    \I__3653\ : Span4Mux_h
    port map (
            O => \N__15865\,
            I => \N__15862\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__15862\,
            I => \N__15859\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__15859\,
            I => \line_buffer.n685\
        );

    \I__3650\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15853\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__15853\,
            I => \N__15850\
        );

    \I__3648\ : Span12Mux_v
    port map (
            O => \N__15850\,
            I => \N__15847\
        );

    \I__3647\ : Span12Mux_h
    port map (
            O => \N__15847\,
            I => \N__15844\
        );

    \I__3646\ : Odrv12
    port map (
            O => \N__15844\,
            I => \line_buffer.n693\
        );

    \I__3645\ : CascadeMux
    port map (
            O => \N__15841\,
            I => \line_buffer.n3155_cascade_\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__15838\,
            I => \N__15831\
        );

    \I__3643\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15827\
        );

    \I__3642\ : CascadeMux
    port map (
            O => \N__15836\,
            I => \N__15822\
        );

    \I__3641\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15819\
        );

    \I__3640\ : InMux
    port map (
            O => \N__15834\,
            I => \N__15814\
        );

    \I__3639\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15814\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__15830\,
            I => \N__15804\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__15827\,
            I => \N__15801\
        );

    \I__3636\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15794\
        );

    \I__3635\ : InMux
    port map (
            O => \N__15825\,
            I => \N__15794\
        );

    \I__3634\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15794\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__15819\,
            I => \N__15789\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__15814\,
            I => \N__15789\
        );

    \I__3631\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15786\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__15812\,
            I => \N__15782\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__15811\,
            I => \N__15778\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__15810\,
            I => \N__15773\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__15809\,
            I => \N__15769\
        );

    \I__3626\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15761\
        );

    \I__3625\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15761\
        );

    \I__3624\ : InMux
    port map (
            O => \N__15804\,
            I => \N__15761\
        );

    \I__3623\ : Span4Mux_h
    port map (
            O => \N__15801\,
            I => \N__15756\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__15794\,
            I => \N__15756\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__15789\,
            I => \N__15751\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__15786\,
            I => \N__15751\
        );

    \I__3619\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15746\
        );

    \I__3618\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15746\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__15781\,
            I => \N__15742\
        );

    \I__3616\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15739\
        );

    \I__3615\ : InMux
    port map (
            O => \N__15777\,
            I => \N__15736\
        );

    \I__3614\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15733\
        );

    \I__3613\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15730\
        );

    \I__3612\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15727\
        );

    \I__3611\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15724\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__15768\,
            I => \N__15720\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__15761\,
            I => \N__15716\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__15756\,
            I => \N__15713\
        );

    \I__3607\ : Span4Mux_v
    port map (
            O => \N__15751\,
            I => \N__15708\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__15746\,
            I => \N__15708\
        );

    \I__3605\ : InMux
    port map (
            O => \N__15745\,
            I => \N__15703\
        );

    \I__3604\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15703\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__15739\,
            I => \N__15700\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__15736\,
            I => \N__15697\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__15733\,
            I => \N__15694\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__15730\,
            I => \N__15691\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__15727\,
            I => \N__15686\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__15724\,
            I => \N__15686\
        );

    \I__3597\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15683\
        );

    \I__3596\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15680\
        );

    \I__3595\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15677\
        );

    \I__3594\ : Span4Mux_h
    port map (
            O => \N__15716\,
            I => \N__15670\
        );

    \I__3593\ : Span4Mux_v
    port map (
            O => \N__15713\,
            I => \N__15670\
        );

    \I__3592\ : Span4Mux_h
    port map (
            O => \N__15708\,
            I => \N__15670\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__15703\,
            I => \N__15665\
        );

    \I__3590\ : Span12Mux_v
    port map (
            O => \N__15700\,
            I => \N__15665\
        );

    \I__3589\ : Span4Mux_h
    port map (
            O => \N__15697\,
            I => \N__15656\
        );

    \I__3588\ : Span4Mux_h
    port map (
            O => \N__15694\,
            I => \N__15656\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__15691\,
            I => \N__15656\
        );

    \I__3586\ : Span4Mux_h
    port map (
            O => \N__15686\,
            I => \N__15656\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__15683\,
            I => \TX_ADDR_12\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__15680\,
            I => \TX_ADDR_12\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__15677\,
            I => \TX_ADDR_12\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__15670\,
            I => \TX_ADDR_12\
        );

    \I__3581\ : Odrv12
    port map (
            O => \N__15665\,
            I => \TX_ADDR_12\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__15656\,
            I => \TX_ADDR_12\
        );

    \I__3579\ : InMux
    port map (
            O => \N__15643\,
            I => \N__15640\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__15640\,
            I => \line_buffer.n3158\
        );

    \I__3577\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15634\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15631\
        );

    \I__3575\ : Span4Mux_h
    port map (
            O => \N__15631\,
            I => \N__15628\
        );

    \I__3574\ : Span4Mux_h
    port map (
            O => \N__15628\,
            I => \N__15625\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__15625\,
            I => \line_buffer.n627\
        );

    \I__3572\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15619\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__15619\,
            I => \N__15616\
        );

    \I__3570\ : Span12Mux_v
    port map (
            O => \N__15616\,
            I => \N__15613\
        );

    \I__3569\ : Odrv12
    port map (
            O => \N__15613\,
            I => \line_buffer.n619\
        );

    \I__3568\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15607\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__15607\,
            I => \N__15604\
        );

    \I__3566\ : Span4Mux_v
    port map (
            O => \N__15604\,
            I => \N__15601\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__15601\,
            I => \line_buffer.n3045\
        );

    \I__3564\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15595\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__15595\,
            I => \N__15592\
        );

    \I__3562\ : Sp12to4
    port map (
            O => \N__15592\,
            I => \N__15589\
        );

    \I__3561\ : Span12Mux_v
    port map (
            O => \N__15589\,
            I => \N__15586\
        );

    \I__3560\ : Odrv12
    port map (
            O => \N__15586\,
            I => \line_buffer.n725\
        );

    \I__3559\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15580\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__15580\,
            I => \N__15577\
        );

    \I__3557\ : Odrv12
    port map (
            O => \N__15577\,
            I => \line_buffer.n717\
        );

    \I__3556\ : InMux
    port map (
            O => \N__15574\,
            I => \N__15571\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__15571\,
            I => \receive_module.n133\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__15568\,
            I => \N__15564\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__15567\,
            I => \N__15561\
        );

    \I__3552\ : CascadeBuf
    port map (
            O => \N__15564\,
            I => \N__15558\
        );

    \I__3551\ : CascadeBuf
    port map (
            O => \N__15561\,
            I => \N__15555\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__15558\,
            I => \N__15552\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__15555\,
            I => \N__15549\
        );

    \I__3548\ : CascadeBuf
    port map (
            O => \N__15552\,
            I => \N__15546\
        );

    \I__3547\ : CascadeBuf
    port map (
            O => \N__15549\,
            I => \N__15543\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__15546\,
            I => \N__15540\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__15543\,
            I => \N__15537\
        );

    \I__3544\ : CascadeBuf
    port map (
            O => \N__15540\,
            I => \N__15534\
        );

    \I__3543\ : CascadeBuf
    port map (
            O => \N__15537\,
            I => \N__15531\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__15534\,
            I => \N__15528\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__15531\,
            I => \N__15525\
        );

    \I__3540\ : CascadeBuf
    port map (
            O => \N__15528\,
            I => \N__15522\
        );

    \I__3539\ : CascadeBuf
    port map (
            O => \N__15525\,
            I => \N__15519\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__15522\,
            I => \N__15516\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__15519\,
            I => \N__15513\
        );

    \I__3536\ : CascadeBuf
    port map (
            O => \N__15516\,
            I => \N__15510\
        );

    \I__3535\ : CascadeBuf
    port map (
            O => \N__15513\,
            I => \N__15507\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__15510\,
            I => \N__15504\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__15507\,
            I => \N__15501\
        );

    \I__3532\ : CascadeBuf
    port map (
            O => \N__15504\,
            I => \N__15498\
        );

    \I__3531\ : CascadeBuf
    port map (
            O => \N__15501\,
            I => \N__15495\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__15498\,
            I => \N__15492\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__15495\,
            I => \N__15489\
        );

    \I__3528\ : CascadeBuf
    port map (
            O => \N__15492\,
            I => \N__15486\
        );

    \I__3527\ : CascadeBuf
    port map (
            O => \N__15489\,
            I => \N__15483\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__15486\,
            I => \N__15480\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__15483\,
            I => \N__15477\
        );

    \I__3524\ : CascadeBuf
    port map (
            O => \N__15480\,
            I => \N__15474\
        );

    \I__3523\ : CascadeBuf
    port map (
            O => \N__15477\,
            I => \N__15471\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__15474\,
            I => \N__15468\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__15471\,
            I => \N__15465\
        );

    \I__3520\ : CascadeBuf
    port map (
            O => \N__15468\,
            I => \N__15462\
        );

    \I__3519\ : CascadeBuf
    port map (
            O => \N__15465\,
            I => \N__15459\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__15462\,
            I => \N__15456\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__15459\,
            I => \N__15453\
        );

    \I__3516\ : CascadeBuf
    port map (
            O => \N__15456\,
            I => \N__15450\
        );

    \I__3515\ : CascadeBuf
    port map (
            O => \N__15453\,
            I => \N__15447\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__15450\,
            I => \N__15444\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__15447\,
            I => \N__15441\
        );

    \I__3512\ : CascadeBuf
    port map (
            O => \N__15444\,
            I => \N__15438\
        );

    \I__3511\ : CascadeBuf
    port map (
            O => \N__15441\,
            I => \N__15435\
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__15438\,
            I => \N__15432\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__15435\,
            I => \N__15429\
        );

    \I__3508\ : CascadeBuf
    port map (
            O => \N__15432\,
            I => \N__15426\
        );

    \I__3507\ : CascadeBuf
    port map (
            O => \N__15429\,
            I => \N__15423\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__15426\,
            I => \N__15420\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__15423\,
            I => \N__15417\
        );

    \I__3504\ : CascadeBuf
    port map (
            O => \N__15420\,
            I => \N__15414\
        );

    \I__3503\ : CascadeBuf
    port map (
            O => \N__15417\,
            I => \N__15411\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__15414\,
            I => \N__15408\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__15411\,
            I => \N__15405\
        );

    \I__3500\ : CascadeBuf
    port map (
            O => \N__15408\,
            I => \N__15402\
        );

    \I__3499\ : CascadeBuf
    port map (
            O => \N__15405\,
            I => \N__15399\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__15402\,
            I => \N__15396\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__15399\,
            I => \N__15393\
        );

    \I__3496\ : CascadeBuf
    port map (
            O => \N__15396\,
            I => \N__15390\
        );

    \I__3495\ : CascadeBuf
    port map (
            O => \N__15393\,
            I => \N__15387\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__15390\,
            I => \N__15384\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__15387\,
            I => \N__15381\
        );

    \I__3492\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15378\
        );

    \I__3491\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15375\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__15378\,
            I => \N__15372\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__15375\,
            I => \N__15369\
        );

    \I__3488\ : Span4Mux_v
    port map (
            O => \N__15372\,
            I => \N__15366\
        );

    \I__3487\ : Span4Mux_v
    port map (
            O => \N__15369\,
            I => \N__15363\
        );

    \I__3486\ : Sp12to4
    port map (
            O => \N__15366\,
            I => \N__15360\
        );

    \I__3485\ : Sp12to4
    port map (
            O => \N__15363\,
            I => \N__15357\
        );

    \I__3484\ : Span12Mux_h
    port map (
            O => \N__15360\,
            I => \N__15350\
        );

    \I__3483\ : Span12Mux_h
    port map (
            O => \N__15357\,
            I => \N__15350\
        );

    \I__3482\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15347\
        );

    \I__3481\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15344\
        );

    \I__3480\ : Span12Mux_v
    port map (
            O => \N__15350\,
            I => \N__15341\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__15347\,
            I => \RX_ADDR_3\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__15344\,
            I => \RX_ADDR_3\
        );

    \I__3477\ : Odrv12
    port map (
            O => \N__15341\,
            I => \RX_ADDR_3\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__15334\,
            I => \N__15331\
        );

    \I__3475\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15328\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__15328\,
            I => \receive_module.n134\
        );

    \I__3473\ : CascadeMux
    port map (
            O => \N__15325\,
            I => \N__15322\
        );

    \I__3472\ : CascadeBuf
    port map (
            O => \N__15322\,
            I => \N__15318\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__15321\,
            I => \N__15315\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__15318\,
            I => \N__15312\
        );

    \I__3469\ : CascadeBuf
    port map (
            O => \N__15315\,
            I => \N__15309\
        );

    \I__3468\ : CascadeBuf
    port map (
            O => \N__15312\,
            I => \N__15306\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__15309\,
            I => \N__15303\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__15306\,
            I => \N__15300\
        );

    \I__3465\ : CascadeBuf
    port map (
            O => \N__15303\,
            I => \N__15297\
        );

    \I__3464\ : CascadeBuf
    port map (
            O => \N__15300\,
            I => \N__15294\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__15297\,
            I => \N__15291\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__15294\,
            I => \N__15288\
        );

    \I__3461\ : CascadeBuf
    port map (
            O => \N__15291\,
            I => \N__15285\
        );

    \I__3460\ : CascadeBuf
    port map (
            O => \N__15288\,
            I => \N__15282\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__15285\,
            I => \N__15279\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__15282\,
            I => \N__15276\
        );

    \I__3457\ : CascadeBuf
    port map (
            O => \N__15279\,
            I => \N__15273\
        );

    \I__3456\ : CascadeBuf
    port map (
            O => \N__15276\,
            I => \N__15270\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__15273\,
            I => \N__15267\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__15270\,
            I => \N__15264\
        );

    \I__3453\ : CascadeBuf
    port map (
            O => \N__15267\,
            I => \N__15261\
        );

    \I__3452\ : CascadeBuf
    port map (
            O => \N__15264\,
            I => \N__15258\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__15261\,
            I => \N__15255\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__15258\,
            I => \N__15252\
        );

    \I__3449\ : CascadeBuf
    port map (
            O => \N__15255\,
            I => \N__15249\
        );

    \I__3448\ : CascadeBuf
    port map (
            O => \N__15252\,
            I => \N__15246\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__15249\,
            I => \N__15243\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__15246\,
            I => \N__15240\
        );

    \I__3445\ : CascadeBuf
    port map (
            O => \N__15243\,
            I => \N__15237\
        );

    \I__3444\ : CascadeBuf
    port map (
            O => \N__15240\,
            I => \N__15234\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__15237\,
            I => \N__15231\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__15234\,
            I => \N__15228\
        );

    \I__3441\ : CascadeBuf
    port map (
            O => \N__15231\,
            I => \N__15225\
        );

    \I__3440\ : CascadeBuf
    port map (
            O => \N__15228\,
            I => \N__15222\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__15225\,
            I => \N__15219\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__15222\,
            I => \N__15216\
        );

    \I__3437\ : CascadeBuf
    port map (
            O => \N__15219\,
            I => \N__15213\
        );

    \I__3436\ : CascadeBuf
    port map (
            O => \N__15216\,
            I => \N__15210\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__15213\,
            I => \N__15207\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__15210\,
            I => \N__15204\
        );

    \I__3433\ : CascadeBuf
    port map (
            O => \N__15207\,
            I => \N__15201\
        );

    \I__3432\ : CascadeBuf
    port map (
            O => \N__15204\,
            I => \N__15198\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__15201\,
            I => \N__15195\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__15198\,
            I => \N__15192\
        );

    \I__3429\ : CascadeBuf
    port map (
            O => \N__15195\,
            I => \N__15189\
        );

    \I__3428\ : CascadeBuf
    port map (
            O => \N__15192\,
            I => \N__15186\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__15189\,
            I => \N__15183\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__15186\,
            I => \N__15180\
        );

    \I__3425\ : CascadeBuf
    port map (
            O => \N__15183\,
            I => \N__15177\
        );

    \I__3424\ : CascadeBuf
    port map (
            O => \N__15180\,
            I => \N__15174\
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__15177\,
            I => \N__15171\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__15174\,
            I => \N__15168\
        );

    \I__3421\ : CascadeBuf
    port map (
            O => \N__15171\,
            I => \N__15165\
        );

    \I__3420\ : CascadeBuf
    port map (
            O => \N__15168\,
            I => \N__15162\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__15165\,
            I => \N__15159\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__15162\,
            I => \N__15156\
        );

    \I__3417\ : CascadeBuf
    port map (
            O => \N__15159\,
            I => \N__15153\
        );

    \I__3416\ : CascadeBuf
    port map (
            O => \N__15156\,
            I => \N__15150\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__15153\,
            I => \N__15147\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__15150\,
            I => \N__15144\
        );

    \I__3413\ : CascadeBuf
    port map (
            O => \N__15147\,
            I => \N__15141\
        );

    \I__3412\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15138\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__15141\,
            I => \N__15135\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__15138\,
            I => \N__15132\
        );

    \I__3409\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15129\
        );

    \I__3408\ : Span4Mux_s3_v
    port map (
            O => \N__15132\,
            I => \N__15126\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__15129\,
            I => \N__15123\
        );

    \I__3406\ : Sp12to4
    port map (
            O => \N__15126\,
            I => \N__15120\
        );

    \I__3405\ : Span12Mux_s5_v
    port map (
            O => \N__15123\,
            I => \N__15115\
        );

    \I__3404\ : Span12Mux_h
    port map (
            O => \N__15120\,
            I => \N__15112\
        );

    \I__3403\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15109\
        );

    \I__3402\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15106\
        );

    \I__3401\ : Span12Mux_v
    port map (
            O => \N__15115\,
            I => \N__15103\
        );

    \I__3400\ : Span12Mux_v
    port map (
            O => \N__15112\,
            I => \N__15100\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__15109\,
            I => \RX_ADDR_2\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__15106\,
            I => \RX_ADDR_2\
        );

    \I__3397\ : Odrv12
    port map (
            O => \N__15103\,
            I => \RX_ADDR_2\
        );

    \I__3396\ : Odrv12
    port map (
            O => \N__15100\,
            I => \RX_ADDR_2\
        );

    \I__3395\ : InMux
    port map (
            O => \N__15091\,
            I => \N__15088\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__15088\,
            I => \receive_module.n135\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__15085\,
            I => \N__15081\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__15084\,
            I => \N__15078\
        );

    \I__3391\ : CascadeBuf
    port map (
            O => \N__15081\,
            I => \N__15075\
        );

    \I__3390\ : CascadeBuf
    port map (
            O => \N__15078\,
            I => \N__15072\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__15075\,
            I => \N__15069\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__15072\,
            I => \N__15066\
        );

    \I__3387\ : CascadeBuf
    port map (
            O => \N__15069\,
            I => \N__15063\
        );

    \I__3386\ : CascadeBuf
    port map (
            O => \N__15066\,
            I => \N__15060\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__15063\,
            I => \N__15057\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__15060\,
            I => \N__15054\
        );

    \I__3383\ : CascadeBuf
    port map (
            O => \N__15057\,
            I => \N__15051\
        );

    \I__3382\ : CascadeBuf
    port map (
            O => \N__15054\,
            I => \N__15048\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__15051\,
            I => \N__15045\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__15048\,
            I => \N__15042\
        );

    \I__3379\ : CascadeBuf
    port map (
            O => \N__15045\,
            I => \N__15039\
        );

    \I__3378\ : CascadeBuf
    port map (
            O => \N__15042\,
            I => \N__15036\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__15039\,
            I => \N__15033\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__15036\,
            I => \N__15030\
        );

    \I__3375\ : CascadeBuf
    port map (
            O => \N__15033\,
            I => \N__15027\
        );

    \I__3374\ : CascadeBuf
    port map (
            O => \N__15030\,
            I => \N__15024\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__15027\,
            I => \N__15021\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__15024\,
            I => \N__15018\
        );

    \I__3371\ : CascadeBuf
    port map (
            O => \N__15021\,
            I => \N__15015\
        );

    \I__3370\ : CascadeBuf
    port map (
            O => \N__15018\,
            I => \N__15012\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__15015\,
            I => \N__15009\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__15012\,
            I => \N__15006\
        );

    \I__3367\ : CascadeBuf
    port map (
            O => \N__15009\,
            I => \N__15003\
        );

    \I__3366\ : CascadeBuf
    port map (
            O => \N__15006\,
            I => \N__15000\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__15003\,
            I => \N__14997\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__15000\,
            I => \N__14994\
        );

    \I__3363\ : CascadeBuf
    port map (
            O => \N__14997\,
            I => \N__14991\
        );

    \I__3362\ : CascadeBuf
    port map (
            O => \N__14994\,
            I => \N__14988\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__14991\,
            I => \N__14985\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__14988\,
            I => \N__14982\
        );

    \I__3359\ : CascadeBuf
    port map (
            O => \N__14985\,
            I => \N__14979\
        );

    \I__3358\ : CascadeBuf
    port map (
            O => \N__14982\,
            I => \N__14976\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__14979\,
            I => \N__14973\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__14976\,
            I => \N__14970\
        );

    \I__3355\ : CascadeBuf
    port map (
            O => \N__14973\,
            I => \N__14967\
        );

    \I__3354\ : CascadeBuf
    port map (
            O => \N__14970\,
            I => \N__14964\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__14967\,
            I => \N__14961\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__14964\,
            I => \N__14958\
        );

    \I__3351\ : CascadeBuf
    port map (
            O => \N__14961\,
            I => \N__14955\
        );

    \I__3350\ : CascadeBuf
    port map (
            O => \N__14958\,
            I => \N__14952\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__14955\,
            I => \N__14949\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__14952\,
            I => \N__14946\
        );

    \I__3347\ : CascadeBuf
    port map (
            O => \N__14949\,
            I => \N__14943\
        );

    \I__3346\ : CascadeBuf
    port map (
            O => \N__14946\,
            I => \N__14940\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__14943\,
            I => \N__14937\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__14940\,
            I => \N__14934\
        );

    \I__3343\ : CascadeBuf
    port map (
            O => \N__14937\,
            I => \N__14931\
        );

    \I__3342\ : CascadeBuf
    port map (
            O => \N__14934\,
            I => \N__14928\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__14931\,
            I => \N__14925\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__14928\,
            I => \N__14922\
        );

    \I__3339\ : CascadeBuf
    port map (
            O => \N__14925\,
            I => \N__14919\
        );

    \I__3338\ : CascadeBuf
    port map (
            O => \N__14922\,
            I => \N__14916\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__14919\,
            I => \N__14913\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__14916\,
            I => \N__14910\
        );

    \I__3335\ : CascadeBuf
    port map (
            O => \N__14913\,
            I => \N__14907\
        );

    \I__3334\ : CascadeBuf
    port map (
            O => \N__14910\,
            I => \N__14904\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__14907\,
            I => \N__14901\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__14904\,
            I => \N__14898\
        );

    \I__3331\ : InMux
    port map (
            O => \N__14901\,
            I => \N__14895\
        );

    \I__3330\ : InMux
    port map (
            O => \N__14898\,
            I => \N__14892\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__14895\,
            I => \N__14889\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__14892\,
            I => \N__14886\
        );

    \I__3327\ : Span4Mux_h
    port map (
            O => \N__14889\,
            I => \N__14883\
        );

    \I__3326\ : Span4Mux_h
    port map (
            O => \N__14886\,
            I => \N__14880\
        );

    \I__3325\ : Sp12to4
    port map (
            O => \N__14883\,
            I => \N__14877\
        );

    \I__3324\ : Sp12to4
    port map (
            O => \N__14880\,
            I => \N__14874\
        );

    \I__3323\ : Span12Mux_s5_v
    port map (
            O => \N__14877\,
            I => \N__14869\
        );

    \I__3322\ : Span12Mux_s5_v
    port map (
            O => \N__14874\,
            I => \N__14866\
        );

    \I__3321\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14863\
        );

    \I__3320\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14860\
        );

    \I__3319\ : Span12Mux_v
    port map (
            O => \N__14869\,
            I => \N__14855\
        );

    \I__3318\ : Span12Mux_v
    port map (
            O => \N__14866\,
            I => \N__14855\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__14863\,
            I => \RX_ADDR_1\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__14860\,
            I => \RX_ADDR_1\
        );

    \I__3315\ : Odrv12
    port map (
            O => \N__14855\,
            I => \RX_ADDR_1\
        );

    \I__3314\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14845\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__14845\,
            I => \N__14842\
        );

    \I__3312\ : Span4Mux_h
    port map (
            O => \N__14842\,
            I => \N__14839\
        );

    \I__3311\ : Span4Mux_h
    port map (
            O => \N__14839\,
            I => \N__14836\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__14836\,
            I => \line_buffer.n628\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__14833\,
            I => \N__14830\
        );

    \I__3308\ : InMux
    port map (
            O => \N__14830\,
            I => \N__14827\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__14827\,
            I => \N__14824\
        );

    \I__3306\ : Span12Mux_h
    port map (
            O => \N__14824\,
            I => \N__14821\
        );

    \I__3305\ : Span12Mux_v
    port map (
            O => \N__14821\,
            I => \N__14818\
        );

    \I__3304\ : Odrv12
    port map (
            O => \N__14818\,
            I => \line_buffer.n620\
        );

    \I__3303\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14812\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__14812\,
            I => \N__14809\
        );

    \I__3301\ : Odrv12
    port map (
            O => \N__14809\,
            I => \line_buffer.n3149\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__14806\,
            I => \line_buffer.n3152_cascade_\
        );

    \I__3299\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14800\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__14800\,
            I => \N__14797\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__14797\,
            I => \N__14794\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__14794\,
            I => \TX_DATA_5\
        );

    \I__3295\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14788\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__14788\,
            I => \N__14785\
        );

    \I__3293\ : Span12Mux_v
    port map (
            O => \N__14785\,
            I => \N__14782\
        );

    \I__3292\ : Odrv12
    port map (
            O => \N__14782\,
            I => \line_buffer.n692\
        );

    \I__3291\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14776\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__14776\,
            I => \N__14773\
        );

    \I__3289\ : Span4Mux_v
    port map (
            O => \N__14773\,
            I => \N__14770\
        );

    \I__3288\ : Span4Mux_h
    port map (
            O => \N__14770\,
            I => \N__14767\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__14767\,
            I => \line_buffer.n684\
        );

    \I__3286\ : InMux
    port map (
            O => \N__14764\,
            I => \N__14761\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__14761\,
            I => \N__14758\
        );

    \I__3284\ : Span4Mux_v
    port map (
            O => \N__14758\,
            I => \N__14755\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__14755\,
            I => \line_buffer.n3024\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__14752\,
            I => \line_buffer.n3131_cascade_\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__14749\,
            I => \N__14745\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__14748\,
            I => \N__14742\
        );

    \I__3279\ : CascadeBuf
    port map (
            O => \N__14745\,
            I => \N__14739\
        );

    \I__3278\ : CascadeBuf
    port map (
            O => \N__14742\,
            I => \N__14736\
        );

    \I__3277\ : CascadeMux
    port map (
            O => \N__14739\,
            I => \N__14733\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__14736\,
            I => \N__14730\
        );

    \I__3275\ : CascadeBuf
    port map (
            O => \N__14733\,
            I => \N__14727\
        );

    \I__3274\ : CascadeBuf
    port map (
            O => \N__14730\,
            I => \N__14724\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__14727\,
            I => \N__14721\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__14724\,
            I => \N__14718\
        );

    \I__3271\ : CascadeBuf
    port map (
            O => \N__14721\,
            I => \N__14715\
        );

    \I__3270\ : CascadeBuf
    port map (
            O => \N__14718\,
            I => \N__14712\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__14715\,
            I => \N__14709\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__14712\,
            I => \N__14706\
        );

    \I__3267\ : CascadeBuf
    port map (
            O => \N__14709\,
            I => \N__14703\
        );

    \I__3266\ : CascadeBuf
    port map (
            O => \N__14706\,
            I => \N__14700\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__14703\,
            I => \N__14697\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__14700\,
            I => \N__14694\
        );

    \I__3263\ : CascadeBuf
    port map (
            O => \N__14697\,
            I => \N__14691\
        );

    \I__3262\ : CascadeBuf
    port map (
            O => \N__14694\,
            I => \N__14688\
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__14691\,
            I => \N__14685\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__14688\,
            I => \N__14682\
        );

    \I__3259\ : CascadeBuf
    port map (
            O => \N__14685\,
            I => \N__14679\
        );

    \I__3258\ : CascadeBuf
    port map (
            O => \N__14682\,
            I => \N__14676\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__14679\,
            I => \N__14673\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__14676\,
            I => \N__14670\
        );

    \I__3255\ : CascadeBuf
    port map (
            O => \N__14673\,
            I => \N__14667\
        );

    \I__3254\ : CascadeBuf
    port map (
            O => \N__14670\,
            I => \N__14664\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__14667\,
            I => \N__14661\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__14664\,
            I => \N__14658\
        );

    \I__3251\ : CascadeBuf
    port map (
            O => \N__14661\,
            I => \N__14655\
        );

    \I__3250\ : CascadeBuf
    port map (
            O => \N__14658\,
            I => \N__14652\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__14655\,
            I => \N__14649\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__14652\,
            I => \N__14646\
        );

    \I__3247\ : CascadeBuf
    port map (
            O => \N__14649\,
            I => \N__14643\
        );

    \I__3246\ : CascadeBuf
    port map (
            O => \N__14646\,
            I => \N__14640\
        );

    \I__3245\ : CascadeMux
    port map (
            O => \N__14643\,
            I => \N__14637\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__14640\,
            I => \N__14634\
        );

    \I__3243\ : CascadeBuf
    port map (
            O => \N__14637\,
            I => \N__14631\
        );

    \I__3242\ : CascadeBuf
    port map (
            O => \N__14634\,
            I => \N__14628\
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__14631\,
            I => \N__14625\
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__14628\,
            I => \N__14622\
        );

    \I__3239\ : CascadeBuf
    port map (
            O => \N__14625\,
            I => \N__14619\
        );

    \I__3238\ : CascadeBuf
    port map (
            O => \N__14622\,
            I => \N__14616\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__14619\,
            I => \N__14613\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__14616\,
            I => \N__14610\
        );

    \I__3235\ : CascadeBuf
    port map (
            O => \N__14613\,
            I => \N__14607\
        );

    \I__3234\ : CascadeBuf
    port map (
            O => \N__14610\,
            I => \N__14604\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__14607\,
            I => \N__14601\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__14604\,
            I => \N__14598\
        );

    \I__3231\ : CascadeBuf
    port map (
            O => \N__14601\,
            I => \N__14595\
        );

    \I__3230\ : CascadeBuf
    port map (
            O => \N__14598\,
            I => \N__14592\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__14595\,
            I => \N__14589\
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__14592\,
            I => \N__14586\
        );

    \I__3227\ : CascadeBuf
    port map (
            O => \N__14589\,
            I => \N__14583\
        );

    \I__3226\ : CascadeBuf
    port map (
            O => \N__14586\,
            I => \N__14580\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__14583\,
            I => \N__14577\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__14580\,
            I => \N__14574\
        );

    \I__3223\ : CascadeBuf
    port map (
            O => \N__14577\,
            I => \N__14571\
        );

    \I__3222\ : CascadeBuf
    port map (
            O => \N__14574\,
            I => \N__14568\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__14571\,
            I => \N__14565\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__14568\,
            I => \N__14562\
        );

    \I__3219\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14559\
        );

    \I__3218\ : InMux
    port map (
            O => \N__14562\,
            I => \N__14556\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__14559\,
            I => \N__14553\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__14556\,
            I => \N__14550\
        );

    \I__3215\ : Span4Mux_s1_v
    port map (
            O => \N__14553\,
            I => \N__14547\
        );

    \I__3214\ : Span4Mux_s1_v
    port map (
            O => \N__14550\,
            I => \N__14544\
        );

    \I__3213\ : Span4Mux_v
    port map (
            O => \N__14547\,
            I => \N__14541\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__14544\,
            I => \N__14538\
        );

    \I__3211\ : Sp12to4
    port map (
            O => \N__14541\,
            I => \N__14535\
        );

    \I__3210\ : Sp12to4
    port map (
            O => \N__14538\,
            I => \N__14532\
        );

    \I__3209\ : Span12Mux_s9_h
    port map (
            O => \N__14535\,
            I => \N__14527\
        );

    \I__3208\ : Span12Mux_s10_h
    port map (
            O => \N__14532\,
            I => \N__14524\
        );

    \I__3207\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14521\
        );

    \I__3206\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14518\
        );

    \I__3205\ : Span12Mux_v
    port map (
            O => \N__14527\,
            I => \N__14513\
        );

    \I__3204\ : Span12Mux_v
    port map (
            O => \N__14524\,
            I => \N__14513\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__14521\,
            I => \RX_ADDR_9\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__14518\,
            I => \RX_ADDR_9\
        );

    \I__3201\ : Odrv12
    port map (
            O => \N__14513\,
            I => \RX_ADDR_9\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__14506\,
            I => \N__14503\
        );

    \I__3199\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14500\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__14500\,
            I => \receive_module.n127\
        );

    \I__3197\ : InMux
    port map (
            O => \N__14497\,
            I => \receive_module.n2735\
        );

    \I__3196\ : InMux
    port map (
            O => \N__14494\,
            I => \receive_module.n2736\
        );

    \I__3195\ : InMux
    port map (
            O => \N__14491\,
            I => \receive_module.n2737\
        );

    \I__3194\ : InMux
    port map (
            O => \N__14488\,
            I => \receive_module.n2738\
        );

    \I__3193\ : InMux
    port map (
            O => \N__14485\,
            I => \receive_module.n2739\
        );

    \I__3192\ : CEMux
    port map (
            O => \N__14482\,
            I => \N__14479\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__14479\,
            I => \N__14476\
        );

    \I__3190\ : Span4Mux_v
    port map (
            O => \N__14476\,
            I => \N__14473\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__14473\,
            I => \receive_module.n3181\
        );

    \I__3188\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14467\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__14467\,
            I => \N__14463\
        );

    \I__3186\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14460\
        );

    \I__3185\ : Span4Mux_h
    port map (
            O => \N__14463\,
            I => \N__14457\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__14460\,
            I => \transmit_module.n388\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__14457\,
            I => \transmit_module.n388\
        );

    \I__3182\ : IoInMux
    port map (
            O => \N__14452\,
            I => \N__14449\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__14449\,
            I => \N__14446\
        );

    \I__3180\ : IoSpan4Mux
    port map (
            O => \N__14446\,
            I => \N__14437\
        );

    \I__3179\ : SRMux
    port map (
            O => \N__14445\,
            I => \N__14431\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__14444\,
            I => \N__14428\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__14443\,
            I => \N__14420\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__14442\,
            I => \N__14417\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__14441\,
            I => \N__14414\
        );

    \I__3174\ : SRMux
    port map (
            O => \N__14440\,
            I => \N__14408\
        );

    \I__3173\ : Span4Mux_s3_h
    port map (
            O => \N__14437\,
            I => \N__14405\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__14436\,
            I => \N__14399\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__14435\,
            I => \N__14394\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__14434\,
            I => \N__14391\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__14431\,
            I => \N__14388\
        );

    \I__3168\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14385\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__14427\,
            I => \N__14381\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__14426\,
            I => \N__14378\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__14425\,
            I => \N__14375\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__14424\,
            I => \N__14372\
        );

    \I__3163\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14369\
        );

    \I__3162\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14362\
        );

    \I__3161\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14362\
        );

    \I__3160\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14362\
        );

    \I__3159\ : SRMux
    port map (
            O => \N__14413\,
            I => \N__14357\
        );

    \I__3158\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14352\
        );

    \I__3157\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14352\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__14408\,
            I => \N__14349\
        );

    \I__3155\ : Span4Mux_h
    port map (
            O => \N__14405\,
            I => \N__14345\
        );

    \I__3154\ : SRMux
    port map (
            O => \N__14404\,
            I => \N__14342\
        );

    \I__3153\ : InMux
    port map (
            O => \N__14403\,
            I => \N__14335\
        );

    \I__3152\ : InMux
    port map (
            O => \N__14402\,
            I => \N__14335\
        );

    \I__3151\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14335\
        );

    \I__3150\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14332\
        );

    \I__3149\ : InMux
    port map (
            O => \N__14397\,
            I => \N__14325\
        );

    \I__3148\ : InMux
    port map (
            O => \N__14394\,
            I => \N__14325\
        );

    \I__3147\ : InMux
    port map (
            O => \N__14391\,
            I => \N__14325\
        );

    \I__3146\ : Span4Mux_v
    port map (
            O => \N__14388\,
            I => \N__14320\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__14385\,
            I => \N__14320\
        );

    \I__3144\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14311\
        );

    \I__3143\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14311\
        );

    \I__3142\ : InMux
    port map (
            O => \N__14378\,
            I => \N__14311\
        );

    \I__3141\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14311\
        );

    \I__3140\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14308\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__14369\,
            I => \N__14303\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__14362\,
            I => \N__14303\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__14361\,
            I => \N__14300\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__14360\,
            I => \N__14297\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14293\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__14352\,
            I => \N__14290\
        );

    \I__3133\ : Span4Mux_v
    port map (
            O => \N__14349\,
            I => \N__14287\
        );

    \I__3132\ : InMux
    port map (
            O => \N__14348\,
            I => \N__14284\
        );

    \I__3131\ : Span4Mux_h
    port map (
            O => \N__14345\,
            I => \N__14279\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14279\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__14335\,
            I => \N__14264\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__14332\,
            I => \N__14264\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__14325\,
            I => \N__14264\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__14320\,
            I => \N__14264\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__14311\,
            I => \N__14264\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__14308\,
            I => \N__14264\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__14303\,
            I => \N__14264\
        );

    \I__3122\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14257\
        );

    \I__3121\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14257\
        );

    \I__3120\ : InMux
    port map (
            O => \N__14296\,
            I => \N__14257\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__14293\,
            I => \N__14254\
        );

    \I__3118\ : Span4Mux_v
    port map (
            O => \N__14290\,
            I => \N__14247\
        );

    \I__3117\ : Span4Mux_h
    port map (
            O => \N__14287\,
            I => \N__14247\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14247\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__14279\,
            I => \N__14242\
        );

    \I__3114\ : Span4Mux_v
    port map (
            O => \N__14264\,
            I => \N__14242\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__14257\,
            I => \ADV_VSYNC_c\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__14254\,
            I => \ADV_VSYNC_c\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__14247\,
            I => \ADV_VSYNC_c\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__14242\,
            I => \ADV_VSYNC_c\
        );

    \I__3109\ : IoInMux
    port map (
            O => \N__14233\,
            I => \N__14230\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__14230\,
            I => \N__14226\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__14229\,
            I => \N__14223\
        );

    \I__3106\ : Span12Mux_s3_h
    port map (
            O => \N__14226\,
            I => \N__14220\
        );

    \I__3105\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14216\
        );

    \I__3104\ : Span12Mux_h
    port map (
            O => \N__14220\,
            I => \N__14213\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__14219\,
            I => \N__14210\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__14216\,
            I => \N__14207\
        );

    \I__3101\ : Span12Mux_v
    port map (
            O => \N__14213\,
            I => \N__14203\
        );

    \I__3100\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14200\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__14207\,
            I => \N__14197\
        );

    \I__3098\ : InMux
    port map (
            O => \N__14206\,
            I => \N__14194\
        );

    \I__3097\ : Odrv12
    port map (
            O => \N__14203\,
            I => \DEBUG_c_0\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__14200\,
            I => \DEBUG_c_0\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__14197\,
            I => \DEBUG_c_0\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__14194\,
            I => \DEBUG_c_0\
        );

    \I__3093\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14168\
        );

    \I__3092\ : SRMux
    port map (
            O => \N__14184\,
            I => \N__14161\
        );

    \I__3091\ : InMux
    port map (
            O => \N__14183\,
            I => \N__14158\
        );

    \I__3090\ : InMux
    port map (
            O => \N__14182\,
            I => \N__14149\
        );

    \I__3089\ : InMux
    port map (
            O => \N__14181\,
            I => \N__14149\
        );

    \I__3088\ : InMux
    port map (
            O => \N__14180\,
            I => \N__14149\
        );

    \I__3087\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14149\
        );

    \I__3086\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14142\
        );

    \I__3085\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14142\
        );

    \I__3084\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14142\
        );

    \I__3083\ : InMux
    port map (
            O => \N__14175\,
            I => \N__14132\
        );

    \I__3082\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14132\
        );

    \I__3081\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14132\
        );

    \I__3080\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14125\
        );

    \I__3079\ : InMux
    port map (
            O => \N__14171\,
            I => \N__14125\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__14168\,
            I => \N__14122\
        );

    \I__3077\ : InMux
    port map (
            O => \N__14167\,
            I => \N__14113\
        );

    \I__3076\ : InMux
    port map (
            O => \N__14166\,
            I => \N__14113\
        );

    \I__3075\ : InMux
    port map (
            O => \N__14165\,
            I => \N__14113\
        );

    \I__3074\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14113\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__14161\,
            I => \N__14110\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__14158\,
            I => \N__14103\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__14149\,
            I => \N__14103\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__14142\,
            I => \N__14103\
        );

    \I__3069\ : InMux
    port map (
            O => \N__14141\,
            I => \N__14096\
        );

    \I__3068\ : InMux
    port map (
            O => \N__14140\,
            I => \N__14096\
        );

    \I__3067\ : InMux
    port map (
            O => \N__14139\,
            I => \N__14093\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__14132\,
            I => \N__14090\
        );

    \I__3065\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14087\
        );

    \I__3064\ : SRMux
    port map (
            O => \N__14130\,
            I => \N__14084\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__14125\,
            I => \N__14073\
        );

    \I__3062\ : Span4Mux_v
    port map (
            O => \N__14122\,
            I => \N__14073\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__14113\,
            I => \N__14073\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__14110\,
            I => \N__14073\
        );

    \I__3059\ : Span4Mux_h
    port map (
            O => \N__14103\,
            I => \N__14073\
        );

    \I__3058\ : SRMux
    port map (
            O => \N__14102\,
            I => \N__14070\
        );

    \I__3057\ : SRMux
    port map (
            O => \N__14101\,
            I => \N__14067\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__14096\,
            I => \VGA_VISIBLE\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__14093\,
            I => \VGA_VISIBLE\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__14090\,
            I => \VGA_VISIBLE\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__14087\,
            I => \VGA_VISIBLE\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__14084\,
            I => \VGA_VISIBLE\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__14073\,
            I => \VGA_VISIBLE\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__14070\,
            I => \VGA_VISIBLE\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__14067\,
            I => \VGA_VISIBLE\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__14050\,
            I => \N__14046\
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__14049\,
            I => \N__14043\
        );

    \I__3046\ : CascadeBuf
    port map (
            O => \N__14046\,
            I => \N__14040\
        );

    \I__3045\ : CascadeBuf
    port map (
            O => \N__14043\,
            I => \N__14037\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__14040\,
            I => \N__14034\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__14037\,
            I => \N__14031\
        );

    \I__3042\ : CascadeBuf
    port map (
            O => \N__14034\,
            I => \N__14028\
        );

    \I__3041\ : CascadeBuf
    port map (
            O => \N__14031\,
            I => \N__14025\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__14028\,
            I => \N__14022\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__14025\,
            I => \N__14019\
        );

    \I__3038\ : CascadeBuf
    port map (
            O => \N__14022\,
            I => \N__14016\
        );

    \I__3037\ : CascadeBuf
    port map (
            O => \N__14019\,
            I => \N__14013\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__14016\,
            I => \N__14010\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__14013\,
            I => \N__14007\
        );

    \I__3034\ : CascadeBuf
    port map (
            O => \N__14010\,
            I => \N__14004\
        );

    \I__3033\ : CascadeBuf
    port map (
            O => \N__14007\,
            I => \N__14001\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__14004\,
            I => \N__13998\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__14001\,
            I => \N__13995\
        );

    \I__3030\ : CascadeBuf
    port map (
            O => \N__13998\,
            I => \N__13992\
        );

    \I__3029\ : CascadeBuf
    port map (
            O => \N__13995\,
            I => \N__13989\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__13992\,
            I => \N__13986\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__13989\,
            I => \N__13983\
        );

    \I__3026\ : CascadeBuf
    port map (
            O => \N__13986\,
            I => \N__13980\
        );

    \I__3025\ : CascadeBuf
    port map (
            O => \N__13983\,
            I => \N__13977\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__13980\,
            I => \N__13974\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__13977\,
            I => \N__13971\
        );

    \I__3022\ : CascadeBuf
    port map (
            O => \N__13974\,
            I => \N__13968\
        );

    \I__3021\ : CascadeBuf
    port map (
            O => \N__13971\,
            I => \N__13965\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__13968\,
            I => \N__13962\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__13965\,
            I => \N__13959\
        );

    \I__3018\ : CascadeBuf
    port map (
            O => \N__13962\,
            I => \N__13956\
        );

    \I__3017\ : CascadeBuf
    port map (
            O => \N__13959\,
            I => \N__13953\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__13956\,
            I => \N__13950\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__13953\,
            I => \N__13947\
        );

    \I__3014\ : CascadeBuf
    port map (
            O => \N__13950\,
            I => \N__13944\
        );

    \I__3013\ : CascadeBuf
    port map (
            O => \N__13947\,
            I => \N__13941\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__13944\,
            I => \N__13938\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__13941\,
            I => \N__13935\
        );

    \I__3010\ : CascadeBuf
    port map (
            O => \N__13938\,
            I => \N__13932\
        );

    \I__3009\ : CascadeBuf
    port map (
            O => \N__13935\,
            I => \N__13929\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__13932\,
            I => \N__13926\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__13929\,
            I => \N__13923\
        );

    \I__3006\ : CascadeBuf
    port map (
            O => \N__13926\,
            I => \N__13920\
        );

    \I__3005\ : CascadeBuf
    port map (
            O => \N__13923\,
            I => \N__13917\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__13920\,
            I => \N__13914\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__13917\,
            I => \N__13911\
        );

    \I__3002\ : CascadeBuf
    port map (
            O => \N__13914\,
            I => \N__13908\
        );

    \I__3001\ : CascadeBuf
    port map (
            O => \N__13911\,
            I => \N__13905\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__13908\,
            I => \N__13902\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__13905\,
            I => \N__13899\
        );

    \I__2998\ : CascadeBuf
    port map (
            O => \N__13902\,
            I => \N__13896\
        );

    \I__2997\ : CascadeBuf
    port map (
            O => \N__13899\,
            I => \N__13893\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__13896\,
            I => \N__13890\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__13893\,
            I => \N__13887\
        );

    \I__2994\ : CascadeBuf
    port map (
            O => \N__13890\,
            I => \N__13884\
        );

    \I__2993\ : CascadeBuf
    port map (
            O => \N__13887\,
            I => \N__13881\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__13884\,
            I => \N__13878\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__13881\,
            I => \N__13875\
        );

    \I__2990\ : CascadeBuf
    port map (
            O => \N__13878\,
            I => \N__13872\
        );

    \I__2989\ : CascadeBuf
    port map (
            O => \N__13875\,
            I => \N__13869\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__13872\,
            I => \N__13866\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__13869\,
            I => \N__13863\
        );

    \I__2986\ : InMux
    port map (
            O => \N__13866\,
            I => \N__13860\
        );

    \I__2985\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13857\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__13860\,
            I => \N__13854\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__13857\,
            I => \N__13851\
        );

    \I__2982\ : Span12Mux_h
    port map (
            O => \N__13854\,
            I => \N__13848\
        );

    \I__2981\ : Span12Mux_s11_h
    port map (
            O => \N__13851\,
            I => \N__13845\
        );

    \I__2980\ : Span12Mux_v
    port map (
            O => \N__13848\,
            I => \N__13842\
        );

    \I__2979\ : Span12Mux_v
    port map (
            O => \N__13845\,
            I => \N__13839\
        );

    \I__2978\ : Odrv12
    port map (
            O => \N__13842\,
            I => n28
        );

    \I__2977\ : Odrv12
    port map (
            O => \N__13839\,
            I => n28
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__13834\,
            I => \N__13831\
        );

    \I__2975\ : InMux
    port map (
            O => \N__13831\,
            I => \N__13828\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__13828\,
            I => \N__13825\
        );

    \I__2973\ : Span4Mux_v
    port map (
            O => \N__13825\,
            I => \N__13822\
        );

    \I__2972\ : Sp12to4
    port map (
            O => \N__13822\,
            I => \N__13819\
        );

    \I__2971\ : Span12Mux_h
    port map (
            O => \N__13819\,
            I => \N__13816\
        );

    \I__2970\ : Span12Mux_v
    port map (
            O => \N__13816\,
            I => \N__13813\
        );

    \I__2969\ : Odrv12
    port map (
            O => \N__13813\,
            I => \line_buffer.n744\
        );

    \I__2968\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13807\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__13807\,
            I => \N__13804\
        );

    \I__2966\ : Span4Mux_v
    port map (
            O => \N__13804\,
            I => \N__13801\
        );

    \I__2965\ : Sp12to4
    port map (
            O => \N__13801\,
            I => \N__13798\
        );

    \I__2964\ : Odrv12
    port map (
            O => \N__13798\,
            I => \line_buffer.n752\
        );

    \I__2963\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13792\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__13792\,
            I => \N__13789\
        );

    \I__2961\ : Span4Mux_v
    port map (
            O => \N__13789\,
            I => \N__13786\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__13786\,
            I => \line_buffer.n3119\
        );

    \I__2959\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13780\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__13780\,
            I => \N__13777\
        );

    \I__2957\ : Odrv12
    port map (
            O => \N__13777\,
            I => \line_buffer.n695\
        );

    \I__2956\ : InMux
    port map (
            O => \N__13774\,
            I => \N__13771\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__13771\,
            I => \N__13768\
        );

    \I__2954\ : Span4Mux_h
    port map (
            O => \N__13768\,
            I => \N__13765\
        );

    \I__2953\ : Sp12to4
    port map (
            O => \N__13765\,
            I => \N__13762\
        );

    \I__2952\ : Span12Mux_v
    port map (
            O => \N__13762\,
            I => \N__13759\
        );

    \I__2951\ : Span12Mux_v
    port map (
            O => \N__13759\,
            I => \N__13756\
        );

    \I__2950\ : Odrv12
    port map (
            O => \N__13756\,
            I => \line_buffer.n687\
        );

    \I__2949\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13750\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__13750\,
            I => \line_buffer.n3027\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__13747\,
            I => \N__13743\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__13746\,
            I => \N__13740\
        );

    \I__2945\ : CascadeBuf
    port map (
            O => \N__13743\,
            I => \N__13737\
        );

    \I__2944\ : CascadeBuf
    port map (
            O => \N__13740\,
            I => \N__13734\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__13737\,
            I => \N__13731\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__13734\,
            I => \N__13728\
        );

    \I__2941\ : CascadeBuf
    port map (
            O => \N__13731\,
            I => \N__13725\
        );

    \I__2940\ : CascadeBuf
    port map (
            O => \N__13728\,
            I => \N__13722\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__13725\,
            I => \N__13719\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__13722\,
            I => \N__13716\
        );

    \I__2937\ : CascadeBuf
    port map (
            O => \N__13719\,
            I => \N__13713\
        );

    \I__2936\ : CascadeBuf
    port map (
            O => \N__13716\,
            I => \N__13710\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__13713\,
            I => \N__13707\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__13710\,
            I => \N__13704\
        );

    \I__2933\ : CascadeBuf
    port map (
            O => \N__13707\,
            I => \N__13701\
        );

    \I__2932\ : CascadeBuf
    port map (
            O => \N__13704\,
            I => \N__13698\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__13701\,
            I => \N__13695\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__13698\,
            I => \N__13692\
        );

    \I__2929\ : CascadeBuf
    port map (
            O => \N__13695\,
            I => \N__13689\
        );

    \I__2928\ : CascadeBuf
    port map (
            O => \N__13692\,
            I => \N__13686\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__13689\,
            I => \N__13683\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__13686\,
            I => \N__13680\
        );

    \I__2925\ : CascadeBuf
    port map (
            O => \N__13683\,
            I => \N__13677\
        );

    \I__2924\ : CascadeBuf
    port map (
            O => \N__13680\,
            I => \N__13674\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__13677\,
            I => \N__13671\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__13674\,
            I => \N__13668\
        );

    \I__2921\ : CascadeBuf
    port map (
            O => \N__13671\,
            I => \N__13665\
        );

    \I__2920\ : CascadeBuf
    port map (
            O => \N__13668\,
            I => \N__13662\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__13665\,
            I => \N__13659\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__13662\,
            I => \N__13656\
        );

    \I__2917\ : CascadeBuf
    port map (
            O => \N__13659\,
            I => \N__13653\
        );

    \I__2916\ : CascadeBuf
    port map (
            O => \N__13656\,
            I => \N__13650\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__13653\,
            I => \N__13647\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__13650\,
            I => \N__13644\
        );

    \I__2913\ : CascadeBuf
    port map (
            O => \N__13647\,
            I => \N__13641\
        );

    \I__2912\ : CascadeBuf
    port map (
            O => \N__13644\,
            I => \N__13638\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__13641\,
            I => \N__13635\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__13638\,
            I => \N__13632\
        );

    \I__2909\ : CascadeBuf
    port map (
            O => \N__13635\,
            I => \N__13629\
        );

    \I__2908\ : CascadeBuf
    port map (
            O => \N__13632\,
            I => \N__13626\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__13629\,
            I => \N__13623\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__13626\,
            I => \N__13620\
        );

    \I__2905\ : CascadeBuf
    port map (
            O => \N__13623\,
            I => \N__13617\
        );

    \I__2904\ : CascadeBuf
    port map (
            O => \N__13620\,
            I => \N__13614\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__13617\,
            I => \N__13611\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__13614\,
            I => \N__13608\
        );

    \I__2901\ : CascadeBuf
    port map (
            O => \N__13611\,
            I => \N__13605\
        );

    \I__2900\ : CascadeBuf
    port map (
            O => \N__13608\,
            I => \N__13602\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__13605\,
            I => \N__13599\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__13602\,
            I => \N__13596\
        );

    \I__2897\ : CascadeBuf
    port map (
            O => \N__13599\,
            I => \N__13593\
        );

    \I__2896\ : CascadeBuf
    port map (
            O => \N__13596\,
            I => \N__13590\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__13593\,
            I => \N__13587\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__13590\,
            I => \N__13584\
        );

    \I__2893\ : CascadeBuf
    port map (
            O => \N__13587\,
            I => \N__13581\
        );

    \I__2892\ : CascadeBuf
    port map (
            O => \N__13584\,
            I => \N__13578\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__13581\,
            I => \N__13575\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__13578\,
            I => \N__13572\
        );

    \I__2889\ : CascadeBuf
    port map (
            O => \N__13575\,
            I => \N__13569\
        );

    \I__2888\ : CascadeBuf
    port map (
            O => \N__13572\,
            I => \N__13566\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__13569\,
            I => \N__13563\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__13566\,
            I => \N__13560\
        );

    \I__2885\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13557\
        );

    \I__2884\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13554\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__13557\,
            I => \N__13551\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__13554\,
            I => \N__13548\
        );

    \I__2881\ : Span4Mux_h
    port map (
            O => \N__13551\,
            I => \N__13545\
        );

    \I__2880\ : Sp12to4
    port map (
            O => \N__13548\,
            I => \N__13541\
        );

    \I__2879\ : Sp12to4
    port map (
            O => \N__13545\,
            I => \N__13538\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__13544\,
            I => \N__13535\
        );

    \I__2877\ : Span12Mux_s5_v
    port map (
            O => \N__13541\,
            I => \N__13531\
        );

    \I__2876\ : Span12Mux_s5_v
    port map (
            O => \N__13538\,
            I => \N__13528\
        );

    \I__2875\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13525\
        );

    \I__2874\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13522\
        );

    \I__2873\ : Span12Mux_v
    port map (
            O => \N__13531\,
            I => \N__13519\
        );

    \I__2872\ : Span12Mux_v
    port map (
            O => \N__13528\,
            I => \N__13516\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__13525\,
            I => \RX_ADDR_0\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__13522\,
            I => \RX_ADDR_0\
        );

    \I__2869\ : Odrv12
    port map (
            O => \N__13519\,
            I => \RX_ADDR_0\
        );

    \I__2868\ : Odrv12
    port map (
            O => \N__13516\,
            I => \RX_ADDR_0\
        );

    \I__2867\ : InMux
    port map (
            O => \N__13507\,
            I => \N__13504\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__13504\,
            I => \receive_module.n136\
        );

    \I__2865\ : InMux
    port map (
            O => \N__13501\,
            I => \bfn_18_14_0_\
        );

    \I__2864\ : InMux
    port map (
            O => \N__13498\,
            I => \receive_module.n2727\
        );

    \I__2863\ : InMux
    port map (
            O => \N__13495\,
            I => \receive_module.n2728\
        );

    \I__2862\ : InMux
    port map (
            O => \N__13492\,
            I => \receive_module.n2729\
        );

    \I__2861\ : InMux
    port map (
            O => \N__13489\,
            I => \receive_module.n2730\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__13486\,
            I => \N__13482\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__13485\,
            I => \N__13479\
        );

    \I__2858\ : CascadeBuf
    port map (
            O => \N__13482\,
            I => \N__13476\
        );

    \I__2857\ : CascadeBuf
    port map (
            O => \N__13479\,
            I => \N__13473\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__13476\,
            I => \N__13470\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__13473\,
            I => \N__13467\
        );

    \I__2854\ : CascadeBuf
    port map (
            O => \N__13470\,
            I => \N__13464\
        );

    \I__2853\ : CascadeBuf
    port map (
            O => \N__13467\,
            I => \N__13461\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__13464\,
            I => \N__13458\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__13461\,
            I => \N__13455\
        );

    \I__2850\ : CascadeBuf
    port map (
            O => \N__13458\,
            I => \N__13452\
        );

    \I__2849\ : CascadeBuf
    port map (
            O => \N__13455\,
            I => \N__13449\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__13452\,
            I => \N__13446\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__13449\,
            I => \N__13443\
        );

    \I__2846\ : CascadeBuf
    port map (
            O => \N__13446\,
            I => \N__13440\
        );

    \I__2845\ : CascadeBuf
    port map (
            O => \N__13443\,
            I => \N__13437\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__13440\,
            I => \N__13434\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__13437\,
            I => \N__13431\
        );

    \I__2842\ : CascadeBuf
    port map (
            O => \N__13434\,
            I => \N__13428\
        );

    \I__2841\ : CascadeBuf
    port map (
            O => \N__13431\,
            I => \N__13425\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__13428\,
            I => \N__13422\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__13425\,
            I => \N__13419\
        );

    \I__2838\ : CascadeBuf
    port map (
            O => \N__13422\,
            I => \N__13416\
        );

    \I__2837\ : CascadeBuf
    port map (
            O => \N__13419\,
            I => \N__13413\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__13416\,
            I => \N__13410\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__13413\,
            I => \N__13407\
        );

    \I__2834\ : CascadeBuf
    port map (
            O => \N__13410\,
            I => \N__13404\
        );

    \I__2833\ : CascadeBuf
    port map (
            O => \N__13407\,
            I => \N__13401\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__13404\,
            I => \N__13398\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__13401\,
            I => \N__13395\
        );

    \I__2830\ : CascadeBuf
    port map (
            O => \N__13398\,
            I => \N__13392\
        );

    \I__2829\ : CascadeBuf
    port map (
            O => \N__13395\,
            I => \N__13389\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__13392\,
            I => \N__13386\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__13389\,
            I => \N__13383\
        );

    \I__2826\ : CascadeBuf
    port map (
            O => \N__13386\,
            I => \N__13380\
        );

    \I__2825\ : CascadeBuf
    port map (
            O => \N__13383\,
            I => \N__13377\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__13380\,
            I => \N__13374\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__13377\,
            I => \N__13371\
        );

    \I__2822\ : CascadeBuf
    port map (
            O => \N__13374\,
            I => \N__13368\
        );

    \I__2821\ : CascadeBuf
    port map (
            O => \N__13371\,
            I => \N__13365\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__13368\,
            I => \N__13362\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__13365\,
            I => \N__13359\
        );

    \I__2818\ : CascadeBuf
    port map (
            O => \N__13362\,
            I => \N__13356\
        );

    \I__2817\ : CascadeBuf
    port map (
            O => \N__13359\,
            I => \N__13353\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__13356\,
            I => \N__13350\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__13353\,
            I => \N__13347\
        );

    \I__2814\ : CascadeBuf
    port map (
            O => \N__13350\,
            I => \N__13344\
        );

    \I__2813\ : CascadeBuf
    port map (
            O => \N__13347\,
            I => \N__13341\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__13344\,
            I => \N__13338\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__13341\,
            I => \N__13335\
        );

    \I__2810\ : CascadeBuf
    port map (
            O => \N__13338\,
            I => \N__13332\
        );

    \I__2809\ : CascadeBuf
    port map (
            O => \N__13335\,
            I => \N__13329\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__13332\,
            I => \N__13326\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__13329\,
            I => \N__13323\
        );

    \I__2806\ : CascadeBuf
    port map (
            O => \N__13326\,
            I => \N__13320\
        );

    \I__2805\ : CascadeBuf
    port map (
            O => \N__13323\,
            I => \N__13317\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__13320\,
            I => \N__13314\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__13317\,
            I => \N__13311\
        );

    \I__2802\ : CascadeBuf
    port map (
            O => \N__13314\,
            I => \N__13308\
        );

    \I__2801\ : CascadeBuf
    port map (
            O => \N__13311\,
            I => \N__13305\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__13308\,
            I => \N__13302\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__13305\,
            I => \N__13299\
        );

    \I__2798\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13296\
        );

    \I__2797\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13293\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__13296\,
            I => \N__13290\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__13293\,
            I => \N__13287\
        );

    \I__2794\ : Span4Mux_s1_v
    port map (
            O => \N__13290\,
            I => \N__13284\
        );

    \I__2793\ : Span4Mux_s1_v
    port map (
            O => \N__13287\,
            I => \N__13281\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__13284\,
            I => \N__13278\
        );

    \I__2791\ : Span4Mux_h
    port map (
            O => \N__13281\,
            I => \N__13275\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__13278\,
            I => \N__13269\
        );

    \I__2789\ : Span4Mux_h
    port map (
            O => \N__13275\,
            I => \N__13269\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__13274\,
            I => \N__13266\
        );

    \I__2787\ : Sp12to4
    port map (
            O => \N__13269\,
            I => \N__13262\
        );

    \I__2786\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13259\
        );

    \I__2785\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13256\
        );

    \I__2784\ : Span12Mux_s11_v
    port map (
            O => \N__13262\,
            I => \N__13253\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__13259\,
            I => \RX_ADDR_5\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__13256\,
            I => \RX_ADDR_5\
        );

    \I__2781\ : Odrv12
    port map (
            O => \N__13253\,
            I => \RX_ADDR_5\
        );

    \I__2780\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13243\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__13243\,
            I => \receive_module.n131\
        );

    \I__2778\ : InMux
    port map (
            O => \N__13240\,
            I => \receive_module.n2731\
        );

    \I__2777\ : InMux
    port map (
            O => \N__13237\,
            I => \receive_module.n2732\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__2775\ : CascadeBuf
    port map (
            O => \N__13231\,
            I => \N__13228\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__13228\,
            I => \N__13224\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__13227\,
            I => \N__13221\
        );

    \I__2772\ : CascadeBuf
    port map (
            O => \N__13224\,
            I => \N__13218\
        );

    \I__2771\ : CascadeBuf
    port map (
            O => \N__13221\,
            I => \N__13215\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__13218\,
            I => \N__13212\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__13215\,
            I => \N__13209\
        );

    \I__2768\ : CascadeBuf
    port map (
            O => \N__13212\,
            I => \N__13206\
        );

    \I__2767\ : CascadeBuf
    port map (
            O => \N__13209\,
            I => \N__13203\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__13206\,
            I => \N__13200\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__13203\,
            I => \N__13197\
        );

    \I__2764\ : CascadeBuf
    port map (
            O => \N__13200\,
            I => \N__13194\
        );

    \I__2763\ : CascadeBuf
    port map (
            O => \N__13197\,
            I => \N__13191\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__13194\,
            I => \N__13188\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__13191\,
            I => \N__13185\
        );

    \I__2760\ : CascadeBuf
    port map (
            O => \N__13188\,
            I => \N__13182\
        );

    \I__2759\ : CascadeBuf
    port map (
            O => \N__13185\,
            I => \N__13179\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__13182\,
            I => \N__13176\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__13179\,
            I => \N__13173\
        );

    \I__2756\ : CascadeBuf
    port map (
            O => \N__13176\,
            I => \N__13170\
        );

    \I__2755\ : CascadeBuf
    port map (
            O => \N__13173\,
            I => \N__13167\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__13170\,
            I => \N__13164\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__13167\,
            I => \N__13161\
        );

    \I__2752\ : CascadeBuf
    port map (
            O => \N__13164\,
            I => \N__13158\
        );

    \I__2751\ : CascadeBuf
    port map (
            O => \N__13161\,
            I => \N__13155\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__13158\,
            I => \N__13152\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__13155\,
            I => \N__13149\
        );

    \I__2748\ : CascadeBuf
    port map (
            O => \N__13152\,
            I => \N__13146\
        );

    \I__2747\ : CascadeBuf
    port map (
            O => \N__13149\,
            I => \N__13143\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__13146\,
            I => \N__13140\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__13143\,
            I => \N__13137\
        );

    \I__2744\ : CascadeBuf
    port map (
            O => \N__13140\,
            I => \N__13134\
        );

    \I__2743\ : CascadeBuf
    port map (
            O => \N__13137\,
            I => \N__13131\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__13134\,
            I => \N__13128\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__13131\,
            I => \N__13125\
        );

    \I__2740\ : CascadeBuf
    port map (
            O => \N__13128\,
            I => \N__13122\
        );

    \I__2739\ : CascadeBuf
    port map (
            O => \N__13125\,
            I => \N__13119\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__13122\,
            I => \N__13116\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__13119\,
            I => \N__13113\
        );

    \I__2736\ : CascadeBuf
    port map (
            O => \N__13116\,
            I => \N__13110\
        );

    \I__2735\ : CascadeBuf
    port map (
            O => \N__13113\,
            I => \N__13107\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__13110\,
            I => \N__13104\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__13107\,
            I => \N__13101\
        );

    \I__2732\ : CascadeBuf
    port map (
            O => \N__13104\,
            I => \N__13098\
        );

    \I__2731\ : CascadeBuf
    port map (
            O => \N__13101\,
            I => \N__13095\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__13098\,
            I => \N__13092\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__13095\,
            I => \N__13089\
        );

    \I__2728\ : CascadeBuf
    port map (
            O => \N__13092\,
            I => \N__13086\
        );

    \I__2727\ : CascadeBuf
    port map (
            O => \N__13089\,
            I => \N__13083\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__13086\,
            I => \N__13080\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__13083\,
            I => \N__13077\
        );

    \I__2724\ : CascadeBuf
    port map (
            O => \N__13080\,
            I => \N__13074\
        );

    \I__2723\ : CascadeBuf
    port map (
            O => \N__13077\,
            I => \N__13071\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__13074\,
            I => \N__13068\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__13071\,
            I => \N__13065\
        );

    \I__2720\ : CascadeBuf
    port map (
            O => \N__13068\,
            I => \N__13062\
        );

    \I__2719\ : CascadeBuf
    port map (
            O => \N__13065\,
            I => \N__13059\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__13062\,
            I => \N__13056\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__13059\,
            I => \N__13053\
        );

    \I__2716\ : InMux
    port map (
            O => \N__13056\,
            I => \N__13050\
        );

    \I__2715\ : CascadeBuf
    port map (
            O => \N__13053\,
            I => \N__13047\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__13050\,
            I => \N__13044\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__13047\,
            I => \N__13041\
        );

    \I__2712\ : Span4Mux_s1_v
    port map (
            O => \N__13044\,
            I => \N__13038\
        );

    \I__2711\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13035\
        );

    \I__2710\ : Span4Mux_h
    port map (
            O => \N__13038\,
            I => \N__13032\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__13035\,
            I => \N__13029\
        );

    \I__2708\ : Sp12to4
    port map (
            O => \N__13032\,
            I => \N__13026\
        );

    \I__2707\ : Sp12to4
    port map (
            O => \N__13029\,
            I => \N__13023\
        );

    \I__2706\ : Span12Mux_s5_v
    port map (
            O => \N__13026\,
            I => \N__13018\
        );

    \I__2705\ : Span12Mux_s5_v
    port map (
            O => \N__13023\,
            I => \N__13015\
        );

    \I__2704\ : InMux
    port map (
            O => \N__13022\,
            I => \N__13012\
        );

    \I__2703\ : InMux
    port map (
            O => \N__13021\,
            I => \N__13009\
        );

    \I__2702\ : Span12Mux_v
    port map (
            O => \N__13018\,
            I => \N__13004\
        );

    \I__2701\ : Span12Mux_v
    port map (
            O => \N__13015\,
            I => \N__13004\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__13012\,
            I => \RX_ADDR_7\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__13009\,
            I => \RX_ADDR_7\
        );

    \I__2698\ : Odrv12
    port map (
            O => \N__13004\,
            I => \RX_ADDR_7\
        );

    \I__2697\ : InMux
    port map (
            O => \N__12997\,
            I => \N__12994\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__12994\,
            I => \receive_module.n129\
        );

    \I__2695\ : InMux
    port map (
            O => \N__12991\,
            I => \receive_module.n2733\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__12988\,
            I => \N__12984\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__12987\,
            I => \N__12981\
        );

    \I__2692\ : CascadeBuf
    port map (
            O => \N__12984\,
            I => \N__12978\
        );

    \I__2691\ : CascadeBuf
    port map (
            O => \N__12981\,
            I => \N__12975\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__12978\,
            I => \N__12972\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__12975\,
            I => \N__12969\
        );

    \I__2688\ : CascadeBuf
    port map (
            O => \N__12972\,
            I => \N__12966\
        );

    \I__2687\ : CascadeBuf
    port map (
            O => \N__12969\,
            I => \N__12963\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__12966\,
            I => \N__12960\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__12963\,
            I => \N__12957\
        );

    \I__2684\ : CascadeBuf
    port map (
            O => \N__12960\,
            I => \N__12954\
        );

    \I__2683\ : CascadeBuf
    port map (
            O => \N__12957\,
            I => \N__12951\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__12954\,
            I => \N__12948\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__12951\,
            I => \N__12945\
        );

    \I__2680\ : CascadeBuf
    port map (
            O => \N__12948\,
            I => \N__12942\
        );

    \I__2679\ : CascadeBuf
    port map (
            O => \N__12945\,
            I => \N__12939\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__12942\,
            I => \N__12936\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__12939\,
            I => \N__12933\
        );

    \I__2676\ : CascadeBuf
    port map (
            O => \N__12936\,
            I => \N__12930\
        );

    \I__2675\ : CascadeBuf
    port map (
            O => \N__12933\,
            I => \N__12927\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__12930\,
            I => \N__12924\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__12927\,
            I => \N__12921\
        );

    \I__2672\ : CascadeBuf
    port map (
            O => \N__12924\,
            I => \N__12918\
        );

    \I__2671\ : CascadeBuf
    port map (
            O => \N__12921\,
            I => \N__12915\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__12918\,
            I => \N__12912\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__12915\,
            I => \N__12909\
        );

    \I__2668\ : CascadeBuf
    port map (
            O => \N__12912\,
            I => \N__12906\
        );

    \I__2667\ : CascadeBuf
    port map (
            O => \N__12909\,
            I => \N__12903\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__12906\,
            I => \N__12900\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__12903\,
            I => \N__12897\
        );

    \I__2664\ : CascadeBuf
    port map (
            O => \N__12900\,
            I => \N__12894\
        );

    \I__2663\ : CascadeBuf
    port map (
            O => \N__12897\,
            I => \N__12891\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__12894\,
            I => \N__12888\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__12891\,
            I => \N__12885\
        );

    \I__2660\ : CascadeBuf
    port map (
            O => \N__12888\,
            I => \N__12882\
        );

    \I__2659\ : CascadeBuf
    port map (
            O => \N__12885\,
            I => \N__12879\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__12882\,
            I => \N__12876\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__12879\,
            I => \N__12873\
        );

    \I__2656\ : CascadeBuf
    port map (
            O => \N__12876\,
            I => \N__12870\
        );

    \I__2655\ : CascadeBuf
    port map (
            O => \N__12873\,
            I => \N__12867\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__12870\,
            I => \N__12864\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__12867\,
            I => \N__12861\
        );

    \I__2652\ : CascadeBuf
    port map (
            O => \N__12864\,
            I => \N__12858\
        );

    \I__2651\ : CascadeBuf
    port map (
            O => \N__12861\,
            I => \N__12855\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__12858\,
            I => \N__12852\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__12855\,
            I => \N__12849\
        );

    \I__2648\ : CascadeBuf
    port map (
            O => \N__12852\,
            I => \N__12846\
        );

    \I__2647\ : CascadeBuf
    port map (
            O => \N__12849\,
            I => \N__12843\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__12846\,
            I => \N__12840\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__12843\,
            I => \N__12837\
        );

    \I__2644\ : CascadeBuf
    port map (
            O => \N__12840\,
            I => \N__12834\
        );

    \I__2643\ : CascadeBuf
    port map (
            O => \N__12837\,
            I => \N__12831\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__12834\,
            I => \N__12828\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__12831\,
            I => \N__12825\
        );

    \I__2640\ : CascadeBuf
    port map (
            O => \N__12828\,
            I => \N__12822\
        );

    \I__2639\ : CascadeBuf
    port map (
            O => \N__12825\,
            I => \N__12819\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__12822\,
            I => \N__12816\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__12819\,
            I => \N__12813\
        );

    \I__2636\ : CascadeBuf
    port map (
            O => \N__12816\,
            I => \N__12810\
        );

    \I__2635\ : CascadeBuf
    port map (
            O => \N__12813\,
            I => \N__12807\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__12810\,
            I => \N__12804\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__12807\,
            I => \N__12801\
        );

    \I__2632\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12798\
        );

    \I__2631\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12795\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__12798\,
            I => \N__12792\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__12795\,
            I => \N__12789\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__12792\,
            I => \N__12786\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__12789\,
            I => \N__12783\
        );

    \I__2626\ : Sp12to4
    port map (
            O => \N__12786\,
            I => \N__12780\
        );

    \I__2625\ : Sp12to4
    port map (
            O => \N__12783\,
            I => \N__12777\
        );

    \I__2624\ : Span12Mux_s5_v
    port map (
            O => \N__12780\,
            I => \N__12772\
        );

    \I__2623\ : Span12Mux_s5_v
    port map (
            O => \N__12777\,
            I => \N__12769\
        );

    \I__2622\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12766\
        );

    \I__2621\ : InMux
    port map (
            O => \N__12775\,
            I => \N__12763\
        );

    \I__2620\ : Span12Mux_v
    port map (
            O => \N__12772\,
            I => \N__12758\
        );

    \I__2619\ : Span12Mux_v
    port map (
            O => \N__12769\,
            I => \N__12758\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__12766\,
            I => \RX_ADDR_8\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__12763\,
            I => \RX_ADDR_8\
        );

    \I__2616\ : Odrv12
    port map (
            O => \N__12758\,
            I => \RX_ADDR_8\
        );

    \I__2615\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12748\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__12748\,
            I => \receive_module.n128\
        );

    \I__2613\ : InMux
    port map (
            O => \N__12745\,
            I => \bfn_18_15_0_\
        );

    \I__2612\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12739\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__12739\,
            I => \N__12736\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__12736\,
            I => \N__12733\
        );

    \I__2609\ : Sp12to4
    port map (
            O => \N__12733\,
            I => \N__12730\
        );

    \I__2608\ : Odrv12
    port map (
            O => \N__12730\,
            I => \line_buffer.n726\
        );

    \I__2607\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12724\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__12724\,
            I => \N__12721\
        );

    \I__2605\ : Span12Mux_v
    port map (
            O => \N__12721\,
            I => \N__12718\
        );

    \I__2604\ : Span12Mux_v
    port map (
            O => \N__12718\,
            I => \N__12715\
        );

    \I__2603\ : Odrv12
    port map (
            O => \N__12715\,
            I => \line_buffer.n718\
        );

    \I__2602\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12709\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__12709\,
            I => \N__12706\
        );

    \I__2600\ : Span12Mux_v
    port map (
            O => \N__12706\,
            I => \N__12703\
        );

    \I__2599\ : Odrv12
    port map (
            O => \N__12703\,
            I => \line_buffer.n629\
        );

    \I__2598\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12697\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__12697\,
            I => \N__12694\
        );

    \I__2596\ : Span4Mux_v
    port map (
            O => \N__12694\,
            I => \N__12691\
        );

    \I__2595\ : Span4Mux_h
    port map (
            O => \N__12691\,
            I => \N__12688\
        );

    \I__2594\ : Span4Mux_h
    port map (
            O => \N__12688\,
            I => \N__12685\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__12685\,
            I => \line_buffer.n621\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__12682\,
            I => \line_buffer.n3161_cascade_\
        );

    \I__2591\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12676\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__12676\,
            I => \line_buffer.n3164\
        );

    \I__2589\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12670\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__12670\,
            I => \N__12667\
        );

    \I__2587\ : Span4Mux_h
    port map (
            O => \N__12667\,
            I => \N__12664\
        );

    \I__2586\ : Span4Mux_h
    port map (
            O => \N__12664\,
            I => \N__12661\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__12661\,
            I => \line_buffer.n630\
        );

    \I__2584\ : InMux
    port map (
            O => \N__12658\,
            I => \N__12655\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__12655\,
            I => \N__12652\
        );

    \I__2582\ : Span4Mux_h
    port map (
            O => \N__12652\,
            I => \N__12649\
        );

    \I__2581\ : Span4Mux_h
    port map (
            O => \N__12649\,
            I => \N__12646\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__12646\,
            I => \N__12643\
        );

    \I__2579\ : Odrv4
    port map (
            O => \N__12643\,
            I => \line_buffer.n622\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12637\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__12637\,
            I => \N__12634\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__12634\,
            I => \line_buffer.n3042\
        );

    \I__2575\ : SRMux
    port map (
            O => \N__12631\,
            I => \N__12628\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__12628\,
            I => \N__12623\
        );

    \I__2573\ : SRMux
    port map (
            O => \N__12627\,
            I => \N__12620\
        );

    \I__2572\ : SRMux
    port map (
            O => \N__12626\,
            I => \N__12617\
        );

    \I__2571\ : Span4Mux_s2_v
    port map (
            O => \N__12623\,
            I => \N__12607\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__12620\,
            I => \N__12607\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__12617\,
            I => \N__12607\
        );

    \I__2568\ : SRMux
    port map (
            O => \N__12616\,
            I => \N__12604\
        );

    \I__2567\ : SRMux
    port map (
            O => \N__12615\,
            I => \N__12601\
        );

    \I__2566\ : SRMux
    port map (
            O => \N__12614\,
            I => \N__12596\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__12607\,
            I => \N__12587\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__12604\,
            I => \N__12587\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__12601\,
            I => \N__12587\
        );

    \I__2562\ : SRMux
    port map (
            O => \N__12600\,
            I => \N__12584\
        );

    \I__2561\ : SRMux
    port map (
            O => \N__12599\,
            I => \N__12581\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__12596\,
            I => \N__12576\
        );

    \I__2559\ : SRMux
    port map (
            O => \N__12595\,
            I => \N__12573\
        );

    \I__2558\ : SRMux
    port map (
            O => \N__12594\,
            I => \N__12570\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__12587\,
            I => \N__12561\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__12584\,
            I => \N__12561\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__12581\,
            I => \N__12561\
        );

    \I__2554\ : SRMux
    port map (
            O => \N__12580\,
            I => \N__12558\
        );

    \I__2553\ : SRMux
    port map (
            O => \N__12579\,
            I => \N__12555\
        );

    \I__2552\ : Span4Mux_s2_v
    port map (
            O => \N__12576\,
            I => \N__12546\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__12573\,
            I => \N__12546\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__12570\,
            I => \N__12546\
        );

    \I__2549\ : SRMux
    port map (
            O => \N__12569\,
            I => \N__12543\
        );

    \I__2548\ : SRMux
    port map (
            O => \N__12568\,
            I => \N__12540\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__12561\,
            I => \N__12529\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__12558\,
            I => \N__12529\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__12555\,
            I => \N__12529\
        );

    \I__2544\ : SRMux
    port map (
            O => \N__12554\,
            I => \N__12526\
        );

    \I__2543\ : SRMux
    port map (
            O => \N__12553\,
            I => \N__12523\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__12546\,
            I => \N__12514\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__12543\,
            I => \N__12514\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__12540\,
            I => \N__12514\
        );

    \I__2539\ : SRMux
    port map (
            O => \N__12539\,
            I => \N__12511\
        );

    \I__2538\ : SRMux
    port map (
            O => \N__12538\,
            I => \N__12508\
        );

    \I__2537\ : IoInMux
    port map (
            O => \N__12537\,
            I => \N__12503\
        );

    \I__2536\ : IoInMux
    port map (
            O => \N__12536\,
            I => \N__12500\
        );

    \I__2535\ : Span4Mux_v
    port map (
            O => \N__12529\,
            I => \N__12493\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__12526\,
            I => \N__12493\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__12523\,
            I => \N__12493\
        );

    \I__2532\ : SRMux
    port map (
            O => \N__12522\,
            I => \N__12490\
        );

    \I__2531\ : SRMux
    port map (
            O => \N__12521\,
            I => \N__12487\
        );

    \I__2530\ : Span4Mux_v
    port map (
            O => \N__12514\,
            I => \N__12478\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__12511\,
            I => \N__12478\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__12508\,
            I => \N__12478\
        );

    \I__2527\ : SRMux
    port map (
            O => \N__12507\,
            I => \N__12475\
        );

    \I__2526\ : SRMux
    port map (
            O => \N__12506\,
            I => \N__12472\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__12503\,
            I => \N__12465\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__12500\,
            I => \N__12465\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__12493\,
            I => \N__12458\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__12490\,
            I => \N__12458\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__12487\,
            I => \N__12458\
        );

    \I__2520\ : SRMux
    port map (
            O => \N__12486\,
            I => \N__12455\
        );

    \I__2519\ : SRMux
    port map (
            O => \N__12485\,
            I => \N__12452\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__12478\,
            I => \N__12444\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__12475\,
            I => \N__12444\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__12472\,
            I => \N__12444\
        );

    \I__2515\ : SRMux
    port map (
            O => \N__12471\,
            I => \N__12441\
        );

    \I__2514\ : SRMux
    port map (
            O => \N__12470\,
            I => \N__12438\
        );

    \I__2513\ : IoSpan4Mux
    port map (
            O => \N__12465\,
            I => \N__12433\
        );

    \I__2512\ : Span4Mux_v
    port map (
            O => \N__12458\,
            I => \N__12426\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__12455\,
            I => \N__12426\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__12452\,
            I => \N__12426\
        );

    \I__2509\ : SRMux
    port map (
            O => \N__12451\,
            I => \N__12423\
        );

    \I__2508\ : Span4Mux_v
    port map (
            O => \N__12444\,
            I => \N__12416\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__12441\,
            I => \N__12416\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__12438\,
            I => \N__12416\
        );

    \I__2505\ : SRMux
    port map (
            O => \N__12437\,
            I => \N__12413\
        );

    \I__2504\ : SRMux
    port map (
            O => \N__12436\,
            I => \N__12410\
        );

    \I__2503\ : Span4Mux_s0_v
    port map (
            O => \N__12433\,
            I => \N__12404\
        );

    \I__2502\ : Span4Mux_v
    port map (
            O => \N__12426\,
            I => \N__12399\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__12423\,
            I => \N__12399\
        );

    \I__2500\ : Span4Mux_v
    port map (
            O => \N__12416\,
            I => \N__12392\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__12413\,
            I => \N__12392\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__12410\,
            I => \N__12392\
        );

    \I__2497\ : SRMux
    port map (
            O => \N__12409\,
            I => \N__12389\
        );

    \I__2496\ : SRMux
    port map (
            O => \N__12408\,
            I => \N__12386\
        );

    \I__2495\ : SRMux
    port map (
            O => \N__12407\,
            I => \N__12383\
        );

    \I__2494\ : Sp12to4
    port map (
            O => \N__12404\,
            I => \N__12380\
        );

    \I__2493\ : Span4Mux_s1_v
    port map (
            O => \N__12399\,
            I => \N__12377\
        );

    \I__2492\ : Span4Mux_v
    port map (
            O => \N__12392\,
            I => \N__12370\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__12389\,
            I => \N__12370\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__12386\,
            I => \N__12370\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12383\,
            I => \N__12367\
        );

    \I__2488\ : Span12Mux_s11_v
    port map (
            O => \N__12380\,
            I => \N__12364\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__12377\,
            I => \N__12361\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__12370\,
            I => \N__12356\
        );

    \I__2485\ : Span4Mux_s1_v
    port map (
            O => \N__12367\,
            I => \N__12356\
        );

    \I__2484\ : Span12Mux_v
    port map (
            O => \N__12364\,
            I => \N__12353\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__12361\,
            I => \N__12348\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__12356\,
            I => \N__12348\
        );

    \I__2481\ : Odrv12
    port map (
            O => \N__12353\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__12348\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2479\ : InMux
    port map (
            O => \N__12343\,
            I => \N__12340\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__12340\,
            I => \N__12337\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__12337\,
            I => \N__12334\
        );

    \I__2476\ : Sp12to4
    port map (
            O => \N__12334\,
            I => \N__12331\
        );

    \I__2475\ : Span12Mux_h
    port map (
            O => \N__12331\,
            I => \N__12328\
        );

    \I__2474\ : Odrv12
    port map (
            O => \N__12328\,
            I => \line_buffer.n623\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__12325\,
            I => \N__12322\
        );

    \I__2472\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12319\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__12319\,
            I => \N__12316\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__12316\,
            I => \N__12313\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__12313\,
            I => \N__12310\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__12310\,
            I => \N__12307\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__12307\,
            I => \line_buffer.n615\
        );

    \I__2466\ : InMux
    port map (
            O => \N__12304\,
            I => \N__12301\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__12301\,
            I => \N__12298\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__12298\,
            I => \N__12295\
        );

    \I__2463\ : Sp12to4
    port map (
            O => \N__12295\,
            I => \N__12292\
        );

    \I__2462\ : Odrv12
    port map (
            O => \N__12292\,
            I => \line_buffer.n720\
        );

    \I__2461\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12286\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__12286\,
            I => \N__12283\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__12283\,
            I => \N__12280\
        );

    \I__2458\ : Span4Mux_v
    port map (
            O => \N__12280\,
            I => \N__12277\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__12277\,
            I => \N__12274\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__12274\,
            I => \line_buffer.n712\
        );

    \I__2455\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12268\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__12268\,
            I => \line_buffer.n3113\
        );

    \I__2453\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12262\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__12262\,
            I => \N__12259\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__12259\,
            I => \N__12256\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__12256\,
            I => \N__12253\
        );

    \I__2449\ : Sp12to4
    port map (
            O => \N__12253\,
            I => \N__12250\
        );

    \I__2448\ : Odrv12
    port map (
            O => \N__12250\,
            I => \line_buffer.n688\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__12247\,
            I => \N__12244\
        );

    \I__2446\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12241\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__12241\,
            I => \N__12238\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__12238\,
            I => \N__12235\
        );

    \I__2443\ : Span4Mux_h
    port map (
            O => \N__12235\,
            I => \N__12232\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__12232\,
            I => \line_buffer.n680\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__12229\,
            I => \line_buffer.n3122_cascade_\
        );

    \I__2440\ : InMux
    port map (
            O => \N__12226\,
            I => \N__12223\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__12223\,
            I => \line_buffer.n3116\
        );

    \I__2438\ : InMux
    port map (
            O => \N__12220\,
            I => \N__12217\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__12217\,
            I => \N__12214\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__12214\,
            I => \N__12211\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__12211\,
            I => \TX_DATA_0\
        );

    \I__2434\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12205\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__12205\,
            I => \N__12202\
        );

    \I__2432\ : Span12Mux_v
    port map (
            O => \N__12202\,
            I => \N__12199\
        );

    \I__2431\ : Span12Mux_v
    port map (
            O => \N__12199\,
            I => \N__12196\
        );

    \I__2430\ : Odrv12
    port map (
            O => \N__12196\,
            I => \line_buffer.n745\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__12193\,
            I => \N__12190\
        );

    \I__2428\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12187\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12184\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__12184\,
            I => \N__12181\
        );

    \I__2425\ : Span4Mux_h
    port map (
            O => \N__12181\,
            I => \N__12178\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__12178\,
            I => \N__12175\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__12175\,
            I => \line_buffer.n753\
        );

    \I__2422\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12169\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__12169\,
            I => \line_buffer.n3137\
        );

    \I__2420\ : SRMux
    port map (
            O => \N__12166\,
            I => \N__12162\
        );

    \I__2419\ : SRMux
    port map (
            O => \N__12165\,
            I => \N__12157\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__12162\,
            I => \N__12154\
        );

    \I__2417\ : SRMux
    port map (
            O => \N__12161\,
            I => \N__12151\
        );

    \I__2416\ : SRMux
    port map (
            O => \N__12160\,
            I => \N__12148\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__12157\,
            I => \N__12145\
        );

    \I__2414\ : Span4Mux_s1_v
    port map (
            O => \N__12154\,
            I => \N__12138\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__12151\,
            I => \N__12138\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__12148\,
            I => \N__12138\
        );

    \I__2411\ : Span4Mux_h
    port map (
            O => \N__12145\,
            I => \N__12135\
        );

    \I__2410\ : Sp12to4
    port map (
            O => \N__12138\,
            I => \N__12132\
        );

    \I__2409\ : Span4Mux_h
    port map (
            O => \N__12135\,
            I => \N__12129\
        );

    \I__2408\ : Span12Mux_v
    port map (
            O => \N__12132\,
            I => \N__12126\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__12129\,
            I => \N__12123\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__12126\,
            I => \line_buffer.n761\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__12123\,
            I => \line_buffer.n761\
        );

    \I__2404\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12115\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__12115\,
            I => \N__12111\
        );

    \I__2402\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12108\
        );

    \I__2401\ : Span4Mux_h
    port map (
            O => \N__12111\,
            I => \N__12105\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__12108\,
            I => \transmit_module.n387\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__12105\,
            I => \transmit_module.n387\
        );

    \I__2398\ : IoInMux
    port map (
            O => \N__12100\,
            I => \N__12097\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__12097\,
            I => \N__12094\
        );

    \I__2396\ : Span12Mux_s10_h
    port map (
            O => \N__12094\,
            I => \N__12090\
        );

    \I__2395\ : InMux
    port map (
            O => \N__12093\,
            I => \N__12087\
        );

    \I__2394\ : Span12Mux_v
    port map (
            O => \N__12090\,
            I => \N__12082\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__12087\,
            I => \N__12079\
        );

    \I__2392\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12076\
        );

    \I__2391\ : InMux
    port map (
            O => \N__12085\,
            I => \N__12073\
        );

    \I__2390\ : Odrv12
    port map (
            O => \N__12082\,
            I => \DEBUG_c_1\
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__12079\,
            I => \DEBUG_c_1\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__12076\,
            I => \DEBUG_c_1\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__12073\,
            I => \DEBUG_c_1\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__12064\,
            I => \N__12060\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__12063\,
            I => \N__12057\
        );

    \I__2384\ : CascadeBuf
    port map (
            O => \N__12060\,
            I => \N__12054\
        );

    \I__2383\ : CascadeBuf
    port map (
            O => \N__12057\,
            I => \N__12051\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__12054\,
            I => \N__12048\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__12051\,
            I => \N__12045\
        );

    \I__2380\ : CascadeBuf
    port map (
            O => \N__12048\,
            I => \N__12042\
        );

    \I__2379\ : CascadeBuf
    port map (
            O => \N__12045\,
            I => \N__12039\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__12042\,
            I => \N__12036\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__12039\,
            I => \N__12033\
        );

    \I__2376\ : CascadeBuf
    port map (
            O => \N__12036\,
            I => \N__12030\
        );

    \I__2375\ : CascadeBuf
    port map (
            O => \N__12033\,
            I => \N__12027\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__12030\,
            I => \N__12024\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__12027\,
            I => \N__12021\
        );

    \I__2372\ : CascadeBuf
    port map (
            O => \N__12024\,
            I => \N__12018\
        );

    \I__2371\ : CascadeBuf
    port map (
            O => \N__12021\,
            I => \N__12015\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__12018\,
            I => \N__12012\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__12015\,
            I => \N__12009\
        );

    \I__2368\ : CascadeBuf
    port map (
            O => \N__12012\,
            I => \N__12006\
        );

    \I__2367\ : CascadeBuf
    port map (
            O => \N__12009\,
            I => \N__12003\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__12006\,
            I => \N__12000\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__12003\,
            I => \N__11997\
        );

    \I__2364\ : CascadeBuf
    port map (
            O => \N__12000\,
            I => \N__11994\
        );

    \I__2363\ : CascadeBuf
    port map (
            O => \N__11997\,
            I => \N__11991\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__11994\,
            I => \N__11988\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__11991\,
            I => \N__11985\
        );

    \I__2360\ : CascadeBuf
    port map (
            O => \N__11988\,
            I => \N__11982\
        );

    \I__2359\ : CascadeBuf
    port map (
            O => \N__11985\,
            I => \N__11979\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__11982\,
            I => \N__11976\
        );

    \I__2357\ : CascadeMux
    port map (
            O => \N__11979\,
            I => \N__11973\
        );

    \I__2356\ : CascadeBuf
    port map (
            O => \N__11976\,
            I => \N__11970\
        );

    \I__2355\ : CascadeBuf
    port map (
            O => \N__11973\,
            I => \N__11967\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__11970\,
            I => \N__11964\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__11967\,
            I => \N__11961\
        );

    \I__2352\ : CascadeBuf
    port map (
            O => \N__11964\,
            I => \N__11958\
        );

    \I__2351\ : CascadeBuf
    port map (
            O => \N__11961\,
            I => \N__11955\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__11958\,
            I => \N__11952\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__11955\,
            I => \N__11949\
        );

    \I__2348\ : CascadeBuf
    port map (
            O => \N__11952\,
            I => \N__11946\
        );

    \I__2347\ : CascadeBuf
    port map (
            O => \N__11949\,
            I => \N__11943\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__11946\,
            I => \N__11940\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__11943\,
            I => \N__11937\
        );

    \I__2344\ : CascadeBuf
    port map (
            O => \N__11940\,
            I => \N__11934\
        );

    \I__2343\ : CascadeBuf
    port map (
            O => \N__11937\,
            I => \N__11931\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__11934\,
            I => \N__11928\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__11931\,
            I => \N__11925\
        );

    \I__2340\ : CascadeBuf
    port map (
            O => \N__11928\,
            I => \N__11922\
        );

    \I__2339\ : CascadeBuf
    port map (
            O => \N__11925\,
            I => \N__11919\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__11922\,
            I => \N__11916\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__11919\,
            I => \N__11913\
        );

    \I__2336\ : CascadeBuf
    port map (
            O => \N__11916\,
            I => \N__11910\
        );

    \I__2335\ : CascadeBuf
    port map (
            O => \N__11913\,
            I => \N__11907\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__11910\,
            I => \N__11904\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__11907\,
            I => \N__11901\
        );

    \I__2332\ : CascadeBuf
    port map (
            O => \N__11904\,
            I => \N__11898\
        );

    \I__2331\ : CascadeBuf
    port map (
            O => \N__11901\,
            I => \N__11895\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__11898\,
            I => \N__11892\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__11895\,
            I => \N__11889\
        );

    \I__2328\ : CascadeBuf
    port map (
            O => \N__11892\,
            I => \N__11886\
        );

    \I__2327\ : CascadeBuf
    port map (
            O => \N__11889\,
            I => \N__11883\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__11886\,
            I => \N__11880\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__11883\,
            I => \N__11877\
        );

    \I__2324\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11874\
        );

    \I__2323\ : InMux
    port map (
            O => \N__11877\,
            I => \N__11871\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__11874\,
            I => \N__11868\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__11871\,
            I => \N__11865\
        );

    \I__2320\ : Span12Mux_s11_h
    port map (
            O => \N__11868\,
            I => \N__11862\
        );

    \I__2319\ : Span12Mux_s8_h
    port map (
            O => \N__11865\,
            I => \N__11859\
        );

    \I__2318\ : Span12Mux_v
    port map (
            O => \N__11862\,
            I => \N__11854\
        );

    \I__2317\ : Span12Mux_v
    port map (
            O => \N__11859\,
            I => \N__11854\
        );

    \I__2316\ : Odrv12
    port map (
            O => \N__11854\,
            I => n27
        );

    \I__2315\ : IoInMux
    port map (
            O => \N__11851\,
            I => \N__11848\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__11848\,
            I => \N__11845\
        );

    \I__2313\ : Span4Mux_s3_h
    port map (
            O => \N__11845\,
            I => \N__11842\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__11842\,
            I => \N__11839\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__11839\,
            I => \N__11836\
        );

    \I__2310\ : Span4Mux_h
    port map (
            O => \N__11836\,
            I => \N__11830\
        );

    \I__2309\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11827\
        );

    \I__2308\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11824\
        );

    \I__2307\ : InMux
    port map (
            O => \N__11833\,
            I => \N__11821\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__11830\,
            I => \DEBUG_c_7\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__11827\,
            I => \DEBUG_c_7\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__11824\,
            I => \DEBUG_c_7\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__11821\,
            I => \DEBUG_c_7\
        );

    \I__2302\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11808\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__11811\,
            I => \N__11805\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__11808\,
            I => \N__11802\
        );

    \I__2299\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11799\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__11802\,
            I => \N__11796\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__11799\,
            I => \transmit_module.n381\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__11796\,
            I => \transmit_module.n381\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__11791\,
            I => \N__11788\
        );

    \I__2294\ : CascadeBuf
    port map (
            O => \N__11788\,
            I => \N__11785\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__11785\,
            I => \N__11781\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__11784\,
            I => \N__11778\
        );

    \I__2291\ : CascadeBuf
    port map (
            O => \N__11781\,
            I => \N__11775\
        );

    \I__2290\ : CascadeBuf
    port map (
            O => \N__11778\,
            I => \N__11772\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__11775\,
            I => \N__11769\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__11772\,
            I => \N__11766\
        );

    \I__2287\ : CascadeBuf
    port map (
            O => \N__11769\,
            I => \N__11763\
        );

    \I__2286\ : CascadeBuf
    port map (
            O => \N__11766\,
            I => \N__11760\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__11763\,
            I => \N__11757\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__11760\,
            I => \N__11754\
        );

    \I__2283\ : CascadeBuf
    port map (
            O => \N__11757\,
            I => \N__11751\
        );

    \I__2282\ : CascadeBuf
    port map (
            O => \N__11754\,
            I => \N__11748\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__11751\,
            I => \N__11745\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__11748\,
            I => \N__11742\
        );

    \I__2279\ : CascadeBuf
    port map (
            O => \N__11745\,
            I => \N__11739\
        );

    \I__2278\ : CascadeBuf
    port map (
            O => \N__11742\,
            I => \N__11736\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__11739\,
            I => \N__11733\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__11736\,
            I => \N__11730\
        );

    \I__2275\ : CascadeBuf
    port map (
            O => \N__11733\,
            I => \N__11727\
        );

    \I__2274\ : CascadeBuf
    port map (
            O => \N__11730\,
            I => \N__11724\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__11727\,
            I => \N__11721\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__11724\,
            I => \N__11718\
        );

    \I__2271\ : CascadeBuf
    port map (
            O => \N__11721\,
            I => \N__11715\
        );

    \I__2270\ : CascadeBuf
    port map (
            O => \N__11718\,
            I => \N__11712\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__11715\,
            I => \N__11709\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__11712\,
            I => \N__11706\
        );

    \I__2267\ : CascadeBuf
    port map (
            O => \N__11709\,
            I => \N__11703\
        );

    \I__2266\ : CascadeBuf
    port map (
            O => \N__11706\,
            I => \N__11700\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__11703\,
            I => \N__11697\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__11700\,
            I => \N__11694\
        );

    \I__2263\ : CascadeBuf
    port map (
            O => \N__11697\,
            I => \N__11691\
        );

    \I__2262\ : CascadeBuf
    port map (
            O => \N__11694\,
            I => \N__11688\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__11691\,
            I => \N__11685\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__11688\,
            I => \N__11682\
        );

    \I__2259\ : CascadeBuf
    port map (
            O => \N__11685\,
            I => \N__11679\
        );

    \I__2258\ : CascadeBuf
    port map (
            O => \N__11682\,
            I => \N__11676\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__11679\,
            I => \N__11673\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__11676\,
            I => \N__11670\
        );

    \I__2255\ : CascadeBuf
    port map (
            O => \N__11673\,
            I => \N__11667\
        );

    \I__2254\ : CascadeBuf
    port map (
            O => \N__11670\,
            I => \N__11664\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__11667\,
            I => \N__11661\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__11664\,
            I => \N__11658\
        );

    \I__2251\ : CascadeBuf
    port map (
            O => \N__11661\,
            I => \N__11655\
        );

    \I__2250\ : CascadeBuf
    port map (
            O => \N__11658\,
            I => \N__11652\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__11655\,
            I => \N__11649\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__11652\,
            I => \N__11646\
        );

    \I__2247\ : CascadeBuf
    port map (
            O => \N__11649\,
            I => \N__11643\
        );

    \I__2246\ : CascadeBuf
    port map (
            O => \N__11646\,
            I => \N__11640\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__11643\,
            I => \N__11637\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__11640\,
            I => \N__11634\
        );

    \I__2243\ : CascadeBuf
    port map (
            O => \N__11637\,
            I => \N__11631\
        );

    \I__2242\ : CascadeBuf
    port map (
            O => \N__11634\,
            I => \N__11628\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__11631\,
            I => \N__11625\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__11628\,
            I => \N__11622\
        );

    \I__2239\ : CascadeBuf
    port map (
            O => \N__11625\,
            I => \N__11619\
        );

    \I__2238\ : CascadeBuf
    port map (
            O => \N__11622\,
            I => \N__11616\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__11619\,
            I => \N__11613\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__11616\,
            I => \N__11610\
        );

    \I__2235\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11607\
        );

    \I__2234\ : CascadeBuf
    port map (
            O => \N__11610\,
            I => \N__11604\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__11607\,
            I => \N__11601\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__11604\,
            I => \N__11598\
        );

    \I__2231\ : Span4Mux_h
    port map (
            O => \N__11601\,
            I => \N__11595\
        );

    \I__2230\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11592\
        );

    \I__2229\ : Sp12to4
    port map (
            O => \N__11595\,
            I => \N__11589\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__11592\,
            I => \N__11586\
        );

    \I__2227\ : Span12Mux_h
    port map (
            O => \N__11589\,
            I => \N__11581\
        );

    \I__2226\ : Span12Mux_s10_h
    port map (
            O => \N__11586\,
            I => \N__11581\
        );

    \I__2225\ : Span12Mux_v
    port map (
            O => \N__11581\,
            I => \N__11578\
        );

    \I__2224\ : Odrv12
    port map (
            O => \N__11578\,
            I => n21
        );

    \I__2223\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11572\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__11572\,
            I => \N__11568\
        );

    \I__2221\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11565\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__11568\,
            I => \N__11562\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__11565\,
            I => \transmit_module.n385\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__11562\,
            I => \transmit_module.n385\
        );

    \I__2217\ : IoInMux
    port map (
            O => \N__11557\,
            I => \N__11554\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__11554\,
            I => \N__11551\
        );

    \I__2215\ : Span4Mux_s3_h
    port map (
            O => \N__11551\,
            I => \N__11548\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__11548\,
            I => \N__11545\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__11545\,
            I => \N__11542\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__11542\,
            I => \N__11537\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__11541\,
            I => \N__11534\
        );

    \I__2210\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11531\
        );

    \I__2209\ : Span4Mux_h
    port map (
            O => \N__11537\,
            I => \N__11527\
        );

    \I__2208\ : InMux
    port map (
            O => \N__11534\,
            I => \N__11524\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__11531\,
            I => \N__11521\
        );

    \I__2206\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11518\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__11527\,
            I => \DEBUG_c_3\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__11524\,
            I => \DEBUG_c_3\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__11521\,
            I => \DEBUG_c_3\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__11518\,
            I => \DEBUG_c_3\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__11509\,
            I => \N__11505\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__11508\,
            I => \N__11502\
        );

    \I__2199\ : CascadeBuf
    port map (
            O => \N__11505\,
            I => \N__11499\
        );

    \I__2198\ : CascadeBuf
    port map (
            O => \N__11502\,
            I => \N__11496\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__11499\,
            I => \N__11493\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__11496\,
            I => \N__11490\
        );

    \I__2195\ : CascadeBuf
    port map (
            O => \N__11493\,
            I => \N__11487\
        );

    \I__2194\ : CascadeBuf
    port map (
            O => \N__11490\,
            I => \N__11484\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__11487\,
            I => \N__11481\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__11484\,
            I => \N__11478\
        );

    \I__2191\ : CascadeBuf
    port map (
            O => \N__11481\,
            I => \N__11475\
        );

    \I__2190\ : CascadeBuf
    port map (
            O => \N__11478\,
            I => \N__11472\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__11475\,
            I => \N__11469\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__11472\,
            I => \N__11466\
        );

    \I__2187\ : CascadeBuf
    port map (
            O => \N__11469\,
            I => \N__11463\
        );

    \I__2186\ : CascadeBuf
    port map (
            O => \N__11466\,
            I => \N__11460\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__11463\,
            I => \N__11457\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__11460\,
            I => \N__11454\
        );

    \I__2183\ : CascadeBuf
    port map (
            O => \N__11457\,
            I => \N__11451\
        );

    \I__2182\ : CascadeBuf
    port map (
            O => \N__11454\,
            I => \N__11448\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__11451\,
            I => \N__11445\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__11448\,
            I => \N__11442\
        );

    \I__2179\ : CascadeBuf
    port map (
            O => \N__11445\,
            I => \N__11439\
        );

    \I__2178\ : CascadeBuf
    port map (
            O => \N__11442\,
            I => \N__11436\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__11439\,
            I => \N__11433\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__11436\,
            I => \N__11430\
        );

    \I__2175\ : CascadeBuf
    port map (
            O => \N__11433\,
            I => \N__11427\
        );

    \I__2174\ : CascadeBuf
    port map (
            O => \N__11430\,
            I => \N__11424\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__11427\,
            I => \N__11421\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__11424\,
            I => \N__11418\
        );

    \I__2171\ : CascadeBuf
    port map (
            O => \N__11421\,
            I => \N__11415\
        );

    \I__2170\ : CascadeBuf
    port map (
            O => \N__11418\,
            I => \N__11412\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__11415\,
            I => \N__11409\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__11412\,
            I => \N__11406\
        );

    \I__2167\ : CascadeBuf
    port map (
            O => \N__11409\,
            I => \N__11403\
        );

    \I__2166\ : CascadeBuf
    port map (
            O => \N__11406\,
            I => \N__11400\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__11403\,
            I => \N__11397\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__11400\,
            I => \N__11394\
        );

    \I__2163\ : CascadeBuf
    port map (
            O => \N__11397\,
            I => \N__11391\
        );

    \I__2162\ : CascadeBuf
    port map (
            O => \N__11394\,
            I => \N__11388\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__11391\,
            I => \N__11385\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__11388\,
            I => \N__11382\
        );

    \I__2159\ : CascadeBuf
    port map (
            O => \N__11385\,
            I => \N__11379\
        );

    \I__2158\ : CascadeBuf
    port map (
            O => \N__11382\,
            I => \N__11376\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__11379\,
            I => \N__11373\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__11376\,
            I => \N__11370\
        );

    \I__2155\ : CascadeBuf
    port map (
            O => \N__11373\,
            I => \N__11367\
        );

    \I__2154\ : CascadeBuf
    port map (
            O => \N__11370\,
            I => \N__11364\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__11367\,
            I => \N__11361\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__11364\,
            I => \N__11358\
        );

    \I__2151\ : CascadeBuf
    port map (
            O => \N__11361\,
            I => \N__11355\
        );

    \I__2150\ : CascadeBuf
    port map (
            O => \N__11358\,
            I => \N__11352\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__11355\,
            I => \N__11349\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__11352\,
            I => \N__11346\
        );

    \I__2147\ : CascadeBuf
    port map (
            O => \N__11349\,
            I => \N__11343\
        );

    \I__2146\ : CascadeBuf
    port map (
            O => \N__11346\,
            I => \N__11340\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__11343\,
            I => \N__11337\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__11340\,
            I => \N__11334\
        );

    \I__2143\ : CascadeBuf
    port map (
            O => \N__11337\,
            I => \N__11331\
        );

    \I__2142\ : CascadeBuf
    port map (
            O => \N__11334\,
            I => \N__11328\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__11331\,
            I => \N__11325\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__11328\,
            I => \N__11322\
        );

    \I__2139\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11319\
        );

    \I__2138\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11316\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__11319\,
            I => \N__11313\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__11316\,
            I => \N__11310\
        );

    \I__2135\ : Span12Mux_h
    port map (
            O => \N__11313\,
            I => \N__11307\
        );

    \I__2134\ : Sp12to4
    port map (
            O => \N__11310\,
            I => \N__11304\
        );

    \I__2133\ : Span12Mux_v
    port map (
            O => \N__11307\,
            I => \N__11299\
        );

    \I__2132\ : Span12Mux_v
    port map (
            O => \N__11304\,
            I => \N__11299\
        );

    \I__2131\ : Odrv12
    port map (
            O => \N__11299\,
            I => n25_adj_573
        );

    \I__2130\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__11293\,
            I => \N__11290\
        );

    \I__2128\ : Odrv12
    port map (
            O => \N__11290\,
            I => \line_buffer.n3028\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__11287\,
            I => \line_buffer.n3125_cascade_\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11281\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__11278\,
            I => \TX_DATA_7\
        );

    \I__2123\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11272\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__2121\ : Span4Mux_v
    port map (
            O => \N__11269\,
            I => \N__11266\
        );

    \I__2120\ : Sp12to4
    port map (
            O => \N__11266\,
            I => \N__11263\
        );

    \I__2119\ : Odrv12
    port map (
            O => \N__11263\,
            I => \line_buffer.n727\
        );

    \I__2118\ : InMux
    port map (
            O => \N__11260\,
            I => \N__11257\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__11257\,
            I => \N__11254\
        );

    \I__2116\ : Span12Mux_v
    port map (
            O => \N__11254\,
            I => \N__11251\
        );

    \I__2115\ : Span12Mux_v
    port map (
            O => \N__11251\,
            I => \N__11248\
        );

    \I__2114\ : Odrv12
    port map (
            O => \N__11248\,
            I => \line_buffer.n719\
        );

    \I__2113\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11242\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__11242\,
            I => \line_buffer.n3043\
        );

    \I__2111\ : InMux
    port map (
            O => \N__11239\,
            I => \N__11236\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__11236\,
            I => \N__11233\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__11233\,
            I => \N__11230\
        );

    \I__2108\ : Span4Mux_h
    port map (
            O => \N__11230\,
            I => \N__11227\
        );

    \I__2107\ : Span4Mux_h
    port map (
            O => \N__11227\,
            I => \N__11224\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__11224\,
            I => \N__11221\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__11221\,
            I => \line_buffer.n689\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__11218\,
            I => \N__11215\
        );

    \I__2103\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11212\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__11212\,
            I => \N__11209\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__11209\,
            I => \N__11206\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__11206\,
            I => \N__11203\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__11203\,
            I => \N__11200\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__11200\,
            I => \line_buffer.n681\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__11197\,
            I => \line_buffer.n3140_cascade_\
        );

    \I__2096\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11191\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__11191\,
            I => \TX_DATA_1\
        );

    \I__2094\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11185\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__11185\,
            I => \N__11182\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__11182\,
            I => \line_buffer.n713\
        );

    \I__2091\ : InMux
    port map (
            O => \N__11179\,
            I => \N__11176\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__11176\,
            I => \N__11173\
        );

    \I__2089\ : Span4Mux_v
    port map (
            O => \N__11173\,
            I => \N__11170\
        );

    \I__2088\ : Span4Mux_h
    port map (
            O => \N__11170\,
            I => \N__11167\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__11167\,
            I => \N__11164\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__11164\,
            I => \line_buffer.n721\
        );

    \I__2085\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11158\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__11158\,
            I => \N__11155\
        );

    \I__2083\ : Span12Mux_v
    port map (
            O => \N__11155\,
            I => \N__11152\
        );

    \I__2082\ : Odrv12
    port map (
            O => \N__11152\,
            I => \line_buffer.n624\
        );

    \I__2081\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11146\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__11146\,
            I => \N__11143\
        );

    \I__2079\ : Span12Mux_v
    port map (
            O => \N__11143\,
            I => \N__11140\
        );

    \I__2078\ : Odrv12
    port map (
            O => \N__11140\,
            I => \line_buffer.n616\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__11137\,
            I => \line_buffer.n3107_cascade_\
        );

    \I__2076\ : InMux
    port map (
            O => \N__11134\,
            I => \N__11131\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__11131\,
            I => \line_buffer.n3110\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__11128\,
            I => \N__11124\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__11127\,
            I => \N__11121\
        );

    \I__2072\ : CascadeBuf
    port map (
            O => \N__11124\,
            I => \N__11118\
        );

    \I__2071\ : CascadeBuf
    port map (
            O => \N__11121\,
            I => \N__11115\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__11118\,
            I => \N__11112\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__11115\,
            I => \N__11109\
        );

    \I__2068\ : CascadeBuf
    port map (
            O => \N__11112\,
            I => \N__11106\
        );

    \I__2067\ : CascadeBuf
    port map (
            O => \N__11109\,
            I => \N__11103\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__11106\,
            I => \N__11100\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__11103\,
            I => \N__11097\
        );

    \I__2064\ : CascadeBuf
    port map (
            O => \N__11100\,
            I => \N__11094\
        );

    \I__2063\ : CascadeBuf
    port map (
            O => \N__11097\,
            I => \N__11091\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__11094\,
            I => \N__11088\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__11091\,
            I => \N__11085\
        );

    \I__2060\ : CascadeBuf
    port map (
            O => \N__11088\,
            I => \N__11082\
        );

    \I__2059\ : CascadeBuf
    port map (
            O => \N__11085\,
            I => \N__11079\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__11082\,
            I => \N__11076\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__11079\,
            I => \N__11073\
        );

    \I__2056\ : CascadeBuf
    port map (
            O => \N__11076\,
            I => \N__11070\
        );

    \I__2055\ : CascadeBuf
    port map (
            O => \N__11073\,
            I => \N__11067\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__11070\,
            I => \N__11064\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__11067\,
            I => \N__11061\
        );

    \I__2052\ : CascadeBuf
    port map (
            O => \N__11064\,
            I => \N__11058\
        );

    \I__2051\ : CascadeBuf
    port map (
            O => \N__11061\,
            I => \N__11055\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__11058\,
            I => \N__11052\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__11055\,
            I => \N__11049\
        );

    \I__2048\ : CascadeBuf
    port map (
            O => \N__11052\,
            I => \N__11046\
        );

    \I__2047\ : CascadeBuf
    port map (
            O => \N__11049\,
            I => \N__11043\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__11046\,
            I => \N__11040\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__11043\,
            I => \N__11037\
        );

    \I__2044\ : CascadeBuf
    port map (
            O => \N__11040\,
            I => \N__11034\
        );

    \I__2043\ : CascadeBuf
    port map (
            O => \N__11037\,
            I => \N__11031\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__11034\,
            I => \N__11028\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__11031\,
            I => \N__11025\
        );

    \I__2040\ : CascadeBuf
    port map (
            O => \N__11028\,
            I => \N__11022\
        );

    \I__2039\ : CascadeBuf
    port map (
            O => \N__11025\,
            I => \N__11019\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__11022\,
            I => \N__11016\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__11019\,
            I => \N__11013\
        );

    \I__2036\ : CascadeBuf
    port map (
            O => \N__11016\,
            I => \N__11010\
        );

    \I__2035\ : CascadeBuf
    port map (
            O => \N__11013\,
            I => \N__11007\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__11010\,
            I => \N__11004\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__11007\,
            I => \N__11001\
        );

    \I__2032\ : CascadeBuf
    port map (
            O => \N__11004\,
            I => \N__10998\
        );

    \I__2031\ : CascadeBuf
    port map (
            O => \N__11001\,
            I => \N__10995\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__10998\,
            I => \N__10992\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__10995\,
            I => \N__10989\
        );

    \I__2028\ : CascadeBuf
    port map (
            O => \N__10992\,
            I => \N__10986\
        );

    \I__2027\ : CascadeBuf
    port map (
            O => \N__10989\,
            I => \N__10983\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__10986\,
            I => \N__10980\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__10983\,
            I => \N__10977\
        );

    \I__2024\ : CascadeBuf
    port map (
            O => \N__10980\,
            I => \N__10974\
        );

    \I__2023\ : CascadeBuf
    port map (
            O => \N__10977\,
            I => \N__10971\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__10974\,
            I => \N__10968\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__10971\,
            I => \N__10965\
        );

    \I__2020\ : CascadeBuf
    port map (
            O => \N__10968\,
            I => \N__10962\
        );

    \I__2019\ : CascadeBuf
    port map (
            O => \N__10965\,
            I => \N__10959\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__10962\,
            I => \N__10956\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__10959\,
            I => \N__10953\
        );

    \I__2016\ : CascadeBuf
    port map (
            O => \N__10956\,
            I => \N__10950\
        );

    \I__2015\ : CascadeBuf
    port map (
            O => \N__10953\,
            I => \N__10947\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__10950\,
            I => \N__10944\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__10947\,
            I => \N__10941\
        );

    \I__2012\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10938\
        );

    \I__2011\ : InMux
    port map (
            O => \N__10941\,
            I => \N__10935\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__10938\,
            I => \N__10932\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__10935\,
            I => \N__10929\
        );

    \I__2008\ : Sp12to4
    port map (
            O => \N__10932\,
            I => \N__10926\
        );

    \I__2007\ : Span12Mux_s8_h
    port map (
            O => \N__10929\,
            I => \N__10923\
        );

    \I__2006\ : Span12Mux_s11_h
    port map (
            O => \N__10926\,
            I => \N__10920\
        );

    \I__2005\ : Span12Mux_v
    port map (
            O => \N__10923\,
            I => \N__10915\
        );

    \I__2004\ : Span12Mux_v
    port map (
            O => \N__10920\,
            I => \N__10915\
        );

    \I__2003\ : Odrv12
    port map (
            O => \N__10915\,
            I => n19
        );

    \I__2002\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10906\
        );

    \I__2001\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10906\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__10906\,
            I => \transmit_module.n379\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__10903\,
            I => \N__10899\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__10902\,
            I => \N__10895\
        );

    \I__1997\ : InMux
    port map (
            O => \N__10899\,
            I => \N__10890\
        );

    \I__1996\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10890\
        );

    \I__1995\ : InMux
    port map (
            O => \N__10895\,
            I => \N__10887\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__10890\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__10887\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__1992\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10877\
        );

    \I__1991\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10874\
        );

    \I__1990\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10871\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__10877\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__10874\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__10871\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__10864\,
            I => \N__10861\
        );

    \I__1985\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10857\
        );

    \I__1984\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10854\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__10857\,
            I => \transmit_module.n380\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__10854\,
            I => \transmit_module.n380\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__10849\,
            I => \N__10846\
        );

    \I__1980\ : CascadeBuf
    port map (
            O => \N__10846\,
            I => \N__10842\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__10845\,
            I => \N__10839\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__10842\,
            I => \N__10836\
        );

    \I__1977\ : CascadeBuf
    port map (
            O => \N__10839\,
            I => \N__10833\
        );

    \I__1976\ : CascadeBuf
    port map (
            O => \N__10836\,
            I => \N__10830\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__10833\,
            I => \N__10827\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__10830\,
            I => \N__10824\
        );

    \I__1973\ : CascadeBuf
    port map (
            O => \N__10827\,
            I => \N__10821\
        );

    \I__1972\ : CascadeBuf
    port map (
            O => \N__10824\,
            I => \N__10818\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__10821\,
            I => \N__10815\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__10818\,
            I => \N__10812\
        );

    \I__1969\ : CascadeBuf
    port map (
            O => \N__10815\,
            I => \N__10809\
        );

    \I__1968\ : CascadeBuf
    port map (
            O => \N__10812\,
            I => \N__10806\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__10809\,
            I => \N__10803\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__10806\,
            I => \N__10800\
        );

    \I__1965\ : CascadeBuf
    port map (
            O => \N__10803\,
            I => \N__10797\
        );

    \I__1964\ : CascadeBuf
    port map (
            O => \N__10800\,
            I => \N__10794\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__10797\,
            I => \N__10791\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__10794\,
            I => \N__10788\
        );

    \I__1961\ : CascadeBuf
    port map (
            O => \N__10791\,
            I => \N__10785\
        );

    \I__1960\ : CascadeBuf
    port map (
            O => \N__10788\,
            I => \N__10782\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__10785\,
            I => \N__10779\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__10782\,
            I => \N__10776\
        );

    \I__1957\ : CascadeBuf
    port map (
            O => \N__10779\,
            I => \N__10773\
        );

    \I__1956\ : CascadeBuf
    port map (
            O => \N__10776\,
            I => \N__10770\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__10773\,
            I => \N__10767\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__10770\,
            I => \N__10764\
        );

    \I__1953\ : CascadeBuf
    port map (
            O => \N__10767\,
            I => \N__10761\
        );

    \I__1952\ : CascadeBuf
    port map (
            O => \N__10764\,
            I => \N__10758\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__10761\,
            I => \N__10755\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__10758\,
            I => \N__10752\
        );

    \I__1949\ : CascadeBuf
    port map (
            O => \N__10755\,
            I => \N__10749\
        );

    \I__1948\ : CascadeBuf
    port map (
            O => \N__10752\,
            I => \N__10746\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__10749\,
            I => \N__10743\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__10746\,
            I => \N__10740\
        );

    \I__1945\ : CascadeBuf
    port map (
            O => \N__10743\,
            I => \N__10737\
        );

    \I__1944\ : CascadeBuf
    port map (
            O => \N__10740\,
            I => \N__10734\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__10737\,
            I => \N__10731\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__10734\,
            I => \N__10728\
        );

    \I__1941\ : CascadeBuf
    port map (
            O => \N__10731\,
            I => \N__10725\
        );

    \I__1940\ : CascadeBuf
    port map (
            O => \N__10728\,
            I => \N__10722\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__10725\,
            I => \N__10719\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__10722\,
            I => \N__10716\
        );

    \I__1937\ : CascadeBuf
    port map (
            O => \N__10719\,
            I => \N__10713\
        );

    \I__1936\ : CascadeBuf
    port map (
            O => \N__10716\,
            I => \N__10710\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__10713\,
            I => \N__10707\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__10710\,
            I => \N__10704\
        );

    \I__1933\ : CascadeBuf
    port map (
            O => \N__10707\,
            I => \N__10701\
        );

    \I__1932\ : CascadeBuf
    port map (
            O => \N__10704\,
            I => \N__10698\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__10698\,
            I => \N__10692\
        );

    \I__1929\ : CascadeBuf
    port map (
            O => \N__10695\,
            I => \N__10689\
        );

    \I__1928\ : CascadeBuf
    port map (
            O => \N__10692\,
            I => \N__10686\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__10689\,
            I => \N__10683\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__10686\,
            I => \N__10680\
        );

    \I__1925\ : CascadeBuf
    port map (
            O => \N__10683\,
            I => \N__10677\
        );

    \I__1924\ : CascadeBuf
    port map (
            O => \N__10680\,
            I => \N__10674\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__10677\,
            I => \N__10671\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__10674\,
            I => \N__10668\
        );

    \I__1921\ : CascadeBuf
    port map (
            O => \N__10671\,
            I => \N__10665\
        );

    \I__1920\ : InMux
    port map (
            O => \N__10668\,
            I => \N__10662\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__10665\,
            I => \N__10659\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__10662\,
            I => \N__10656\
        );

    \I__1917\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10653\
        );

    \I__1916\ : Span12Mux_h
    port map (
            O => \N__10656\,
            I => \N__10650\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__10653\,
            I => \N__10647\
        );

    \I__1914\ : Span12Mux_v
    port map (
            O => \N__10650\,
            I => \N__10642\
        );

    \I__1913\ : Span12Mux_v
    port map (
            O => \N__10647\,
            I => \N__10642\
        );

    \I__1912\ : Odrv12
    port map (
            O => \N__10642\,
            I => n20
        );

    \I__1911\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10636\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__10636\,
            I => \N__10631\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__10635\,
            I => \N__10628\
        );

    \I__1908\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10625\
        );

    \I__1907\ : Span4Mux_v
    port map (
            O => \N__10631\,
            I => \N__10622\
        );

    \I__1906\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10619\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__10625\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__10622\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__10619\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__10612\,
            I => \N__10609\
        );

    \I__1901\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10605\
        );

    \I__1900\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10602\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__10605\,
            I => \transmit_module.n378\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__10602\,
            I => \transmit_module.n378\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__10597\,
            I => \N__10594\
        );

    \I__1896\ : CascadeBuf
    port map (
            O => \N__10594\,
            I => \N__10590\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__10593\,
            I => \N__10587\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__10590\,
            I => \N__10584\
        );

    \I__1893\ : CascadeBuf
    port map (
            O => \N__10587\,
            I => \N__10581\
        );

    \I__1892\ : CascadeBuf
    port map (
            O => \N__10584\,
            I => \N__10578\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__10581\,
            I => \N__10575\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__10578\,
            I => \N__10572\
        );

    \I__1889\ : CascadeBuf
    port map (
            O => \N__10575\,
            I => \N__10569\
        );

    \I__1888\ : CascadeBuf
    port map (
            O => \N__10572\,
            I => \N__10566\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__10569\,
            I => \N__10563\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__10566\,
            I => \N__10560\
        );

    \I__1885\ : CascadeBuf
    port map (
            O => \N__10563\,
            I => \N__10557\
        );

    \I__1884\ : CascadeBuf
    port map (
            O => \N__10560\,
            I => \N__10554\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__10557\,
            I => \N__10551\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__10554\,
            I => \N__10548\
        );

    \I__1881\ : CascadeBuf
    port map (
            O => \N__10551\,
            I => \N__10545\
        );

    \I__1880\ : CascadeBuf
    port map (
            O => \N__10548\,
            I => \N__10542\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__10545\,
            I => \N__10539\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__10542\,
            I => \N__10536\
        );

    \I__1877\ : CascadeBuf
    port map (
            O => \N__10539\,
            I => \N__10533\
        );

    \I__1876\ : CascadeBuf
    port map (
            O => \N__10536\,
            I => \N__10530\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__10533\,
            I => \N__10527\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__10530\,
            I => \N__10524\
        );

    \I__1873\ : CascadeBuf
    port map (
            O => \N__10527\,
            I => \N__10521\
        );

    \I__1872\ : CascadeBuf
    port map (
            O => \N__10524\,
            I => \N__10518\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__10521\,
            I => \N__10515\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__10518\,
            I => \N__10512\
        );

    \I__1869\ : CascadeBuf
    port map (
            O => \N__10515\,
            I => \N__10509\
        );

    \I__1868\ : CascadeBuf
    port map (
            O => \N__10512\,
            I => \N__10506\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__10509\,
            I => \N__10503\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__10506\,
            I => \N__10500\
        );

    \I__1865\ : CascadeBuf
    port map (
            O => \N__10503\,
            I => \N__10497\
        );

    \I__1864\ : CascadeBuf
    port map (
            O => \N__10500\,
            I => \N__10494\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__10497\,
            I => \N__10491\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__10494\,
            I => \N__10488\
        );

    \I__1861\ : CascadeBuf
    port map (
            O => \N__10491\,
            I => \N__10485\
        );

    \I__1860\ : CascadeBuf
    port map (
            O => \N__10488\,
            I => \N__10482\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__10485\,
            I => \N__10479\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__10482\,
            I => \N__10476\
        );

    \I__1857\ : CascadeBuf
    port map (
            O => \N__10479\,
            I => \N__10473\
        );

    \I__1856\ : CascadeBuf
    port map (
            O => \N__10476\,
            I => \N__10470\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__10473\,
            I => \N__10467\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__10470\,
            I => \N__10464\
        );

    \I__1853\ : CascadeBuf
    port map (
            O => \N__10467\,
            I => \N__10461\
        );

    \I__1852\ : CascadeBuf
    port map (
            O => \N__10464\,
            I => \N__10458\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__10461\,
            I => \N__10455\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__10458\,
            I => \N__10452\
        );

    \I__1849\ : CascadeBuf
    port map (
            O => \N__10455\,
            I => \N__10449\
        );

    \I__1848\ : CascadeBuf
    port map (
            O => \N__10452\,
            I => \N__10446\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__10449\,
            I => \N__10443\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__10446\,
            I => \N__10440\
        );

    \I__1845\ : CascadeBuf
    port map (
            O => \N__10443\,
            I => \N__10437\
        );

    \I__1844\ : CascadeBuf
    port map (
            O => \N__10440\,
            I => \N__10434\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__10437\,
            I => \N__10431\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__10434\,
            I => \N__10428\
        );

    \I__1841\ : CascadeBuf
    port map (
            O => \N__10431\,
            I => \N__10425\
        );

    \I__1840\ : CascadeBuf
    port map (
            O => \N__10428\,
            I => \N__10422\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__10425\,
            I => \N__10419\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__10422\,
            I => \N__10416\
        );

    \I__1837\ : CascadeBuf
    port map (
            O => \N__10419\,
            I => \N__10413\
        );

    \I__1836\ : InMux
    port map (
            O => \N__10416\,
            I => \N__10410\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__10413\,
            I => \N__10407\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__10410\,
            I => \N__10404\
        );

    \I__1833\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10401\
        );

    \I__1832\ : Sp12to4
    port map (
            O => \N__10404\,
            I => \N__10398\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__10401\,
            I => \N__10395\
        );

    \I__1830\ : Span12Mux_h
    port map (
            O => \N__10398\,
            I => \N__10392\
        );

    \I__1829\ : Span12Mux_v
    port map (
            O => \N__10395\,
            I => \N__10387\
        );

    \I__1828\ : Span12Mux_v
    port map (
            O => \N__10392\,
            I => \N__10387\
        );

    \I__1827\ : Odrv12
    port map (
            O => \N__10387\,
            I => n18
        );

    \I__1826\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10381\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__10381\,
            I => \N__10378\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__10378\,
            I => \line_buffer.n3104\
        );

    \I__1823\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10372\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__10372\,
            I => \N__10369\
        );

    \I__1821\ : Odrv12
    port map (
            O => \N__10369\,
            I => \TX_DATA_6\
        );

    \I__1820\ : IoInMux
    port map (
            O => \N__10366\,
            I => \N__10363\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__10363\,
            I => \N__10360\
        );

    \I__1818\ : IoSpan4Mux
    port map (
            O => \N__10360\,
            I => \N__10357\
        );

    \I__1817\ : Span4Mux_s0_v
    port map (
            O => \N__10357\,
            I => \N__10354\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__10354\,
            I => \GB_BUFFER_TVP_CLK_c_THRU_CO\
        );

    \I__1815\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10348\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__10348\,
            I => \receive_module.old_VS\
        );

    \I__1813\ : CEMux
    port map (
            O => \N__10345\,
            I => \N__10342\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__10342\,
            I => \N__10338\
        );

    \I__1811\ : CEMux
    port map (
            O => \N__10341\,
            I => \N__10335\
        );

    \I__1810\ : Span4Mux_h
    port map (
            O => \N__10338\,
            I => \N__10331\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__10335\,
            I => \N__10328\
        );

    \I__1808\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10325\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__10331\,
            I => \receive_module.n252\
        );

    \I__1806\ : Odrv12
    port map (
            O => \N__10328\,
            I => \receive_module.n252\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__10325\,
            I => \receive_module.n252\
        );

    \I__1804\ : IoInMux
    port map (
            O => \N__10318\,
            I => \N__10315\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__10315\,
            I => \N__10312\
        );

    \I__1802\ : Span4Mux_s3_h
    port map (
            O => \N__10312\,
            I => \N__10307\
        );

    \I__1801\ : IoInMux
    port map (
            O => \N__10311\,
            I => \N__10304\
        );

    \I__1800\ : IoInMux
    port map (
            O => \N__10310\,
            I => \N__10301\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__10307\,
            I => \N__10298\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__10304\,
            I => \N__10295\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__10301\,
            I => \N__10292\
        );

    \I__1796\ : Span4Mux_h
    port map (
            O => \N__10298\,
            I => \N__10289\
        );

    \I__1795\ : Span4Mux_s3_v
    port map (
            O => \N__10295\,
            I => \N__10286\
        );

    \I__1794\ : Span12Mux_s3_v
    port map (
            O => \N__10292\,
            I => \N__10283\
        );

    \I__1793\ : Span4Mux_h
    port map (
            O => \N__10289\,
            I => \N__10280\
        );

    \I__1792\ : Sp12to4
    port map (
            O => \N__10286\,
            I => \N__10277\
        );

    \I__1791\ : Span12Mux_h
    port map (
            O => \N__10283\,
            I => \N__10270\
        );

    \I__1790\ : Sp12to4
    port map (
            O => \N__10280\,
            I => \N__10270\
        );

    \I__1789\ : Span12Mux_h
    port map (
            O => \N__10277\,
            I => \N__10270\
        );

    \I__1788\ : Span12Mux_v
    port map (
            O => \N__10270\,
            I => \N__10267\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__10267\,
            I => n1950
        );

    \I__1786\ : IoInMux
    port map (
            O => \N__10264\,
            I => \N__10261\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__10261\,
            I => \N__10258\
        );

    \I__1784\ : IoSpan4Mux
    port map (
            O => \N__10258\,
            I => \N__10253\
        );

    \I__1783\ : IoInMux
    port map (
            O => \N__10257\,
            I => \N__10250\
        );

    \I__1782\ : IoInMux
    port map (
            O => \N__10256\,
            I => \N__10247\
        );

    \I__1781\ : Span4Mux_s1_v
    port map (
            O => \N__10253\,
            I => \N__10244\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__10250\,
            I => \N__10241\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__10247\,
            I => \N__10238\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__10244\,
            I => \N__10233\
        );

    \I__1777\ : Span4Mux_s3_h
    port map (
            O => \N__10241\,
            I => \N__10233\
        );

    \I__1776\ : Span4Mux_s3_v
    port map (
            O => \N__10238\,
            I => \N__10230\
        );

    \I__1775\ : Sp12to4
    port map (
            O => \N__10233\,
            I => \N__10227\
        );

    \I__1774\ : Span4Mux_v
    port map (
            O => \N__10230\,
            I => \N__10224\
        );

    \I__1773\ : Span12Mux_s7_v
    port map (
            O => \N__10227\,
            I => \N__10221\
        );

    \I__1772\ : Span4Mux_v
    port map (
            O => \N__10224\,
            I => \N__10218\
        );

    \I__1771\ : Span12Mux_h
    port map (
            O => \N__10221\,
            I => \N__10215\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__10218\,
            I => \N__10212\
        );

    \I__1769\ : Odrv12
    port map (
            O => \N__10215\,
            I => n1954
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__10212\,
            I => n1954
        );

    \I__1767\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10204\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__10204\,
            I => \N__10201\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__10201\,
            I => \TX_DATA_3\
        );

    \I__1764\ : IoInMux
    port map (
            O => \N__10198\,
            I => \N__10193\
        );

    \I__1763\ : IoInMux
    port map (
            O => \N__10197\,
            I => \N__10190\
        );

    \I__1762\ : IoInMux
    port map (
            O => \N__10196\,
            I => \N__10187\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__10193\,
            I => \N__10184\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__10190\,
            I => \N__10181\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10178\
        );

    \I__1758\ : Span4Mux_s3_v
    port map (
            O => \N__10184\,
            I => \N__10175\
        );

    \I__1757\ : Span4Mux_s3_v
    port map (
            O => \N__10181\,
            I => \N__10172\
        );

    \I__1756\ : Span4Mux_s3_h
    port map (
            O => \N__10178\,
            I => \N__10169\
        );

    \I__1755\ : Sp12to4
    port map (
            O => \N__10175\,
            I => \N__10166\
        );

    \I__1754\ : Sp12to4
    port map (
            O => \N__10172\,
            I => \N__10163\
        );

    \I__1753\ : Sp12to4
    port map (
            O => \N__10169\,
            I => \N__10160\
        );

    \I__1752\ : Span12Mux_s8_h
    port map (
            O => \N__10166\,
            I => \N__10157\
        );

    \I__1751\ : Span12Mux_s11_h
    port map (
            O => \N__10163\,
            I => \N__10154\
        );

    \I__1750\ : Span12Mux_v
    port map (
            O => \N__10160\,
            I => \N__10151\
        );

    \I__1749\ : Span12Mux_v
    port map (
            O => \N__10157\,
            I => \N__10146\
        );

    \I__1748\ : Span12Mux_v
    port map (
            O => \N__10154\,
            I => \N__10146\
        );

    \I__1747\ : Span12Mux_h
    port map (
            O => \N__10151\,
            I => \N__10143\
        );

    \I__1746\ : Odrv12
    port map (
            O => \N__10146\,
            I => n1952
        );

    \I__1745\ : Odrv12
    port map (
            O => \N__10143\,
            I => n1952
        );

    \I__1744\ : IoInMux
    port map (
            O => \N__10138\,
            I => \N__10134\
        );

    \I__1743\ : IoInMux
    port map (
            O => \N__10137\,
            I => \N__10131\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__10134\,
            I => \N__10128\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__10131\,
            I => \N__10124\
        );

    \I__1740\ : IoSpan4Mux
    port map (
            O => \N__10128\,
            I => \N__10121\
        );

    \I__1739\ : IoInMux
    port map (
            O => \N__10127\,
            I => \N__10118\
        );

    \I__1738\ : IoSpan4Mux
    port map (
            O => \N__10124\,
            I => \N__10115\
        );

    \I__1737\ : Span4Mux_s3_v
    port map (
            O => \N__10121\,
            I => \N__10112\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__10118\,
            I => \N__10109\
        );

    \I__1735\ : Span4Mux_s3_v
    port map (
            O => \N__10115\,
            I => \N__10106\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__10112\,
            I => \N__10101\
        );

    \I__1733\ : Span4Mux_s3_h
    port map (
            O => \N__10109\,
            I => \N__10101\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__10106\,
            I => \N__10098\
        );

    \I__1731\ : Sp12to4
    port map (
            O => \N__10101\,
            I => \N__10095\
        );

    \I__1730\ : Sp12to4
    port map (
            O => \N__10098\,
            I => \N__10092\
        );

    \I__1729\ : Span12Mux_v
    port map (
            O => \N__10095\,
            I => \N__10089\
        );

    \I__1728\ : Span12Mux_v
    port map (
            O => \N__10092\,
            I => \N__10084\
        );

    \I__1727\ : Span12Mux_h
    port map (
            O => \N__10089\,
            I => \N__10084\
        );

    \I__1726\ : Odrv12
    port map (
            O => \N__10084\,
            I => n1951
        );

    \I__1725\ : IoInMux
    port map (
            O => \N__10081\,
            I => \N__10078\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__10078\,
            I => \N__10073\
        );

    \I__1723\ : IoInMux
    port map (
            O => \N__10077\,
            I => \N__10070\
        );

    \I__1722\ : IoInMux
    port map (
            O => \N__10076\,
            I => \N__10067\
        );

    \I__1721\ : IoSpan4Mux
    port map (
            O => \N__10073\,
            I => \N__10064\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__10070\,
            I => \N__10061\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__10067\,
            I => \N__10058\
        );

    \I__1718\ : Span4Mux_s1_h
    port map (
            O => \N__10064\,
            I => \N__10055\
        );

    \I__1717\ : Span4Mux_s3_v
    port map (
            O => \N__10061\,
            I => \N__10052\
        );

    \I__1716\ : Span12Mux_s3_v
    port map (
            O => \N__10058\,
            I => \N__10049\
        );

    \I__1715\ : Sp12to4
    port map (
            O => \N__10055\,
            I => \N__10046\
        );

    \I__1714\ : Span4Mux_h
    port map (
            O => \N__10052\,
            I => \N__10043\
        );

    \I__1713\ : Span12Mux_v
    port map (
            O => \N__10049\,
            I => \N__10040\
        );

    \I__1712\ : Span12Mux_v
    port map (
            O => \N__10046\,
            I => \N__10037\
        );

    \I__1711\ : Sp12to4
    port map (
            O => \N__10043\,
            I => \N__10034\
        );

    \I__1710\ : Span12Mux_h
    port map (
            O => \N__10040\,
            I => \N__10031\
        );

    \I__1709\ : Span12Mux_h
    port map (
            O => \N__10037\,
            I => \N__10026\
        );

    \I__1708\ : Span12Mux_v
    port map (
            O => \N__10034\,
            I => \N__10026\
        );

    \I__1707\ : Odrv12
    port map (
            O => \N__10031\,
            I => n1949
        );

    \I__1706\ : Odrv12
    port map (
            O => \N__10026\,
            I => n1949
        );

    \I__1705\ : IoInMux
    port map (
            O => \N__10021\,
            I => \N__10016\
        );

    \I__1704\ : IoInMux
    port map (
            O => \N__10020\,
            I => \N__10013\
        );

    \I__1703\ : IoInMux
    port map (
            O => \N__10019\,
            I => \N__10010\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__10016\,
            I => \N__10007\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__10013\,
            I => \N__10004\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__10010\,
            I => \N__10001\
        );

    \I__1699\ : Span4Mux_s3_v
    port map (
            O => \N__10007\,
            I => \N__9998\
        );

    \I__1698\ : Span4Mux_s0_h
    port map (
            O => \N__10004\,
            I => \N__9995\
        );

    \I__1697\ : Span4Mux_s3_v
    port map (
            O => \N__10001\,
            I => \N__9992\
        );

    \I__1696\ : Sp12to4
    port map (
            O => \N__9998\,
            I => \N__9989\
        );

    \I__1695\ : Sp12to4
    port map (
            O => \N__9995\,
            I => \N__9986\
        );

    \I__1694\ : Sp12to4
    port map (
            O => \N__9992\,
            I => \N__9983\
        );

    \I__1693\ : Span12Mux_s7_h
    port map (
            O => \N__9989\,
            I => \N__9980\
        );

    \I__1692\ : Span12Mux_v
    port map (
            O => \N__9986\,
            I => \N__9977\
        );

    \I__1691\ : Span12Mux_h
    port map (
            O => \N__9983\,
            I => \N__9974\
        );

    \I__1690\ : Span12Mux_v
    port map (
            O => \N__9980\,
            I => \N__9967\
        );

    \I__1689\ : Span12Mux_h
    port map (
            O => \N__9977\,
            I => \N__9967\
        );

    \I__1688\ : Span12Mux_v
    port map (
            O => \N__9974\,
            I => \N__9967\
        );

    \I__1687\ : Odrv12
    port map (
            O => \N__9967\,
            I => \ADV_B_c\
        );

    \I__1686\ : InMux
    port map (
            O => \N__9964\,
            I => \transmit_module.n2752\
        );

    \I__1685\ : CEMux
    port map (
            O => \N__9961\,
            I => \N__9957\
        );

    \I__1684\ : CEMux
    port map (
            O => \N__9960\,
            I => \N__9952\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__9957\,
            I => \N__9949\
        );

    \I__1682\ : CEMux
    port map (
            O => \N__9956\,
            I => \N__9946\
        );

    \I__1681\ : CEMux
    port map (
            O => \N__9955\,
            I => \N__9943\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__9952\,
            I => \transmit_module.n2200\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__9949\,
            I => \transmit_module.n2200\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__9946\,
            I => \transmit_module.n2200\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__9943\,
            I => \transmit_module.n2200\
        );

    \I__1676\ : IoInMux
    port map (
            O => \N__9934\,
            I => \N__9931\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__9931\,
            I => \N__9926\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__9930\,
            I => \N__9923\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__9929\,
            I => \N__9919\
        );

    \I__1672\ : Span12Mux_s5_h
    port map (
            O => \N__9926\,
            I => \N__9916\
        );

    \I__1671\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9913\
        );

    \I__1670\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9910\
        );

    \I__1669\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9907\
        );

    \I__1668\ : Odrv12
    port map (
            O => \N__9916\,
            I => \DEBUG_c_6\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__9913\,
            I => \DEBUG_c_6\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__9910\,
            I => \DEBUG_c_6\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__9907\,
            I => \DEBUG_c_6\
        );

    \I__1664\ : InMux
    port map (
            O => \N__9898\,
            I => \N__9894\
        );

    \I__1663\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9891\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__9894\,
            I => \N__9888\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__9891\,
            I => \transmit_module.n382\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__9888\,
            I => \transmit_module.n382\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__9883\,
            I => \N__9879\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__9882\,
            I => \N__9876\
        );

    \I__1657\ : CascadeBuf
    port map (
            O => \N__9879\,
            I => \N__9873\
        );

    \I__1656\ : CascadeBuf
    port map (
            O => \N__9876\,
            I => \N__9870\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__9873\,
            I => \N__9867\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__9870\,
            I => \N__9864\
        );

    \I__1653\ : CascadeBuf
    port map (
            O => \N__9867\,
            I => \N__9861\
        );

    \I__1652\ : CascadeBuf
    port map (
            O => \N__9864\,
            I => \N__9858\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__9861\,
            I => \N__9855\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__9858\,
            I => \N__9852\
        );

    \I__1649\ : CascadeBuf
    port map (
            O => \N__9855\,
            I => \N__9849\
        );

    \I__1648\ : CascadeBuf
    port map (
            O => \N__9852\,
            I => \N__9846\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__9849\,
            I => \N__9843\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__9846\,
            I => \N__9840\
        );

    \I__1645\ : CascadeBuf
    port map (
            O => \N__9843\,
            I => \N__9837\
        );

    \I__1644\ : CascadeBuf
    port map (
            O => \N__9840\,
            I => \N__9834\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__9837\,
            I => \N__9831\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__9834\,
            I => \N__9828\
        );

    \I__1641\ : CascadeBuf
    port map (
            O => \N__9831\,
            I => \N__9825\
        );

    \I__1640\ : CascadeBuf
    port map (
            O => \N__9828\,
            I => \N__9822\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__9825\,
            I => \N__9819\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__9822\,
            I => \N__9816\
        );

    \I__1637\ : CascadeBuf
    port map (
            O => \N__9819\,
            I => \N__9813\
        );

    \I__1636\ : CascadeBuf
    port map (
            O => \N__9816\,
            I => \N__9810\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__9813\,
            I => \N__9807\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__9810\,
            I => \N__9804\
        );

    \I__1633\ : CascadeBuf
    port map (
            O => \N__9807\,
            I => \N__9801\
        );

    \I__1632\ : CascadeBuf
    port map (
            O => \N__9804\,
            I => \N__9798\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__9801\,
            I => \N__9795\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__9798\,
            I => \N__9792\
        );

    \I__1629\ : CascadeBuf
    port map (
            O => \N__9795\,
            I => \N__9789\
        );

    \I__1628\ : CascadeBuf
    port map (
            O => \N__9792\,
            I => \N__9786\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__9789\,
            I => \N__9783\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__9786\,
            I => \N__9780\
        );

    \I__1625\ : CascadeBuf
    port map (
            O => \N__9783\,
            I => \N__9777\
        );

    \I__1624\ : CascadeBuf
    port map (
            O => \N__9780\,
            I => \N__9774\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__9777\,
            I => \N__9771\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__9774\,
            I => \N__9768\
        );

    \I__1621\ : CascadeBuf
    port map (
            O => \N__9771\,
            I => \N__9765\
        );

    \I__1620\ : CascadeBuf
    port map (
            O => \N__9768\,
            I => \N__9762\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__9765\,
            I => \N__9759\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__9762\,
            I => \N__9756\
        );

    \I__1617\ : CascadeBuf
    port map (
            O => \N__9759\,
            I => \N__9753\
        );

    \I__1616\ : CascadeBuf
    port map (
            O => \N__9756\,
            I => \N__9750\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__9753\,
            I => \N__9747\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__9750\,
            I => \N__9744\
        );

    \I__1613\ : CascadeBuf
    port map (
            O => \N__9747\,
            I => \N__9741\
        );

    \I__1612\ : CascadeBuf
    port map (
            O => \N__9744\,
            I => \N__9738\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__9741\,
            I => \N__9735\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__9738\,
            I => \N__9732\
        );

    \I__1609\ : CascadeBuf
    port map (
            O => \N__9735\,
            I => \N__9729\
        );

    \I__1608\ : CascadeBuf
    port map (
            O => \N__9732\,
            I => \N__9726\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__9729\,
            I => \N__9723\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__9726\,
            I => \N__9720\
        );

    \I__1605\ : CascadeBuf
    port map (
            O => \N__9723\,
            I => \N__9717\
        );

    \I__1604\ : CascadeBuf
    port map (
            O => \N__9720\,
            I => \N__9714\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__9717\,
            I => \N__9711\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__9714\,
            I => \N__9708\
        );

    \I__1601\ : CascadeBuf
    port map (
            O => \N__9711\,
            I => \N__9705\
        );

    \I__1600\ : CascadeBuf
    port map (
            O => \N__9708\,
            I => \N__9702\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__9705\,
            I => \N__9699\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__9702\,
            I => \N__9696\
        );

    \I__1597\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9693\
        );

    \I__1596\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9690\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__9693\,
            I => \N__9687\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__9690\,
            I => \N__9684\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__9687\,
            I => \N__9681\
        );

    \I__1592\ : Span4Mux_h
    port map (
            O => \N__9684\,
            I => \N__9678\
        );

    \I__1591\ : Span4Mux_h
    port map (
            O => \N__9681\,
            I => \N__9675\
        );

    \I__1590\ : Sp12to4
    port map (
            O => \N__9678\,
            I => \N__9672\
        );

    \I__1589\ : Span4Mux_v
    port map (
            O => \N__9675\,
            I => \N__9669\
        );

    \I__1588\ : Span12Mux_v
    port map (
            O => \N__9672\,
            I => \N__9666\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__9669\,
            I => \N__9663\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__9666\,
            I => n22
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__9663\,
            I => n22
        );

    \I__1584\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9654\
        );

    \I__1583\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9651\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__9654\,
            I => \N__9648\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__9651\,
            I => \transmit_module.n383\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__9648\,
            I => \transmit_module.n383\
        );

    \I__1579\ : IoInMux
    port map (
            O => \N__9643\,
            I => \N__9640\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__9640\,
            I => \N__9637\
        );

    \I__1577\ : Span4Mux_s2_h
    port map (
            O => \N__9637\,
            I => \N__9634\
        );

    \I__1576\ : Span4Mux_h
    port map (
            O => \N__9634\,
            I => \N__9631\
        );

    \I__1575\ : Span4Mux_h
    port map (
            O => \N__9631\,
            I => \N__9627\
        );

    \I__1574\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9623\
        );

    \I__1573\ : Span4Mux_h
    port map (
            O => \N__9627\,
            I => \N__9619\
        );

    \I__1572\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9616\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__9623\,
            I => \N__9613\
        );

    \I__1570\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9610\
        );

    \I__1569\ : Odrv4
    port map (
            O => \N__9619\,
            I => \DEBUG_c_5\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__9616\,
            I => \DEBUG_c_5\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__9613\,
            I => \DEBUG_c_5\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__9610\,
            I => \DEBUG_c_5\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__9601\,
            I => \N__9597\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__9600\,
            I => \N__9594\
        );

    \I__1563\ : CascadeBuf
    port map (
            O => \N__9597\,
            I => \N__9591\
        );

    \I__1562\ : CascadeBuf
    port map (
            O => \N__9594\,
            I => \N__9588\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__9591\,
            I => \N__9585\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__9588\,
            I => \N__9582\
        );

    \I__1559\ : CascadeBuf
    port map (
            O => \N__9585\,
            I => \N__9579\
        );

    \I__1558\ : CascadeBuf
    port map (
            O => \N__9582\,
            I => \N__9576\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__9579\,
            I => \N__9573\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__9576\,
            I => \N__9570\
        );

    \I__1555\ : CascadeBuf
    port map (
            O => \N__9573\,
            I => \N__9567\
        );

    \I__1554\ : CascadeBuf
    port map (
            O => \N__9570\,
            I => \N__9564\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__9567\,
            I => \N__9561\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__9564\,
            I => \N__9558\
        );

    \I__1551\ : CascadeBuf
    port map (
            O => \N__9561\,
            I => \N__9555\
        );

    \I__1550\ : CascadeBuf
    port map (
            O => \N__9558\,
            I => \N__9552\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__9555\,
            I => \N__9549\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__9552\,
            I => \N__9546\
        );

    \I__1547\ : CascadeBuf
    port map (
            O => \N__9549\,
            I => \N__9543\
        );

    \I__1546\ : CascadeBuf
    port map (
            O => \N__9546\,
            I => \N__9540\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__9543\,
            I => \N__9537\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__9540\,
            I => \N__9534\
        );

    \I__1543\ : CascadeBuf
    port map (
            O => \N__9537\,
            I => \N__9531\
        );

    \I__1542\ : CascadeBuf
    port map (
            O => \N__9534\,
            I => \N__9528\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__9531\,
            I => \N__9525\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__9528\,
            I => \N__9522\
        );

    \I__1539\ : CascadeBuf
    port map (
            O => \N__9525\,
            I => \N__9519\
        );

    \I__1538\ : CascadeBuf
    port map (
            O => \N__9522\,
            I => \N__9516\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__9519\,
            I => \N__9513\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__9516\,
            I => \N__9510\
        );

    \I__1535\ : CascadeBuf
    port map (
            O => \N__9513\,
            I => \N__9507\
        );

    \I__1534\ : CascadeBuf
    port map (
            O => \N__9510\,
            I => \N__9504\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__9507\,
            I => \N__9501\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__9504\,
            I => \N__9498\
        );

    \I__1531\ : CascadeBuf
    port map (
            O => \N__9501\,
            I => \N__9495\
        );

    \I__1530\ : CascadeBuf
    port map (
            O => \N__9498\,
            I => \N__9492\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__9495\,
            I => \N__9489\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__9492\,
            I => \N__9486\
        );

    \I__1527\ : CascadeBuf
    port map (
            O => \N__9489\,
            I => \N__9483\
        );

    \I__1526\ : CascadeBuf
    port map (
            O => \N__9486\,
            I => \N__9480\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__9483\,
            I => \N__9477\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__9480\,
            I => \N__9474\
        );

    \I__1523\ : CascadeBuf
    port map (
            O => \N__9477\,
            I => \N__9471\
        );

    \I__1522\ : CascadeBuf
    port map (
            O => \N__9474\,
            I => \N__9468\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__9471\,
            I => \N__9465\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__9468\,
            I => \N__9462\
        );

    \I__1519\ : CascadeBuf
    port map (
            O => \N__9465\,
            I => \N__9459\
        );

    \I__1518\ : CascadeBuf
    port map (
            O => \N__9462\,
            I => \N__9456\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__9459\,
            I => \N__9453\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__9456\,
            I => \N__9450\
        );

    \I__1515\ : CascadeBuf
    port map (
            O => \N__9453\,
            I => \N__9447\
        );

    \I__1514\ : CascadeBuf
    port map (
            O => \N__9450\,
            I => \N__9444\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__9447\,
            I => \N__9441\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__9444\,
            I => \N__9438\
        );

    \I__1511\ : CascadeBuf
    port map (
            O => \N__9441\,
            I => \N__9435\
        );

    \I__1510\ : CascadeBuf
    port map (
            O => \N__9438\,
            I => \N__9432\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__9435\,
            I => \N__9429\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__9432\,
            I => \N__9426\
        );

    \I__1507\ : CascadeBuf
    port map (
            O => \N__9429\,
            I => \N__9423\
        );

    \I__1506\ : CascadeBuf
    port map (
            O => \N__9426\,
            I => \N__9420\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__9423\,
            I => \N__9417\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__9420\,
            I => \N__9414\
        );

    \I__1503\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9411\
        );

    \I__1502\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9408\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__9411\,
            I => \N__9405\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__9408\,
            I => \N__9402\
        );

    \I__1499\ : Span12Mux_s11_h
    port map (
            O => \N__9405\,
            I => \N__9399\
        );

    \I__1498\ : Span12Mux_s8_h
    port map (
            O => \N__9402\,
            I => \N__9396\
        );

    \I__1497\ : Span12Mux_v
    port map (
            O => \N__9399\,
            I => \N__9391\
        );

    \I__1496\ : Span12Mux_v
    port map (
            O => \N__9396\,
            I => \N__9391\
        );

    \I__1495\ : Odrv12
    port map (
            O => \N__9391\,
            I => n23
        );

    \I__1494\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9385\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__9385\,
            I => \N__9381\
        );

    \I__1492\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9378\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__9381\,
            I => \N__9375\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__9378\,
            I => \transmit_module.n384\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__9375\,
            I => \transmit_module.n384\
        );

    \I__1488\ : IoInMux
    port map (
            O => \N__9370\,
            I => \N__9367\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__9367\,
            I => \N__9363\
        );

    \I__1486\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9359\
        );

    \I__1485\ : Span12Mux_s9_h
    port map (
            O => \N__9363\,
            I => \N__9355\
        );

    \I__1484\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9352\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__9359\,
            I => \N__9349\
        );

    \I__1482\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9346\
        );

    \I__1481\ : Odrv12
    port map (
            O => \N__9355\,
            I => \DEBUG_c_4\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__9352\,
            I => \DEBUG_c_4\
        );

    \I__1479\ : Odrv12
    port map (
            O => \N__9349\,
            I => \DEBUG_c_4\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__9346\,
            I => \DEBUG_c_4\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__9337\,
            I => \N__9333\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__9336\,
            I => \N__9330\
        );

    \I__1475\ : CascadeBuf
    port map (
            O => \N__9333\,
            I => \N__9327\
        );

    \I__1474\ : CascadeBuf
    port map (
            O => \N__9330\,
            I => \N__9324\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__9327\,
            I => \N__9321\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__9324\,
            I => \N__9318\
        );

    \I__1471\ : CascadeBuf
    port map (
            O => \N__9321\,
            I => \N__9315\
        );

    \I__1470\ : CascadeBuf
    port map (
            O => \N__9318\,
            I => \N__9312\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__9315\,
            I => \N__9309\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__9312\,
            I => \N__9306\
        );

    \I__1467\ : CascadeBuf
    port map (
            O => \N__9309\,
            I => \N__9303\
        );

    \I__1466\ : CascadeBuf
    port map (
            O => \N__9306\,
            I => \N__9300\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__9303\,
            I => \N__9297\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__9300\,
            I => \N__9294\
        );

    \I__1463\ : CascadeBuf
    port map (
            O => \N__9297\,
            I => \N__9291\
        );

    \I__1462\ : CascadeBuf
    port map (
            O => \N__9294\,
            I => \N__9288\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__9291\,
            I => \N__9285\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__9288\,
            I => \N__9282\
        );

    \I__1459\ : CascadeBuf
    port map (
            O => \N__9285\,
            I => \N__9279\
        );

    \I__1458\ : CascadeBuf
    port map (
            O => \N__9282\,
            I => \N__9276\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__9279\,
            I => \N__9273\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__9276\,
            I => \N__9270\
        );

    \I__1455\ : CascadeBuf
    port map (
            O => \N__9273\,
            I => \N__9267\
        );

    \I__1454\ : CascadeBuf
    port map (
            O => \N__9270\,
            I => \N__9264\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__9267\,
            I => \N__9261\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__9264\,
            I => \N__9258\
        );

    \I__1451\ : CascadeBuf
    port map (
            O => \N__9261\,
            I => \N__9255\
        );

    \I__1450\ : CascadeBuf
    port map (
            O => \N__9258\,
            I => \N__9252\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__9255\,
            I => \N__9249\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__9252\,
            I => \N__9246\
        );

    \I__1447\ : CascadeBuf
    port map (
            O => \N__9249\,
            I => \N__9243\
        );

    \I__1446\ : CascadeBuf
    port map (
            O => \N__9246\,
            I => \N__9240\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__9243\,
            I => \N__9237\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__9240\,
            I => \N__9234\
        );

    \I__1443\ : CascadeBuf
    port map (
            O => \N__9237\,
            I => \N__9231\
        );

    \I__1442\ : CascadeBuf
    port map (
            O => \N__9234\,
            I => \N__9228\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__9231\,
            I => \N__9225\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__9228\,
            I => \N__9222\
        );

    \I__1439\ : CascadeBuf
    port map (
            O => \N__9225\,
            I => \N__9219\
        );

    \I__1438\ : CascadeBuf
    port map (
            O => \N__9222\,
            I => \N__9216\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__9219\,
            I => \N__9213\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__9216\,
            I => \N__9210\
        );

    \I__1435\ : CascadeBuf
    port map (
            O => \N__9213\,
            I => \N__9207\
        );

    \I__1434\ : CascadeBuf
    port map (
            O => \N__9210\,
            I => \N__9204\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__9207\,
            I => \N__9201\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__9204\,
            I => \N__9198\
        );

    \I__1431\ : CascadeBuf
    port map (
            O => \N__9201\,
            I => \N__9195\
        );

    \I__1430\ : CascadeBuf
    port map (
            O => \N__9198\,
            I => \N__9192\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__9195\,
            I => \N__9189\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__9192\,
            I => \N__9186\
        );

    \I__1427\ : CascadeBuf
    port map (
            O => \N__9189\,
            I => \N__9183\
        );

    \I__1426\ : CascadeBuf
    port map (
            O => \N__9186\,
            I => \N__9180\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__9183\,
            I => \N__9177\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__9180\,
            I => \N__9174\
        );

    \I__1423\ : CascadeBuf
    port map (
            O => \N__9177\,
            I => \N__9171\
        );

    \I__1422\ : CascadeBuf
    port map (
            O => \N__9174\,
            I => \N__9168\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__9171\,
            I => \N__9165\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__9168\,
            I => \N__9162\
        );

    \I__1419\ : CascadeBuf
    port map (
            O => \N__9165\,
            I => \N__9159\
        );

    \I__1418\ : CascadeBuf
    port map (
            O => \N__9162\,
            I => \N__9156\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__9159\,
            I => \N__9153\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__9156\,
            I => \N__9150\
        );

    \I__1415\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9147\
        );

    \I__1414\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9144\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__9147\,
            I => \N__9141\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__9144\,
            I => \N__9138\
        );

    \I__1411\ : Span12Mux_h
    port map (
            O => \N__9141\,
            I => \N__9133\
        );

    \I__1410\ : Span12Mux_h
    port map (
            O => \N__9138\,
            I => \N__9133\
        );

    \I__1409\ : Span12Mux_v
    port map (
            O => \N__9133\,
            I => \N__9130\
        );

    \I__1408\ : Odrv12
    port map (
            O => \N__9130\,
            I => n24
        );

    \I__1407\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9123\
        );

    \I__1406\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9120\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__9123\,
            I => \N__9117\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__9120\,
            I => \transmit_module.n386\
        );

    \I__1403\ : Odrv12
    port map (
            O => \N__9117\,
            I => \transmit_module.n386\
        );

    \I__1402\ : IoInMux
    port map (
            O => \N__9112\,
            I => \N__9109\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__1400\ : Span4Mux_s1_h
    port map (
            O => \N__9106\,
            I => \N__9103\
        );

    \I__1399\ : Sp12to4
    port map (
            O => \N__9103\,
            I => \N__9099\
        );

    \I__1398\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9096\
        );

    \I__1397\ : Span12Mux_v
    port map (
            O => \N__9099\,
            I => \N__9093\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__9096\,
            I => \N__9089\
        );

    \I__1395\ : Span12Mux_h
    port map (
            O => \N__9093\,
            I => \N__9085\
        );

    \I__1394\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9082\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__9089\,
            I => \N__9079\
        );

    \I__1392\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9076\
        );

    \I__1391\ : Odrv12
    port map (
            O => \N__9085\,
            I => \DEBUG_c_2\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__9082\,
            I => \DEBUG_c_2\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__9079\,
            I => \DEBUG_c_2\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__9076\,
            I => \DEBUG_c_2\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__9067\,
            I => \N__9064\
        );

    \I__1386\ : CascadeBuf
    port map (
            O => \N__9064\,
            I => \N__9061\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__9061\,
            I => \N__9057\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__9060\,
            I => \N__9054\
        );

    \I__1383\ : CascadeBuf
    port map (
            O => \N__9057\,
            I => \N__9051\
        );

    \I__1382\ : CascadeBuf
    port map (
            O => \N__9054\,
            I => \N__9048\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__9051\,
            I => \N__9045\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__9048\,
            I => \N__9042\
        );

    \I__1379\ : CascadeBuf
    port map (
            O => \N__9045\,
            I => \N__9039\
        );

    \I__1378\ : CascadeBuf
    port map (
            O => \N__9042\,
            I => \N__9036\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__9039\,
            I => \N__9033\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__9036\,
            I => \N__9030\
        );

    \I__1375\ : CascadeBuf
    port map (
            O => \N__9033\,
            I => \N__9027\
        );

    \I__1374\ : CascadeBuf
    port map (
            O => \N__9030\,
            I => \N__9024\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__9027\,
            I => \N__9021\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__9024\,
            I => \N__9018\
        );

    \I__1371\ : CascadeBuf
    port map (
            O => \N__9021\,
            I => \N__9015\
        );

    \I__1370\ : CascadeBuf
    port map (
            O => \N__9018\,
            I => \N__9012\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__9015\,
            I => \N__9009\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__9012\,
            I => \N__9006\
        );

    \I__1367\ : CascadeBuf
    port map (
            O => \N__9009\,
            I => \N__9003\
        );

    \I__1366\ : CascadeBuf
    port map (
            O => \N__9006\,
            I => \N__9000\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__9003\,
            I => \N__8997\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__9000\,
            I => \N__8994\
        );

    \I__1363\ : CascadeBuf
    port map (
            O => \N__8997\,
            I => \N__8991\
        );

    \I__1362\ : CascadeBuf
    port map (
            O => \N__8994\,
            I => \N__8988\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__8991\,
            I => \N__8985\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__8988\,
            I => \N__8982\
        );

    \I__1359\ : CascadeBuf
    port map (
            O => \N__8985\,
            I => \N__8979\
        );

    \I__1358\ : CascadeBuf
    port map (
            O => \N__8982\,
            I => \N__8976\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__8979\,
            I => \N__8973\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__8976\,
            I => \N__8970\
        );

    \I__1355\ : CascadeBuf
    port map (
            O => \N__8973\,
            I => \N__8967\
        );

    \I__1354\ : CascadeBuf
    port map (
            O => \N__8970\,
            I => \N__8964\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__8967\,
            I => \N__8961\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__8964\,
            I => \N__8958\
        );

    \I__1351\ : CascadeBuf
    port map (
            O => \N__8961\,
            I => \N__8955\
        );

    \I__1350\ : CascadeBuf
    port map (
            O => \N__8958\,
            I => \N__8952\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__8955\,
            I => \N__8949\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__8952\,
            I => \N__8946\
        );

    \I__1347\ : CascadeBuf
    port map (
            O => \N__8949\,
            I => \N__8943\
        );

    \I__1346\ : CascadeBuf
    port map (
            O => \N__8946\,
            I => \N__8940\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__8943\,
            I => \N__8937\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__8940\,
            I => \N__8934\
        );

    \I__1343\ : CascadeBuf
    port map (
            O => \N__8937\,
            I => \N__8931\
        );

    \I__1342\ : CascadeBuf
    port map (
            O => \N__8934\,
            I => \N__8928\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__8931\,
            I => \N__8925\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__8928\,
            I => \N__8922\
        );

    \I__1339\ : CascadeBuf
    port map (
            O => \N__8925\,
            I => \N__8919\
        );

    \I__1338\ : CascadeBuf
    port map (
            O => \N__8922\,
            I => \N__8916\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__8919\,
            I => \N__8913\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__8916\,
            I => \N__8910\
        );

    \I__1335\ : CascadeBuf
    port map (
            O => \N__8913\,
            I => \N__8907\
        );

    \I__1334\ : CascadeBuf
    port map (
            O => \N__8910\,
            I => \N__8904\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__8907\,
            I => \N__8901\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__8904\,
            I => \N__8898\
        );

    \I__1331\ : CascadeBuf
    port map (
            O => \N__8901\,
            I => \N__8895\
        );

    \I__1330\ : CascadeBuf
    port map (
            O => \N__8898\,
            I => \N__8892\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__8895\,
            I => \N__8889\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__8892\,
            I => \N__8886\
        );

    \I__1327\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8883\
        );

    \I__1326\ : CascadeBuf
    port map (
            O => \N__8886\,
            I => \N__8880\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__8883\,
            I => \N__8877\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__8880\,
            I => \N__8874\
        );

    \I__1323\ : Span4Mux_h
    port map (
            O => \N__8877\,
            I => \N__8871\
        );

    \I__1322\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8868\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__8871\,
            I => \N__8865\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__8868\,
            I => \N__8862\
        );

    \I__1319\ : Sp12to4
    port map (
            O => \N__8865\,
            I => \N__8859\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__8862\,
            I => \N__8856\
        );

    \I__1317\ : Span12Mux_s9_v
    port map (
            O => \N__8859\,
            I => \N__8851\
        );

    \I__1316\ : Span12Mux_s9_v
    port map (
            O => \N__8856\,
            I => \N__8851\
        );

    \I__1315\ : Odrv12
    port map (
            O => \N__8851\,
            I => n26
        );

    \I__1314\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8843\
        );

    \I__1313\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8840\
        );

    \I__1312\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8837\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__8843\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__8840\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__8837\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__1308\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8827\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__8827\,
            I => \receive_module.rx_counter.n10_adj_570\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__8824\,
            I => \N__8821\
        );

    \I__1305\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8816\
        );

    \I__1304\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8813\
        );

    \I__1303\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8810\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__8816\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__8813\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__8810\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__1299\ : IoInMux
    port map (
            O => \N__8803\,
            I => \N__8800\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__8800\,
            I => \N__8797\
        );

    \I__1297\ : IoSpan4Mux
    port map (
            O => \N__8797\,
            I => \N__8794\
        );

    \I__1296\ : Sp12to4
    port map (
            O => \N__8794\,
            I => \N__8791\
        );

    \I__1295\ : Span12Mux_s9_v
    port map (
            O => \N__8791\,
            I => \N__8787\
        );

    \I__1294\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8784\
        );

    \I__1293\ : Odrv12
    port map (
            O => \N__8787\,
            I => \LED_c\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__8784\,
            I => \LED_c\
        );

    \I__1291\ : InMux
    port map (
            O => \N__8779\,
            I => \transmit_module.n2743\
        );

    \I__1290\ : InMux
    port map (
            O => \N__8776\,
            I => \transmit_module.n2744\
        );

    \I__1289\ : InMux
    port map (
            O => \N__8773\,
            I => \transmit_module.n2745\
        );

    \I__1288\ : InMux
    port map (
            O => \N__8770\,
            I => \transmit_module.n2746\
        );

    \I__1287\ : InMux
    port map (
            O => \N__8767\,
            I => \bfn_15_18_0_\
        );

    \I__1286\ : InMux
    port map (
            O => \N__8764\,
            I => \transmit_module.n2748\
        );

    \I__1285\ : InMux
    port map (
            O => \N__8761\,
            I => \transmit_module.n2749\
        );

    \I__1284\ : InMux
    port map (
            O => \N__8758\,
            I => \transmit_module.n2750\
        );

    \I__1283\ : InMux
    port map (
            O => \N__8755\,
            I => \transmit_module.n2751\
        );

    \I__1282\ : InMux
    port map (
            O => \N__8752\,
            I => \N__8747\
        );

    \I__1281\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8744\
        );

    \I__1280\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8741\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8738\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__8744\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__8741\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__8738\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1275\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8728\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__8728\,
            I => \transmit_module.video_signal_controller.n3183\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__8725\,
            I => \N__8721\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__8724\,
            I => \N__8718\
        );

    \I__1271\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8714\
        );

    \I__1270\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8711\
        );

    \I__1269\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8708\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8705\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__8711\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__8708\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__8705\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1264\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8695\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__8695\,
            I => \transmit_module.video_signal_controller.n6\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__8692\,
            I => \N__8688\
        );

    \I__1261\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8683\
        );

    \I__1260\ : InMux
    port map (
            O => \N__8688\,
            I => \N__8680\
        );

    \I__1259\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8677\
        );

    \I__1258\ : InMux
    port map (
            O => \N__8686\,
            I => \N__8674\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__8683\,
            I => \N__8671\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__8680\,
            I => \N__8668\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__8677\,
            I => \N__8665\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__8674\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__8671\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__8668\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__8665\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1250\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8650\
        );

    \I__1249\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8647\
        );

    \I__1248\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8644\
        );

    \I__1247\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8641\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__8650\,
            I => \N__8636\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__8647\,
            I => \N__8636\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__8644\,
            I => \N__8633\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__8641\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__8636\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__8633\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__8626\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_558_cascade_\
        );

    \I__1239\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8620\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__8620\,
            I => \transmit_module.video_signal_controller.n18\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__8617\,
            I => \VGA_VISIBLE_cascade_\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__8614\,
            I => \N__8610\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8607\
        );

    \I__1234\ : InMux
    port map (
            O => \N__8610\,
            I => \N__8604\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__8607\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__8604\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__1231\ : InMux
    port map (
            O => \N__8599\,
            I => \transmit_module.n2740\
        );

    \I__1230\ : InMux
    port map (
            O => \N__8596\,
            I => \transmit_module.n2741\
        );

    \I__1229\ : InMux
    port map (
            O => \N__8593\,
            I => \transmit_module.n2742\
        );

    \I__1228\ : InMux
    port map (
            O => \N__8590\,
            I => \bfn_15_11_0_\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__8587\,
            I => \N__8583\
        );

    \I__1226\ : InMux
    port map (
            O => \N__8586\,
            I => \N__8580\
        );

    \I__1225\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8577\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__8580\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__8577\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__1222\ : InMux
    port map (
            O => \N__8572\,
            I => \receive_module.rx_counter.n2753\
        );

    \I__1221\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8565\
        );

    \I__1220\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8562\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__8565\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__8562\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__1217\ : InMux
    port map (
            O => \N__8557\,
            I => \receive_module.rx_counter.n2754\
        );

    \I__1216\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8550\
        );

    \I__1215\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8547\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__8550\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__8547\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__1212\ : InMux
    port map (
            O => \N__8542\,
            I => \receive_module.rx_counter.n2755\
        );

    \I__1211\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8535\
        );

    \I__1210\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8532\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__8535\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__8532\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__1207\ : InMux
    port map (
            O => \N__8527\,
            I => \receive_module.rx_counter.n2756\
        );

    \I__1206\ : InMux
    port map (
            O => \N__8524\,
            I => \receive_module.rx_counter.n2757\
        );

    \I__1205\ : SRMux
    port map (
            O => \N__8521\,
            I => \N__8518\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8515\
        );

    \I__1203\ : Span4Mux_h
    port map (
            O => \N__8515\,
            I => \N__8512\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__8512\,
            I => \receive_module.rx_counter.n2227\
        );

    \I__1201\ : IoInMux
    port map (
            O => \N__8509\,
            I => \N__8506\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8503\
        );

    \I__1199\ : IoSpan4Mux
    port map (
            O => \N__8503\,
            I => \N__8499\
        );

    \I__1198\ : IoInMux
    port map (
            O => \N__8502\,
            I => \N__8495\
        );

    \I__1197\ : Span4Mux_s2_v
    port map (
            O => \N__8499\,
            I => \N__8492\
        );

    \I__1196\ : IoInMux
    port map (
            O => \N__8498\,
            I => \N__8489\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__8495\,
            I => \N__8486\
        );

    \I__1194\ : Span4Mux_v
    port map (
            O => \N__8492\,
            I => \N__8483\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8480\
        );

    \I__1192\ : Span4Mux_s2_v
    port map (
            O => \N__8486\,
            I => \N__8477\
        );

    \I__1191\ : Sp12to4
    port map (
            O => \N__8483\,
            I => \N__8472\
        );

    \I__1190\ : Span12Mux_s2_h
    port map (
            O => \N__8480\,
            I => \N__8472\
        );

    \I__1189\ : Span4Mux_h
    port map (
            O => \N__8477\,
            I => \N__8469\
        );

    \I__1188\ : Span12Mux_v
    port map (
            O => \N__8472\,
            I => \N__8466\
        );

    \I__1187\ : Sp12to4
    port map (
            O => \N__8469\,
            I => \N__8463\
        );

    \I__1186\ : Span12Mux_h
    port map (
            O => \N__8466\,
            I => \N__8460\
        );

    \I__1185\ : Span12Mux_s9_v
    port map (
            O => \N__8463\,
            I => \N__8457\
        );

    \I__1184\ : Odrv12
    port map (
            O => \N__8460\,
            I => n1955
        );

    \I__1183\ : Odrv12
    port map (
            O => \N__8457\,
            I => n1955
        );

    \I__1182\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8449\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__8449\,
            I => \N__8446\
        );

    \I__1180\ : Span4Mux_h
    port map (
            O => \N__8446\,
            I => \N__8443\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__8443\,
            I => \TX_DATA_2\
        );

    \I__1178\ : IoInMux
    port map (
            O => \N__8440\,
            I => \N__8437\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__8437\,
            I => \N__8434\
        );

    \I__1176\ : IoSpan4Mux
    port map (
            O => \N__8434\,
            I => \N__8430\
        );

    \I__1175\ : IoInMux
    port map (
            O => \N__8433\,
            I => \N__8426\
        );

    \I__1174\ : IoSpan4Mux
    port map (
            O => \N__8430\,
            I => \N__8423\
        );

    \I__1173\ : IoInMux
    port map (
            O => \N__8429\,
            I => \N__8420\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__8426\,
            I => \N__8417\
        );

    \I__1171\ : Span4Mux_s3_v
    port map (
            O => \N__8423\,
            I => \N__8414\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8411\
        );

    \I__1169\ : Span12Mux_s5_v
    port map (
            O => \N__8417\,
            I => \N__8408\
        );

    \I__1168\ : Sp12to4
    port map (
            O => \N__8414\,
            I => \N__8405\
        );

    \I__1167\ : Span12Mux_s2_h
    port map (
            O => \N__8411\,
            I => \N__8402\
        );

    \I__1166\ : Span12Mux_v
    port map (
            O => \N__8408\,
            I => \N__8399\
        );

    \I__1165\ : Span12Mux_s10_v
    port map (
            O => \N__8405\,
            I => \N__8394\
        );

    \I__1164\ : Span12Mux_h
    port map (
            O => \N__8402\,
            I => \N__8394\
        );

    \I__1163\ : Odrv12
    port map (
            O => \N__8399\,
            I => n1953
        );

    \I__1162\ : Odrv12
    port map (
            O => \N__8394\,
            I => n1953
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__8389\,
            I => \line_buffer.n3031_cascade_\
        );

    \I__1160\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8383\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__8383\,
            I => \N__8380\
        );

    \I__1158\ : Odrv12
    port map (
            O => \N__8380\,
            I => \line_buffer.n3030\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__8377\,
            I => \line_buffer.n3095_cascade_\
        );

    \I__1156\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8371\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8368\
        );

    \I__1154\ : Span4Mux_h
    port map (
            O => \N__8368\,
            I => \N__8365\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__8365\,
            I => \line_buffer.n3040\
        );

    \I__1152\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8359\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8356\
        );

    \I__1150\ : Span4Mux_v
    port map (
            O => \N__8356\,
            I => \N__8353\
        );

    \I__1149\ : Span4Mux_h
    port map (
            O => \N__8353\,
            I => \N__8350\
        );

    \I__1148\ : Span4Mux_h
    port map (
            O => \N__8350\,
            I => \N__8347\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__8347\,
            I => \line_buffer.n625\
        );

    \I__1146\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8341\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__8341\,
            I => \N__8338\
        );

    \I__1144\ : Span4Mux_v
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__1143\ : Sp12to4
    port map (
            O => \N__8335\,
            I => \N__8332\
        );

    \I__1142\ : Span12Mux_h
    port map (
            O => \N__8332\,
            I => \N__8329\
        );

    \I__1141\ : Span12Mux_v
    port map (
            O => \N__8329\,
            I => \N__8326\
        );

    \I__1140\ : Odrv12
    port map (
            O => \N__8326\,
            I => \line_buffer.n617\
        );

    \I__1139\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8320\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__8320\,
            I => \N__8317\
        );

    \I__1137\ : Odrv12
    port map (
            O => \N__8317\,
            I => \line_buffer.n3089\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__8314\,
            I => \line_buffer.n3092_cascade_\
        );

    \I__1135\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8308\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__8308\,
            I => \line_buffer.n3146\
        );

    \I__1133\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8302\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__8302\,
            I => \N__8299\
        );

    \I__1131\ : Span12Mux_h
    port map (
            O => \N__8299\,
            I => \N__8296\
        );

    \I__1130\ : Odrv12
    port map (
            O => \N__8296\,
            I => \line_buffer.n626\
        );

    \I__1129\ : InMux
    port map (
            O => \N__8293\,
            I => \N__8290\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1127\ : Span4Mux_h
    port map (
            O => \N__8287\,
            I => \N__8284\
        );

    \I__1126\ : Span4Mux_h
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__1125\ : Sp12to4
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1124\ : Odrv12
    port map (
            O => \N__8278\,
            I => \line_buffer.n618\
        );

    \I__1123\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__8272\,
            I => \N__8269\
        );

    \I__1121\ : Odrv12
    port map (
            O => \N__8269\,
            I => \line_buffer.n3039\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__8266\,
            I => \receive_module.rx_counter.n10_adj_570_cascade_\
        );

    \I__1119\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8258\
        );

    \I__1118\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8255\
        );

    \I__1117\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8252\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__8258\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__8255\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__8252\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1113\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8240\
        );

    \I__1112\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8235\
        );

    \I__1111\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8235\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__8240\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__8235\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1108\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8227\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__8227\,
            I => \transmit_module.X_DELTA_PATTERN_1\
        );

    \I__1106\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8221\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__8221\,
            I => \transmit_module.X_DELTA_PATTERN_2\
        );

    \I__1104\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__8215\,
            I => \transmit_module.X_DELTA_PATTERN_6\
        );

    \I__1102\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__8209\,
            I => \transmit_module.X_DELTA_PATTERN_5\
        );

    \I__1100\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8203\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__8203\,
            I => \transmit_module.X_DELTA_PATTERN_4\
        );

    \I__1098\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__8197\,
            I => \transmit_module.X_DELTA_PATTERN_3\
        );

    \I__1096\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8191\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__8191\,
            I => \N__8188\
        );

    \I__1094\ : Odrv12
    port map (
            O => \N__8188\,
            I => \line_buffer.n755\
        );

    \I__1093\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8182\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__8182\,
            I => \N__8179\
        );

    \I__1091\ : Span12Mux_h
    port map (
            O => \N__8179\,
            I => \N__8176\
        );

    \I__1090\ : Span12Mux_v
    port map (
            O => \N__8176\,
            I => \N__8173\
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__8173\,
            I => \line_buffer.n747\
        );

    \I__1088\ : InMux
    port map (
            O => \N__8170\,
            I => \transmit_module.video_signal_controller.n2778\
        );

    \I__1087\ : InMux
    port map (
            O => \N__8167\,
            I => \transmit_module.video_signal_controller.n2779\
        );

    \I__1086\ : InMux
    port map (
            O => \N__8164\,
            I => \transmit_module.video_signal_controller.n2780\
        );

    \I__1085\ : InMux
    port map (
            O => \N__8161\,
            I => \transmit_module.video_signal_controller.n2781\
        );

    \I__1084\ : SRMux
    port map (
            O => \N__8158\,
            I => \N__8154\
        );

    \I__1083\ : SRMux
    port map (
            O => \N__8157\,
            I => \N__8150\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__8154\,
            I => \N__8147\
        );

    \I__1081\ : CEMux
    port map (
            O => \N__8153\,
            I => \N__8144\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__8150\,
            I => \N__8141\
        );

    \I__1079\ : Span4Mux_h
    port map (
            O => \N__8147\,
            I => \N__8138\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__8144\,
            I => n2147
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__8141\,
            I => n2147
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__8138\,
            I => n2147
        );

    \I__1075\ : SRMux
    port map (
            O => \N__8131\,
            I => \N__8128\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__8128\,
            I => \transmit_module.video_signal_controller.n2262\
        );

    \I__1073\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8121\
        );

    \I__1072\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8118\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__8121\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__8118\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__8113\,
            I => \transmit_module.video_signal_controller.n3022_cascade_\
        );

    \I__1068\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8105\
        );

    \I__1067\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8102\
        );

    \I__1066\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8098\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__8105\,
            I => \N__8093\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__8102\,
            I => \N__8093\
        );

    \I__1063\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8090\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__8098\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__8093\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__8090\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1059\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8076\
        );

    \I__1058\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8073\
        );

    \I__1057\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8068\
        );

    \I__1056\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8068\
        );

    \I__1055\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8065\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__8076\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__8073\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__8068\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__8065\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__1049\ : InMux
    port map (
            O => \N__8053\,
            I => \N__8046\
        );

    \I__1048\ : InMux
    port map (
            O => \N__8052\,
            I => \N__8043\
        );

    \I__1047\ : InMux
    port map (
            O => \N__8051\,
            I => \N__8036\
        );

    \I__1046\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8036\
        );

    \I__1045\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8036\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__8046\,
            I => \N__8033\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__8043\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__8036\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__8033\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1040\ : InMux
    port map (
            O => \N__8026\,
            I => \N__8019\
        );

    \I__1039\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8016\
        );

    \I__1038\ : InMux
    port map (
            O => \N__8024\,
            I => \N__8011\
        );

    \I__1037\ : InMux
    port map (
            O => \N__8023\,
            I => \N__8011\
        );

    \I__1036\ : InMux
    port map (
            O => \N__8022\,
            I => \N__8008\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__8019\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__8016\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__8011\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__8008\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1031\ : InMux
    port map (
            O => \N__7999\,
            I => \N__7994\
        );

    \I__1030\ : InMux
    port map (
            O => \N__7998\,
            I => \N__7989\
        );

    \I__1029\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7989\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__7994\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__7989\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1026\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7979\
        );

    \I__1025\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7976\
        );

    \I__1024\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7973\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__7979\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__7976\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__7973\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1020\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7963\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__7963\,
            I => \transmit_module.X_DELTA_PATTERN_15\
        );

    \I__1018\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7957\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__7957\,
            I => \transmit_module.X_DELTA_PATTERN_14\
        );

    \I__1016\ : InMux
    port map (
            O => \N__7954\,
            I => \N__7951\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__7951\,
            I => \N__7948\
        );

    \I__1014\ : Odrv12
    port map (
            O => \N__7948\,
            I => \line_buffer.n754\
        );

    \I__1013\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7942\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__7942\,
            I => \N__7939\
        );

    \I__1011\ : Span12Mux_h
    port map (
            O => \N__7939\,
            I => \N__7936\
        );

    \I__1010\ : Span12Mux_v
    port map (
            O => \N__7936\,
            I => \N__7933\
        );

    \I__1009\ : Odrv12
    port map (
            O => \N__7933\,
            I => \line_buffer.n746\
        );

    \I__1008\ : InMux
    port map (
            O => \N__7930\,
            I => \N__7927\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__7927\,
            I => \N__7924\
        );

    \I__1006\ : Span12Mux_v
    port map (
            O => \N__7924\,
            I => \N__7921\
        );

    \I__1005\ : Span12Mux_h
    port map (
            O => \N__7921\,
            I => \N__7918\
        );

    \I__1004\ : Odrv12
    port map (
            O => \N__7918\,
            I => \line_buffer.n682\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__7915\,
            I => \line_buffer.n3143_cascade_\
        );

    \I__1002\ : InMux
    port map (
            O => \N__7912\,
            I => \N__7909\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1000\ : Span4Mux_v
    port map (
            O => \N__7906\,
            I => \N__7903\
        );

    \I__999\ : Span4Mux_h
    port map (
            O => \N__7903\,
            I => \N__7900\
        );

    \I__998\ : Span4Mux_v
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__997\ : Span4Mux_v
    port map (
            O => \N__7897\,
            I => \N__7894\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__7894\,
            I => \line_buffer.n690\
        );

    \I__995\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7888\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__7888\,
            I => \N__7885\
        );

    \I__993\ : Span4Mux_h
    port map (
            O => \N__7885\,
            I => \N__7882\
        );

    \I__992\ : Span4Mux_h
    port map (
            O => \N__7882\,
            I => \N__7879\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__7879\,
            I => \line_buffer.n694\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__7876\,
            I => \N__7873\
        );

    \I__989\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7870\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7867\
        );

    \I__987\ : Span12Mux_v
    port map (
            O => \N__7867\,
            I => \N__7864\
        );

    \I__986\ : Span12Mux_v
    port map (
            O => \N__7864\,
            I => \N__7861\
        );

    \I__985\ : Span12Mux_h
    port map (
            O => \N__7861\,
            I => \N__7858\
        );

    \I__984\ : Odrv12
    port map (
            O => \N__7858\,
            I => \line_buffer.n686\
        );

    \I__983\ : InMux
    port map (
            O => \N__7855\,
            I => \N__7852\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__7852\,
            I => \line_buffer.n3101\
        );

    \I__981\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7846\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__7846\,
            I => \N__7843\
        );

    \I__979\ : Span4Mux_h
    port map (
            O => \N__7843\,
            I => \N__7840\
        );

    \I__978\ : Span4Mux_h
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__7837\,
            I => \N__7834\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__7834\,
            I => \line_buffer.n691\
        );

    \I__975\ : InMux
    port map (
            O => \N__7831\,
            I => \N__7828\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__7828\,
            I => \N__7825\
        );

    \I__973\ : Span12Mux_h
    port map (
            O => \N__7825\,
            I => \N__7822\
        );

    \I__972\ : Odrv12
    port map (
            O => \N__7822\,
            I => \line_buffer.n683\
        );

    \I__971\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7816\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__7816\,
            I => \N__7813\
        );

    \I__969\ : Span4Mux_h
    port map (
            O => \N__7813\,
            I => \N__7810\
        );

    \I__968\ : Span4Mux_h
    port map (
            O => \N__7810\,
            I => \N__7807\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__7807\,
            I => \line_buffer.n722\
        );

    \I__966\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7801\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__7801\,
            I => \N__7798\
        );

    \I__964\ : Span4Mux_v
    port map (
            O => \N__7798\,
            I => \N__7795\
        );

    \I__963\ : Span4Mux_h
    port map (
            O => \N__7795\,
            I => \N__7792\
        );

    \I__962\ : Span4Mux_h
    port map (
            O => \N__7792\,
            I => \N__7789\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__7789\,
            I => \line_buffer.n714\
        );

    \I__960\ : InMux
    port map (
            O => \N__7786\,
            I => \bfn_14_14_0_\
        );

    \I__959\ : InMux
    port map (
            O => \N__7783\,
            I => \transmit_module.video_signal_controller.n2776\
        );

    \I__958\ : InMux
    port map (
            O => \N__7780\,
            I => \transmit_module.video_signal_controller.n2777\
        );

    \I__957\ : InMux
    port map (
            O => \N__7777\,
            I => \bfn_13_16_0_\
        );

    \I__956\ : InMux
    port map (
            O => \N__7774\,
            I => \transmit_module.video_signal_controller.n2774\
        );

    \I__955\ : InMux
    port map (
            O => \N__7771\,
            I => \transmit_module.video_signal_controller.n2775\
        );

    \I__954\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7765\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__7765\,
            I => \transmit_module.X_DELTA_PATTERN_13\
        );

    \I__952\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7759\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__7759\,
            I => \transmit_module.X_DELTA_PATTERN_10\
        );

    \I__950\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7753\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__7753\,
            I => \transmit_module.X_DELTA_PATTERN_12\
        );

    \I__948\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7747\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__7747\,
            I => \transmit_module.X_DELTA_PATTERN_11\
        );

    \I__946\ : InMux
    port map (
            O => \N__7744\,
            I => \N__7741\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__7741\,
            I => \transmit_module.X_DELTA_PATTERN_7\
        );

    \I__944\ : InMux
    port map (
            O => \N__7738\,
            I => \N__7734\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__7737\,
            I => \N__7729\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__7734\,
            I => \N__7726\
        );

    \I__941\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7723\
        );

    \I__940\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7720\
        );

    \I__939\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7717\
        );

    \I__938\ : Odrv4
    port map (
            O => \N__7726\,
            I => \Y_0\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__7723\,
            I => \Y_0\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__7720\,
            I => \Y_0\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__7717\,
            I => \Y_0\
        );

    \I__934\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7705\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__7705\,
            I => \N__7699\
        );

    \I__932\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7696\
        );

    \I__931\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7693\
        );

    \I__930\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7690\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__7699\,
            I => \Y_1\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__7696\,
            I => \Y_1\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__7693\,
            I => \Y_1\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__7690\,
            I => \Y_1\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__7681\,
            I => \n5_cascade_\
        );

    \I__924\ : InMux
    port map (
            O => \N__7678\,
            I => \N__7675\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__7675\,
            I => n3009
        );

    \I__922\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7668\
        );

    \I__921\ : InMux
    port map (
            O => \N__7671\,
            I => \N__7665\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__7668\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__7665\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__918\ : InMux
    port map (
            O => \N__7660\,
            I => \bfn_13_15_0_\
        );

    \I__917\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7653\
        );

    \I__916\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7650\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__7653\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__7650\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__913\ : InMux
    port map (
            O => \N__7645\,
            I => \transmit_module.video_signal_controller.n2766\
        );

    \I__912\ : InMux
    port map (
            O => \N__7642\,
            I => \N__7638\
        );

    \I__911\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7635\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__7638\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__7635\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__908\ : InMux
    port map (
            O => \N__7630\,
            I => \transmit_module.video_signal_controller.n2767\
        );

    \I__907\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7622\
        );

    \I__906\ : InMux
    port map (
            O => \N__7626\,
            I => \N__7619\
        );

    \I__905\ : InMux
    port map (
            O => \N__7625\,
            I => \N__7616\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__7622\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__7619\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__7616\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__901\ : InMux
    port map (
            O => \N__7609\,
            I => \transmit_module.video_signal_controller.n2768\
        );

    \I__900\ : InMux
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__899\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7593\
        );

    \I__898\ : InMux
    port map (
            O => \N__7604\,
            I => \N__7593\
        );

    \I__897\ : InMux
    port map (
            O => \N__7603\,
            I => \N__7593\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__7600\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__7593\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__894\ : InMux
    port map (
            O => \N__7588\,
            I => \transmit_module.video_signal_controller.n2769\
        );

    \I__893\ : InMux
    port map (
            O => \N__7585\,
            I => \transmit_module.video_signal_controller.n2770\
        );

    \I__892\ : InMux
    port map (
            O => \N__7582\,
            I => \transmit_module.video_signal_controller.n2771\
        );

    \I__891\ : InMux
    port map (
            O => \N__7579\,
            I => \transmit_module.video_signal_controller.n2772\
        );

    \I__890\ : InMux
    port map (
            O => \N__7576\,
            I => \N__7573\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__7573\,
            I => \transmit_module.X_DELTA_PATTERN_9\
        );

    \I__888\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7567\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__7567\,
            I => \transmit_module.X_DELTA_PATTERN_8\
        );

    \I__886\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7561\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__7561\,
            I => \N__7558\
        );

    \I__884\ : Span12Mux_v
    port map (
            O => \N__7558\,
            I => \N__7555\
        );

    \I__883\ : Odrv12
    port map (
            O => \N__7555\,
            I => \line_buffer.n758\
        );

    \I__882\ : InMux
    port map (
            O => \N__7552\,
            I => \N__7549\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__7549\,
            I => \N__7546\
        );

    \I__880\ : Span4Mux_v
    port map (
            O => \N__7546\,
            I => \N__7543\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__7543\,
            I => \line_buffer.n750\
        );

    \I__878\ : CEMux
    port map (
            O => \N__7540\,
            I => \N__7536\
        );

    \I__877\ : CEMux
    port map (
            O => \N__7539\,
            I => \N__7533\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__7536\,
            I => \receive_module.n2152\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__7533\,
            I => \receive_module.n2152\
        );

    \I__874\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7525\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__7525\,
            I => \N__7520\
        );

    \I__872\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7515\
        );

    \I__871\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7515\
        );

    \I__870\ : Span4Mux_v
    port map (
            O => \N__7520\,
            I => \N__7512\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__7515\,
            I => \N__7509\
        );

    \I__868\ : Span4Mux_h
    port map (
            O => \N__7512\,
            I => \N__7506\
        );

    \I__867\ : Span4Mux_v
    port map (
            O => \N__7509\,
            I => \N__7503\
        );

    \I__866\ : Span4Mux_h
    port map (
            O => \N__7506\,
            I => \N__7500\
        );

    \I__865\ : Sp12to4
    port map (
            O => \N__7503\,
            I => \N__7497\
        );

    \I__864\ : Sp12to4
    port map (
            O => \N__7500\,
            I => \N__7492\
        );

    \I__863\ : Span12Mux_h
    port map (
            O => \N__7497\,
            I => \N__7492\
        );

    \I__862\ : Odrv12
    port map (
            O => \N__7492\,
            I => \TVP_HSYNC_c\
        );

    \I__861\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7486\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__7486\,
            I => \receive_module.old_HS\
        );

    \I__859\ : InMux
    port map (
            O => \N__7483\,
            I => \N__7480\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__7480\,
            I => \transmit_module.video_signal_controller.n2484\
        );

    \I__857\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7471\
        );

    \I__856\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7468\
        );

    \I__855\ : InMux
    port map (
            O => \N__7475\,
            I => \N__7463\
        );

    \I__854\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7463\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__7471\,
            I => \N__7460\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__7468\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__7463\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__7460\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__7453\,
            I => \n2147_cascade_\
        );

    \I__848\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7444\
        );

    \I__847\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7441\
        );

    \I__846\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7436\
        );

    \I__845\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7436\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__7444\,
            I => \N__7433\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__7441\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__7436\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__7433\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__840\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7420\
        );

    \I__839\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7417\
        );

    \I__838\ : InMux
    port map (
            O => \N__7424\,
            I => \N__7412\
        );

    \I__837\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7412\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__7420\,
            I => \N__7409\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__7417\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__7412\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__7409\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__832\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7396\
        );

    \I__831\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7393\
        );

    \I__830\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7390\
        );

    \I__829\ : InMux
    port map (
            O => \N__7399\,
            I => \N__7387\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__7396\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__7393\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__7390\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__7387\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__7378\,
            I => \receive_module.rx_counter.n6_cascade_\
        );

    \I__823\ : InMux
    port map (
            O => \N__7375\,
            I => \N__7369\
        );

    \I__822\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7366\
        );

    \I__821\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7361\
        );

    \I__820\ : InMux
    port map (
            O => \N__7372\,
            I => \N__7361\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__7369\,
            I => \N__7358\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__7366\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__7361\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__7358\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__815\ : InMux
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__7348\,
            I => \N__7345\
        );

    \I__813\ : Span12Mux_v
    port map (
            O => \N__7345\,
            I => \N__7342\
        );

    \I__812\ : Odrv12
    port map (
            O => \N__7342\,
            I => \line_buffer.n723\
        );

    \I__811\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7336\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__809\ : Span12Mux_h
    port map (
            O => \N__7333\,
            I => \N__7330\
        );

    \I__808\ : Odrv12
    port map (
            O => \N__7330\,
            I => \line_buffer.n715\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__7327\,
            I => \N__7324\
        );

    \I__806\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7321\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__7321\,
            I => \transmit_module.video_signal_controller.n2972\
        );

    \I__804\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7315\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__7315\,
            I => \transmit_module.video_signal_controller.n3014\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__7312\,
            I => \transmit_module.video_signal_controller.n3186_cascade_\
        );

    \I__801\ : IoInMux
    port map (
            O => \N__7309\,
            I => \N__7306\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__7306\,
            I => \N__7303\
        );

    \I__799\ : Span4Mux_s3_h
    port map (
            O => \N__7303\,
            I => \N__7300\
        );

    \I__798\ : Sp12to4
    port map (
            O => \N__7300\,
            I => \N__7297\
        );

    \I__797\ : Span12Mux_v
    port map (
            O => \N__7297\,
            I => \N__7294\
        );

    \I__796\ : Odrv12
    port map (
            O => \N__7294\,
            I => \ADV_HSYNC_c\
        );

    \I__795\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7288\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__7288\,
            I => \transmit_module.video_signal_controller.n12\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__7285\,
            I => \transmit_module.video_signal_controller.n3182_cascade_\
        );

    \I__792\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7279\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__7279\,
            I => \transmit_module.video_signal_controller.n8\
        );

    \I__790\ : InMux
    port map (
            O => \N__7276\,
            I => \receive_module.rx_counter.n2759\
        );

    \I__789\ : InMux
    port map (
            O => \N__7273\,
            I => \receive_module.rx_counter.n2760\
        );

    \I__788\ : InMux
    port map (
            O => \N__7270\,
            I => \receive_module.rx_counter.n2761\
        );

    \I__787\ : InMux
    port map (
            O => \N__7267\,
            I => \receive_module.rx_counter.n2762\
        );

    \I__786\ : InMux
    port map (
            O => \N__7264\,
            I => \receive_module.rx_counter.n2763\
        );

    \I__785\ : InMux
    port map (
            O => \N__7261\,
            I => \receive_module.rx_counter.n2764\
        );

    \I__784\ : InMux
    port map (
            O => \N__7258\,
            I => \bfn_12_13_0_\
        );

    \I__783\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7252\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__7252\,
            I => \N__7246\
        );

    \I__781\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7243\
        );

    \I__780\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7238\
        );

    \I__779\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7238\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__7246\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__7243\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__7238\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__775\ : InMux
    port map (
            O => \N__7231\,
            I => \N__7225\
        );

    \I__774\ : InMux
    port map (
            O => \N__7230\,
            I => \N__7222\
        );

    \I__773\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7217\
        );

    \I__772\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7217\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__7225\,
            I => \N__7214\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__7222\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__7217\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__7214\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__7207\,
            I => \receive_module.rx_counter.n4_cascade_\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__7204\,
            I => \receive_module.rx_counter.n2986_cascade_\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__7201\,
            I => \receive_module.rx_counter.n2989_cascade_\
        );

    \I__764\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7195\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__7195\,
            I => \receive_module.rx_counter.n31_adj_572\
        );

    \I__762\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7189\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__7189\,
            I => \receive_module.rx_counter.n7\
        );

    \I__760\ : InMux
    port map (
            O => \N__7186\,
            I => \N__7183\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__7183\,
            I => \receive_module.rx_counter.n3166\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__7180\,
            I => \receive_module.rx_counter.n2978_cascade_\
        );

    \I__757\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7174\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__7174\,
            I => \receive_module.rx_counter.n4_adj_571\
        );

    \I__755\ : InMux
    port map (
            O => \N__7171\,
            I => \bfn_12_12_0_\
        );

    \I__754\ : InMux
    port map (
            O => \N__7168\,
            I => \receive_module.rx_counter.n2758\
        );

    \I__753\ : InMux
    port map (
            O => \N__7165\,
            I => \N__7161\
        );

    \I__752\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7158\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__7161\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__7158\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__749\ : InMux
    port map (
            O => \N__7153\,
            I => \receive_module.rx_counter.n2784\
        );

    \I__748\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7146\
        );

    \I__747\ : InMux
    port map (
            O => \N__7149\,
            I => \N__7143\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__7146\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__7143\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__744\ : InMux
    port map (
            O => \N__7138\,
            I => \receive_module.rx_counter.n2785\
        );

    \I__743\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7131\
        );

    \I__742\ : InMux
    port map (
            O => \N__7134\,
            I => \N__7128\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__7131\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__7128\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__739\ : InMux
    port map (
            O => \N__7123\,
            I => \receive_module.rx_counter.n2786\
        );

    \I__738\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7115\
        );

    \I__737\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7110\
        );

    \I__736\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7110\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__7115\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__7110\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__733\ : InMux
    port map (
            O => \N__7105\,
            I => \receive_module.rx_counter.n2787\
        );

    \I__732\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7095\
        );

    \I__731\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7095\
        );

    \I__730\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7092\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__7095\,
            I => \N__7089\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__7092\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__727\ : Odrv4
    port map (
            O => \N__7089\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__726\ : InMux
    port map (
            O => \N__7084\,
            I => \receive_module.rx_counter.n2788\
        );

    \I__725\ : InMux
    port map (
            O => \N__7081\,
            I => \N__7077\
        );

    \I__724\ : InMux
    port map (
            O => \N__7080\,
            I => \N__7074\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__7077\,
            I => \N__7071\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__7074\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__7071\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__720\ : InMux
    port map (
            O => \N__7066\,
            I => \bfn_10_15_0_\
        );

    \I__719\ : InMux
    port map (
            O => \N__7063\,
            I => \receive_module.rx_counter.n2790\
        );

    \I__718\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7056\
        );

    \I__717\ : InMux
    port map (
            O => \N__7059\,
            I => \N__7053\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7050\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__7053\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__7050\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__713\ : SRMux
    port map (
            O => \N__7045\,
            I => \N__7041\
        );

    \I__712\ : SRMux
    port map (
            O => \N__7044\,
            I => \N__7038\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__7041\,
            I => \N__7035\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__7038\,
            I => \N__7032\
        );

    \I__709\ : Sp12to4
    port map (
            O => \N__7035\,
            I => \N__7029\
        );

    \I__708\ : Span4Mux_v
    port map (
            O => \N__7032\,
            I => \N__7026\
        );

    \I__707\ : Odrv12
    port map (
            O => \N__7029\,
            I => n3184
        );

    \I__706\ : Odrv4
    port map (
            O => \N__7026\,
            I => n3184
        );

    \I__705\ : InMux
    port map (
            O => \N__7021\,
            I => \N__7018\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__7018\,
            I => \N__7015\
        );

    \I__703\ : Span4Mux_v
    port map (
            O => \N__7015\,
            I => \N__7012\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__7012\,
            I => \line_buffer.n759\
        );

    \I__701\ : InMux
    port map (
            O => \N__7009\,
            I => \N__7006\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__7006\,
            I => \N__7003\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__7003\,
            I => \N__7000\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__7000\,
            I => \line_buffer.n751\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__6997\,
            I => \receive_module.rx_counter.n2975_cascade_\
        );

    \I__696\ : SRMux
    port map (
            O => \N__6994\,
            I => \N__6989\
        );

    \I__695\ : SRMux
    port map (
            O => \N__6993\,
            I => \N__6986\
        );

    \I__694\ : SRMux
    port map (
            O => \N__6992\,
            I => \N__6982\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__6989\,
            I => \N__6977\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__6986\,
            I => \N__6977\
        );

    \I__691\ : SRMux
    port map (
            O => \N__6985\,
            I => \N__6974\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__6982\,
            I => \N__6971\
        );

    \I__689\ : Span4Mux_v
    port map (
            O => \N__6977\,
            I => \N__6966\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__6974\,
            I => \N__6966\
        );

    \I__687\ : Span4Mux_v
    port map (
            O => \N__6971\,
            I => \N__6963\
        );

    \I__686\ : Span4Mux_v
    port map (
            O => \N__6966\,
            I => \N__6960\
        );

    \I__685\ : Span4Mux_v
    port map (
            O => \N__6963\,
            I => \N__6957\
        );

    \I__684\ : Span4Mux_v
    port map (
            O => \N__6960\,
            I => \N__6952\
        );

    \I__683\ : Span4Mux_v
    port map (
            O => \N__6957\,
            I => \N__6952\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__6952\,
            I => \line_buffer.n698\
        );

    \I__681\ : InMux
    port map (
            O => \N__6949\,
            I => \N__6946\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__6946\,
            I => \receive_module.rx_counter.n2900\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__6943\,
            I => \receive_module.rx_counter.n2900_cascade_\
        );

    \I__678\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6937\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__6937\,
            I => \receive_module.rx_counter.n2943\
        );

    \I__676\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6931\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__6931\,
            I => \receive_module.rx_counter.n10\
        );

    \I__674\ : InMux
    port map (
            O => \N__6928\,
            I => \bfn_10_14_0_\
        );

    \I__673\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6922\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__6922\,
            I => \receive_module.rx_counter.n9\
        );

    \I__671\ : InMux
    port map (
            O => \N__6919\,
            I => \receive_module.rx_counter.n2782\
        );

    \I__670\ : InMux
    port map (
            O => \N__6916\,
            I => \N__6913\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__6913\,
            I => \receive_module.rx_counter.n8\
        );

    \I__668\ : InMux
    port map (
            O => \N__6910\,
            I => \receive_module.rx_counter.n2783\
        );

    \I__667\ : InMux
    port map (
            O => \N__6907\,
            I => \N__6904\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__6904\,
            I => \N__6901\
        );

    \I__665\ : Span4Mux_s2_v
    port map (
            O => \N__6901\,
            I => \N__6897\
        );

    \I__664\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6894\
        );

    \I__663\ : Span4Mux_v
    port map (
            O => \N__6897\,
            I => \N__6889\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__6894\,
            I => \N__6889\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__6889\,
            I => \N__6885\
        );

    \I__660\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6882\
        );

    \I__659\ : Span4Mux_v
    port map (
            O => \N__6885\,
            I => \N__6876\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__6882\,
            I => \N__6876\
        );

    \I__657\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6873\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__6876\,
            I => \N__6868\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__6873\,
            I => \N__6868\
        );

    \I__654\ : Span4Mux_v
    port map (
            O => \N__6868\,
            I => \N__6863\
        );

    \I__653\ : InMux
    port map (
            O => \N__6867\,
            I => \N__6860\
        );

    \I__652\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6857\
        );

    \I__651\ : Span4Mux_v
    port map (
            O => \N__6863\,
            I => \N__6852\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__6860\,
            I => \N__6852\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__6857\,
            I => \N__6849\
        );

    \I__648\ : Span4Mux_h
    port map (
            O => \N__6852\,
            I => \N__6845\
        );

    \I__647\ : Span4Mux_h
    port map (
            O => \N__6849\,
            I => \N__6842\
        );

    \I__646\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6839\
        );

    \I__645\ : Span4Mux_h
    port map (
            O => \N__6845\,
            I => \N__6836\
        );

    \I__644\ : Span4Mux_v
    port map (
            O => \N__6842\,
            I => \N__6832\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__6839\,
            I => \N__6829\
        );

    \I__642\ : Span4Mux_h
    port map (
            O => \N__6836\,
            I => \N__6826\
        );

    \I__641\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6823\
        );

    \I__640\ : Span4Mux_v
    port map (
            O => \N__6832\,
            I => \N__6818\
        );

    \I__639\ : Span4Mux_h
    port map (
            O => \N__6829\,
            I => \N__6818\
        );

    \I__638\ : Span4Mux_h
    port map (
            O => \N__6826\,
            I => \N__6813\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__6823\,
            I => \N__6813\
        );

    \I__636\ : Span4Mux_v
    port map (
            O => \N__6818\,
            I => \N__6810\
        );

    \I__635\ : Span4Mux_h
    port map (
            O => \N__6813\,
            I => \N__6807\
        );

    \I__634\ : Span4Mux_v
    port map (
            O => \N__6810\,
            I => \N__6804\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__6807\,
            I => \N__6801\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__6804\,
            I => \TVP_VIDEO_c_2\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__6801\,
            I => \TVP_VIDEO_c_2\
        );

    \I__630\ : SRMux
    port map (
            O => \N__6796\,
            I => \N__6792\
        );

    \I__629\ : SRMux
    port map (
            O => \N__6795\,
            I => \N__6789\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__6792\,
            I => \N__6785\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__6789\,
            I => \N__6782\
        );

    \I__626\ : SRMux
    port map (
            O => \N__6788\,
            I => \N__6779\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__6785\,
            I => \N__6776\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__6782\,
            I => \N__6771\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6771\
        );

    \I__622\ : Span4Mux_v
    port map (
            O => \N__6776\,
            I => \N__6768\
        );

    \I__621\ : Span4Mux_v
    port map (
            O => \N__6771\,
            I => \N__6765\
        );

    \I__620\ : Span4Mux_v
    port map (
            O => \N__6768\,
            I => \N__6759\
        );

    \I__619\ : Span4Mux_h
    port map (
            O => \N__6765\,
            I => \N__6759\
        );

    \I__618\ : SRMux
    port map (
            O => \N__6764\,
            I => \N__6756\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__6759\,
            I => \line_buffer.n730\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__6756\,
            I => \line_buffer.n730\
        );

    \I__615\ : SRMux
    port map (
            O => \N__6751\,
            I => \N__6748\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__6748\,
            I => \N__6743\
        );

    \I__613\ : SRMux
    port map (
            O => \N__6747\,
            I => \N__6740\
        );

    \I__612\ : SRMux
    port map (
            O => \N__6746\,
            I => \N__6737\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__6743\,
            I => \N__6733\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__6740\,
            I => \N__6728\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__6737\,
            I => \N__6728\
        );

    \I__608\ : SRMux
    port map (
            O => \N__6736\,
            I => \N__6725\
        );

    \I__607\ : Span4Mux_h
    port map (
            O => \N__6733\,
            I => \N__6722\
        );

    \I__606\ : Span4Mux_v
    port map (
            O => \N__6728\,
            I => \N__6717\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__6725\,
            I => \N__6717\
        );

    \I__604\ : Sp12to4
    port map (
            O => \N__6722\,
            I => \N__6714\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__6717\,
            I => \N__6711\
        );

    \I__602\ : Span12Mux_h
    port map (
            O => \N__6714\,
            I => \N__6708\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__6711\,
            I => \N__6705\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__6708\,
            I => \line_buffer.n632\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__6705\,
            I => \line_buffer.n632\
        );

    \I__598\ : SRMux
    port map (
            O => \N__6700\,
            I => \N__6697\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__6697\,
            I => \N__6693\
        );

    \I__596\ : SRMux
    port map (
            O => \N__6696\,
            I => \N__6688\
        );

    \I__595\ : Span4Mux_v
    port map (
            O => \N__6693\,
            I => \N__6685\
        );

    \I__594\ : SRMux
    port map (
            O => \N__6692\,
            I => \N__6682\
        );

    \I__593\ : SRMux
    port map (
            O => \N__6691\,
            I => \N__6679\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__6688\,
            I => \N__6676\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__6685\,
            I => \N__6671\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__6682\,
            I => \N__6671\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__6679\,
            I => \N__6668\
        );

    \I__588\ : Span4Mux_v
    port map (
            O => \N__6676\,
            I => \N__6663\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__6671\,
            I => \N__6663\
        );

    \I__586\ : Span4Mux_h
    port map (
            O => \N__6668\,
            I => \N__6660\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__6663\,
            I => \line_buffer.n762\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__6660\,
            I => \line_buffer.n762\
        );

    \I__583\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6651\
        );

    \I__582\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6648\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__6651\,
            I => \N__6641\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__6648\,
            I => \N__6641\
        );

    \I__579\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6638\
        );

    \I__578\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6635\
        );

    \I__577\ : Span4Mux_v
    port map (
            O => \N__6641\,
            I => \N__6627\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__6638\,
            I => \N__6627\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__6635\,
            I => \N__6627\
        );

    \I__574\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6623\
        );

    \I__573\ : Span4Mux_v
    port map (
            O => \N__6627\,
            I => \N__6620\
        );

    \I__572\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6617\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__6623\,
            I => \N__6614\
        );

    \I__570\ : Span4Mux_v
    port map (
            O => \N__6620\,
            I => \N__6609\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__6617\,
            I => \N__6609\
        );

    \I__568\ : Span4Mux_v
    port map (
            O => \N__6614\,
            I => \N__6604\
        );

    \I__567\ : Span4Mux_v
    port map (
            O => \N__6609\,
            I => \N__6601\
        );

    \I__566\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6598\
        );

    \I__565\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6595\
        );

    \I__564\ : Sp12to4
    port map (
            O => \N__6604\,
            I => \N__6592\
        );

    \I__563\ : Span4Mux_h
    port map (
            O => \N__6601\,
            I => \N__6589\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__6598\,
            I => \N__6586\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__6595\,
            I => \N__6583\
        );

    \I__560\ : Span12Mux_h
    port map (
            O => \N__6592\,
            I => \N__6580\
        );

    \I__559\ : Span4Mux_h
    port map (
            O => \N__6589\,
            I => \N__6577\
        );

    \I__558\ : Span4Mux_h
    port map (
            O => \N__6586\,
            I => \N__6574\
        );

    \I__557\ : Span4Mux_h
    port map (
            O => \N__6583\,
            I => \N__6571\
        );

    \I__556\ : Span12Mux_v
    port map (
            O => \N__6580\,
            I => \N__6566\
        );

    \I__555\ : Sp12to4
    port map (
            O => \N__6577\,
            I => \N__6566\
        );

    \I__554\ : IoSpan4Mux
    port map (
            O => \N__6574\,
            I => \N__6563\
        );

    \I__553\ : Span4Mux_h
    port map (
            O => \N__6571\,
            I => \N__6560\
        );

    \I__552\ : Span12Mux_v
    port map (
            O => \N__6566\,
            I => \N__6557\
        );

    \I__551\ : IoSpan4Mux
    port map (
            O => \N__6563\,
            I => \N__6554\
        );

    \I__550\ : Span4Mux_h
    port map (
            O => \N__6560\,
            I => \N__6551\
        );

    \I__549\ : Odrv12
    port map (
            O => \N__6557\,
            I => \TVP_VIDEO_c_8\
        );

    \I__548\ : Odrv4
    port map (
            O => \N__6554\,
            I => \TVP_VIDEO_c_8\
        );

    \I__547\ : Odrv4
    port map (
            O => \N__6551\,
            I => \TVP_VIDEO_c_8\
        );

    \I__546\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6540\
        );

    \I__545\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6537\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__6540\,
            I => \N__6531\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__6537\,
            I => \N__6531\
        );

    \I__542\ : InMux
    port map (
            O => \N__6536\,
            I => \N__6528\
        );

    \I__541\ : Span4Mux_v
    port map (
            O => \N__6531\,
            I => \N__6523\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__6528\,
            I => \N__6523\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__6523\,
            I => \N__6518\
        );

    \I__538\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6515\
        );

    \I__537\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6511\
        );

    \I__536\ : Span4Mux_v
    port map (
            O => \N__6518\,
            I => \N__6506\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__6515\,
            I => \N__6506\
        );

    \I__534\ : InMux
    port map (
            O => \N__6514\,
            I => \N__6503\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__6511\,
            I => \N__6500\
        );

    \I__532\ : Span4Mux_h
    port map (
            O => \N__6506\,
            I => \N__6497\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__6503\,
            I => \N__6494\
        );

    \I__530\ : Span12Mux_s11_h
    port map (
            O => \N__6500\,
            I => \N__6490\
        );

    \I__529\ : Sp12to4
    port map (
            O => \N__6497\,
            I => \N__6487\
        );

    \I__528\ : Span12Mux_s8_h
    port map (
            O => \N__6494\,
            I => \N__6484\
        );

    \I__527\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6481\
        );

    \I__526\ : Span12Mux_h
    port map (
            O => \N__6490\,
            I => \N__6478\
        );

    \I__525\ : Span12Mux_v
    port map (
            O => \N__6487\,
            I => \N__6475\
        );

    \I__524\ : Span12Mux_v
    port map (
            O => \N__6484\,
            I => \N__6472\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__6481\,
            I => \N__6469\
        );

    \I__522\ : Span12Mux_v
    port map (
            O => \N__6478\,
            I => \N__6465\
        );

    \I__521\ : Span12Mux_h
    port map (
            O => \N__6475\,
            I => \N__6462\
        );

    \I__520\ : Span12Mux_v
    port map (
            O => \N__6472\,
            I => \N__6459\
        );

    \I__519\ : Span4Mux_h
    port map (
            O => \N__6469\,
            I => \N__6456\
        );

    \I__518\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6453\
        );

    \I__517\ : Odrv12
    port map (
            O => \N__6465\,
            I => \TVP_VIDEO_c_9\
        );

    \I__516\ : Odrv12
    port map (
            O => \N__6462\,
            I => \TVP_VIDEO_c_9\
        );

    \I__515\ : Odrv12
    port map (
            O => \N__6459\,
            I => \TVP_VIDEO_c_9\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__6456\,
            I => \TVP_VIDEO_c_9\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__6453\,
            I => \TVP_VIDEO_c_9\
        );

    \I__512\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6437\
        );

    \I__511\ : InMux
    port map (
            O => \N__6441\,
            I => \N__6433\
        );

    \I__510\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6429\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__6437\,
            I => \N__6426\
        );

    \I__508\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6423\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6420\
        );

    \I__506\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6417\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__6429\,
            I => \N__6414\
        );

    \I__504\ : Span4Mux_h
    port map (
            O => \N__6426\,
            I => \N__6411\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__6423\,
            I => \N__6408\
        );

    \I__502\ : Span4Mux_v
    port map (
            O => \N__6420\,
            I => \N__6403\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__6417\,
            I => \N__6403\
        );

    \I__500\ : Span4Mux_v
    port map (
            O => \N__6414\,
            I => \N__6399\
        );

    \I__499\ : Span4Mux_h
    port map (
            O => \N__6411\,
            I => \N__6396\
        );

    \I__498\ : Span4Mux_h
    port map (
            O => \N__6408\,
            I => \N__6393\
        );

    \I__497\ : Span4Mux_v
    port map (
            O => \N__6403\,
            I => \N__6390\
        );

    \I__496\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6385\
        );

    \I__495\ : Sp12to4
    port map (
            O => \N__6399\,
            I => \N__6382\
        );

    \I__494\ : Sp12to4
    port map (
            O => \N__6396\,
            I => \N__6379\
        );

    \I__493\ : Span4Mux_h
    port map (
            O => \N__6393\,
            I => \N__6376\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__6390\,
            I => \N__6373\
        );

    \I__491\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6370\
        );

    \I__490\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6367\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__6385\,
            I => \N__6364\
        );

    \I__488\ : Span12Mux_h
    port map (
            O => \N__6382\,
            I => \N__6359\
        );

    \I__487\ : Span12Mux_s9_v
    port map (
            O => \N__6379\,
            I => \N__6359\
        );

    \I__486\ : Sp12to4
    port map (
            O => \N__6376\,
            I => \N__6356\
        );

    \I__485\ : Sp12to4
    port map (
            O => \N__6373\,
            I => \N__6351\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__6370\,
            I => \N__6351\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__6367\,
            I => \N__6348\
        );

    \I__482\ : Span4Mux_h
    port map (
            O => \N__6364\,
            I => \N__6345\
        );

    \I__481\ : Span12Mux_v
    port map (
            O => \N__6359\,
            I => \N__6342\
        );

    \I__480\ : Span12Mux_v
    port map (
            O => \N__6356\,
            I => \N__6335\
        );

    \I__479\ : Span12Mux_h
    port map (
            O => \N__6351\,
            I => \N__6335\
        );

    \I__478\ : Span12Mux_h
    port map (
            O => \N__6348\,
            I => \N__6335\
        );

    \I__477\ : Span4Mux_h
    port map (
            O => \N__6345\,
            I => \N__6332\
        );

    \I__476\ : Odrv12
    port map (
            O => \N__6342\,
            I => \TVP_VIDEO_c_7\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__6335\,
            I => \TVP_VIDEO_c_7\
        );

    \I__474\ : Odrv4
    port map (
            O => \N__6332\,
            I => \TVP_VIDEO_c_7\
        );

    \I__473\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6321\
        );

    \I__472\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6318\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__6321\,
            I => \N__6315\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__6318\,
            I => \N__6311\
        );

    \I__469\ : Span4Mux_v
    port map (
            O => \N__6315\,
            I => \N__6308\
        );

    \I__468\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6305\
        );

    \I__467\ : Span4Mux_v
    port map (
            O => \N__6311\,
            I => \N__6301\
        );

    \I__466\ : Span4Mux_v
    port map (
            O => \N__6308\,
            I => \N__6296\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__6305\,
            I => \N__6296\
        );

    \I__464\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6293\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__6301\,
            I => \N__6290\
        );

    \I__462\ : Span4Mux_v
    port map (
            O => \N__6296\,
            I => \N__6284\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__6293\,
            I => \N__6284\
        );

    \I__460\ : Span4Mux_v
    port map (
            O => \N__6290\,
            I => \N__6280\
        );

    \I__459\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6277\
        );

    \I__458\ : Span4Mux_v
    port map (
            O => \N__6284\,
            I => \N__6273\
        );

    \I__457\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6270\
        );

    \I__456\ : Span4Mux_v
    port map (
            O => \N__6280\,
            I => \N__6265\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6265\
        );

    \I__454\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6262\
        );

    \I__453\ : Span4Mux_v
    port map (
            O => \N__6273\,
            I => \N__6257\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__6270\,
            I => \N__6257\
        );

    \I__451\ : Span4Mux_v
    port map (
            O => \N__6265\,
            I => \N__6252\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__6262\,
            I => \N__6252\
        );

    \I__449\ : Span4Mux_v
    port map (
            O => \N__6257\,
            I => \N__6248\
        );

    \I__448\ : Span4Mux_v
    port map (
            O => \N__6252\,
            I => \N__6245\
        );

    \I__447\ : InMux
    port map (
            O => \N__6251\,
            I => \N__6242\
        );

    \I__446\ : Sp12to4
    port map (
            O => \N__6248\,
            I => \N__6239\
        );

    \I__445\ : Span4Mux_v
    port map (
            O => \N__6245\,
            I => \N__6234\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__6242\,
            I => \N__6234\
        );

    \I__443\ : Span12Mux_h
    port map (
            O => \N__6239\,
            I => \N__6231\
        );

    \I__442\ : Span4Mux_h
    port map (
            O => \N__6234\,
            I => \N__6228\
        );

    \I__441\ : Odrv12
    port map (
            O => \N__6231\,
            I => \TVP_VIDEO_c_6\
        );

    \I__440\ : Odrv4
    port map (
            O => \N__6228\,
            I => \TVP_VIDEO_c_6\
        );

    \I__439\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6219\
        );

    \I__438\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6216\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__6219\,
            I => \N__6212\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__6216\,
            I => \N__6209\
        );

    \I__435\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6206\
        );

    \I__434\ : Sp12to4
    port map (
            O => \N__6212\,
            I => \N__6202\
        );

    \I__433\ : Span4Mux_h
    port map (
            O => \N__6209\,
            I => \N__6199\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__6206\,
            I => \N__6196\
        );

    \I__431\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6192\
        );

    \I__430\ : Span12Mux_h
    port map (
            O => \N__6202\,
            I => \N__6187\
        );

    \I__429\ : Span4Mux_h
    port map (
            O => \N__6199\,
            I => \N__6184\
        );

    \I__428\ : Span4Mux_v
    port map (
            O => \N__6196\,
            I => \N__6181\
        );

    \I__427\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6178\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__6192\,
            I => \N__6175\
        );

    \I__425\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6172\
        );

    \I__424\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6168\
        );

    \I__423\ : Span12Mux_v
    port map (
            O => \N__6187\,
            I => \N__6163\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__6184\,
            I => \N__6163\
        );

    \I__421\ : Sp12to4
    port map (
            O => \N__6181\,
            I => \N__6160\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__6178\,
            I => \N__6157\
        );

    \I__419\ : Span12Mux_h
    port map (
            O => \N__6175\,
            I => \N__6154\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__6172\,
            I => \N__6151\
        );

    \I__417\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6148\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6145\
        );

    \I__415\ : Span12Mux_v
    port map (
            O => \N__6163\,
            I => \N__6140\
        );

    \I__414\ : Span12Mux_h
    port map (
            O => \N__6160\,
            I => \N__6140\
        );

    \I__413\ : Span12Mux_h
    port map (
            O => \N__6157\,
            I => \N__6137\
        );

    \I__412\ : Span12Mux_v
    port map (
            O => \N__6154\,
            I => \N__6130\
        );

    \I__411\ : Span12Mux_h
    port map (
            O => \N__6151\,
            I => \N__6130\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__6148\,
            I => \N__6130\
        );

    \I__409\ : Span4Mux_h
    port map (
            O => \N__6145\,
            I => \N__6127\
        );

    \I__408\ : Span12Mux_h
    port map (
            O => \N__6140\,
            I => \N__6122\
        );

    \I__407\ : Span12Mux_v
    port map (
            O => \N__6137\,
            I => \N__6122\
        );

    \I__406\ : Span12Mux_h
    port map (
            O => \N__6130\,
            I => \N__6117\
        );

    \I__405\ : Sp12to4
    port map (
            O => \N__6127\,
            I => \N__6117\
        );

    \I__404\ : Odrv12
    port map (
            O => \N__6122\,
            I => \TVP_VIDEO_c_3\
        );

    \I__403\ : Odrv12
    port map (
            O => \N__6117\,
            I => \TVP_VIDEO_c_3\
        );

    \I__402\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6108\
        );

    \I__401\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6105\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__6108\,
            I => \N__6102\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__6105\,
            I => \N__6098\
        );

    \I__398\ : Span4Mux_v
    port map (
            O => \N__6102\,
            I => \N__6095\
        );

    \I__397\ : InMux
    port map (
            O => \N__6101\,
            I => \N__6092\
        );

    \I__396\ : Span4Mux_v
    port map (
            O => \N__6098\,
            I => \N__6089\
        );

    \I__395\ : Span4Mux_v
    port map (
            O => \N__6095\,
            I => \N__6083\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__6092\,
            I => \N__6083\
        );

    \I__393\ : Span4Mux_v
    port map (
            O => \N__6089\,
            I => \N__6079\
        );

    \I__392\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6076\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__6083\,
            I => \N__6073\
        );

    \I__390\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6070\
        );

    \I__389\ : Span4Mux_v
    port map (
            O => \N__6079\,
            I => \N__6064\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__6076\,
            I => \N__6064\
        );

    \I__387\ : Span4Mux_v
    port map (
            O => \N__6073\,
            I => \N__6058\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6058\
        );

    \I__385\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6055\
        );

    \I__384\ : Span4Mux_v
    port map (
            O => \N__6064\,
            I => \N__6052\
        );

    \I__383\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6049\
        );

    \I__382\ : Span4Mux_v
    port map (
            O => \N__6058\,
            I => \N__6044\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__6055\,
            I => \N__6044\
        );

    \I__380\ : Span4Mux_v
    port map (
            O => \N__6052\,
            I => \N__6039\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__6049\,
            I => \N__6039\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__6044\,
            I => \N__6035\
        );

    \I__377\ : Span4Mux_v
    port map (
            O => \N__6039\,
            I => \N__6032\
        );

    \I__376\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6029\
        );

    \I__375\ : Sp12to4
    port map (
            O => \N__6035\,
            I => \N__6026\
        );

    \I__374\ : Span4Mux_v
    port map (
            O => \N__6032\,
            I => \N__6021\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__6029\,
            I => \N__6021\
        );

    \I__372\ : Span12Mux_h
    port map (
            O => \N__6026\,
            I => \N__6018\
        );

    \I__371\ : Span4Mux_h
    port map (
            O => \N__6021\,
            I => \N__6015\
        );

    \I__370\ : Odrv12
    port map (
            O => \N__6018\,
            I => \TVP_VIDEO_c_5\
        );

    \I__369\ : Odrv4
    port map (
            O => \N__6015\,
            I => \TVP_VIDEO_c_5\
        );

    \I__368\ : InMux
    port map (
            O => \N__6010\,
            I => \N__6007\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__6007\,
            I => \N__6004\
        );

    \I__366\ : Span4Mux_v
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__365\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5995\
        );

    \I__364\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5991\
        );

    \I__363\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5987\
        );

    \I__362\ : Span4Mux_v
    port map (
            O => \N__5998\,
            I => \N__5982\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__5995\,
            I => \N__5982\
        );

    \I__360\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5979\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__5991\,
            I => \N__5976\
        );

    \I__358\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5973\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__5987\,
            I => \N__5970\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__5982\,
            I => \N__5965\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__5979\,
            I => \N__5965\
        );

    \I__354\ : Span4Mux_h
    port map (
            O => \N__5976\,
            I => \N__5962\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__5973\,
            I => \N__5959\
        );

    \I__352\ : Span4Mux_s1_v
    port map (
            O => \N__5970\,
            I => \N__5955\
        );

    \I__351\ : Span4Mux_v
    port map (
            O => \N__5965\,
            I => \N__5952\
        );

    \I__350\ : Span4Mux_h
    port map (
            O => \N__5962\,
            I => \N__5949\
        );

    \I__349\ : Span4Mux_h
    port map (
            O => \N__5959\,
            I => \N__5946\
        );

    \I__348\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5943\
        );

    \I__347\ : Sp12to4
    port map (
            O => \N__5955\,
            I => \N__5940\
        );

    \I__346\ : Sp12to4
    port map (
            O => \N__5952\,
            I => \N__5937\
        );

    \I__345\ : Span4Mux_h
    port map (
            O => \N__5949\,
            I => \N__5934\
        );

    \I__344\ : Span4Mux_v
    port map (
            O => \N__5946\,
            I => \N__5931\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__5943\,
            I => \N__5928\
        );

    \I__342\ : Span12Mux_s10_h
    port map (
            O => \N__5940\,
            I => \N__5924\
        );

    \I__341\ : Span12Mux_s9_h
    port map (
            O => \N__5937\,
            I => \N__5921\
        );

    \I__340\ : Span4Mux_h
    port map (
            O => \N__5934\,
            I => \N__5914\
        );

    \I__339\ : Span4Mux_v
    port map (
            O => \N__5931\,
            I => \N__5914\
        );

    \I__338\ : Span4Mux_h
    port map (
            O => \N__5928\,
            I => \N__5914\
        );

    \I__337\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5911\
        );

    \I__336\ : Span12Mux_v
    port map (
            O => \N__5924\,
            I => \N__5908\
        );

    \I__335\ : Span12Mux_v
    port map (
            O => \N__5921\,
            I => \N__5905\
        );

    \I__334\ : Span4Mux_v
    port map (
            O => \N__5914\,
            I => \N__5902\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__5911\,
            I => \N__5899\
        );

    \I__332\ : Span12Mux_v
    port map (
            O => \N__5908\,
            I => \N__5896\
        );

    \I__331\ : Span12Mux_h
    port map (
            O => \N__5905\,
            I => \N__5893\
        );

    \I__330\ : Span4Mux_v
    port map (
            O => \N__5902\,
            I => \N__5890\
        );

    \I__329\ : Span4Mux_h
    port map (
            O => \N__5899\,
            I => \N__5887\
        );

    \I__328\ : Odrv12
    port map (
            O => \N__5896\,
            I => \TVP_VIDEO_c_4\
        );

    \I__327\ : Odrv12
    port map (
            O => \N__5893\,
            I => \TVP_VIDEO_c_4\
        );

    \I__326\ : Odrv4
    port map (
            O => \N__5890\,
            I => \TVP_VIDEO_c_4\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__5887\,
            I => \TVP_VIDEO_c_4\
        );

    \INVADV_R__i2C\ : INV
    port map (
            O => \INVADV_R__i2C_net\,
            I => \N__17333\
        );

    \INVADV_R__i6C\ : INV
    port map (
            O => \INVADV_R__i6C_net\,
            I => \N__17196\
        );

    \INVADV_R__i3C\ : INV
    port map (
            O => \INVADV_R__i3C_net\,
            I => \N__17411\
        );

    \INVADV_R__i1C\ : INV
    port map (
            O => \INVADV_R__i1C_net\,
            I => \N__17495\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n2773\,
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.n2747\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n2765\,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n2789\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.n2734\,
            carryinitout => \bfn_18_15_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__18151\,
            in1 => \N__18070\,
            in2 => \N__17972\,
            in3 => \N__17780\,
            lcout => \line_buffer.n730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1639_2_lut_3_lut_4_lut_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17812\,
            in1 => \N__18139\,
            in2 => \N__17971\,
            in3 => \N__18068\,
            lcout => \line_buffer.n632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18069\,
            in1 => \N__17952\,
            in2 => \N__18149\,
            in3 => \N__17811\,
            lcout => \line_buffer.n762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1584_3_lut_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18474\,
            in1 => \N__7021\,
            in2 => \_gnd_net_\,
            in3 => \N__7009\,
            lcout => \line_buffer.n3028\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7101\,
            in1 => \N__7118\,
            in2 => \_gnd_net_\,
            in3 => \N__6949\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n2975_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i38_4_lut_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010111001"
        )
    port map (
            in0 => \N__7060\,
            in1 => \N__7081\,
            in2 => \N__6997\,
            in3 => \N__6940\,
            lcout => \receive_module.rx_counter.n31_adj_572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18150\,
            in1 => \N__18067\,
            in2 => \N__17980\,
            in3 => \N__17762\,
            lcout => \line_buffer.n698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_adj_19_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7164\,
            in1 => \N__7134\,
            in2 => \_gnd_net_\,
            in3 => \N__7149\,
            lcout => \receive_module.rx_counter.n2900\,
            ltout => \receive_module.rx_counter.n2900_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1499_3_lut_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__7119\,
            in1 => \_gnd_net_\,
            in2 => \N__6943\,
            in3 => \N__7102\,
            lcout => \receive_module.rx_counter.n2943\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.X_284__i0_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6934\,
            in2 => \_gnd_net_\,
            in3 => \N__6928\,
            lcout => \receive_module.rx_counter.n10\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \receive_module.rx_counter.n2782\,
            clk => \N__16101\,
            ce => 'H',
            sr => \N__7044\
        );

    \receive_module.rx_counter.X_284__i1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6925\,
            in2 => \_gnd_net_\,
            in3 => \N__6919\,
            lcout => \receive_module.rx_counter.n9\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2782\,
            carryout => \receive_module.rx_counter.n2783\,
            clk => \N__16101\,
            ce => 'H',
            sr => \N__7044\
        );

    \receive_module.rx_counter.X_284__i2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6916\,
            in2 => \_gnd_net_\,
            in3 => \N__6910\,
            lcout => \receive_module.rx_counter.n8\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2783\,
            carryout => \receive_module.rx_counter.n2784\,
            clk => \N__16101\,
            ce => 'H',
            sr => \N__7044\
        );

    \receive_module.rx_counter.X_284__i3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7165\,
            in2 => \_gnd_net_\,
            in3 => \N__7153\,
            lcout => \receive_module.rx_counter.X_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2784\,
            carryout => \receive_module.rx_counter.n2785\,
            clk => \N__16101\,
            ce => 'H',
            sr => \N__7044\
        );

    \receive_module.rx_counter.X_284__i4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7150\,
            in2 => \_gnd_net_\,
            in3 => \N__7138\,
            lcout => \receive_module.rx_counter.X_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2785\,
            carryout => \receive_module.rx_counter.n2786\,
            clk => \N__16101\,
            ce => 'H',
            sr => \N__7044\
        );

    \receive_module.rx_counter.X_284__i5_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7135\,
            in2 => \_gnd_net_\,
            in3 => \N__7123\,
            lcout => \receive_module.rx_counter.X_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2786\,
            carryout => \receive_module.rx_counter.n2787\,
            clk => \N__16101\,
            ce => 'H',
            sr => \N__7044\
        );

    \receive_module.rx_counter.X_284__i6_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7120\,
            in2 => \_gnd_net_\,
            in3 => \N__7105\,
            lcout => \receive_module.rx_counter.X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2787\,
            carryout => \receive_module.rx_counter.n2788\,
            clk => \N__16101\,
            ce => 'H',
            sr => \N__7044\
        );

    \receive_module.rx_counter.X_284__i7_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7100\,
            in2 => \_gnd_net_\,
            in3 => \N__7084\,
            lcout => \receive_module.rx_counter.X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2788\,
            carryout => \receive_module.rx_counter.n2789\,
            clk => \N__16101\,
            ce => 'H',
            sr => \N__7044\
        );

    \receive_module.rx_counter.X_284__i8_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7080\,
            in2 => \_gnd_net_\,
            in3 => \N__7066\,
            lcout => \receive_module.rx_counter.X_8\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \receive_module.rx_counter.n2790\,
            clk => \N__16103\,
            ce => 'H',
            sr => \N__7045\
        );

    \receive_module.rx_counter.X_284__i9_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7059\,
            in2 => \_gnd_net_\,
            in3 => \N__7063\,
            lcout => \receive_module.rx_counter.X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16103\,
            ce => 'H',
            sr => \N__7045\
        );

    \i27_1_lut_rep_20_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n3184,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7372\,
            in2 => \_gnd_net_\,
            in3 => \N__7228\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_adj_17_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__7732\,
            in1 => \N__7702\,
            in2 => \N__7207\,
            in3 => \N__7423\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n2986_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i4_4_lut_adj_18_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7475\,
            in1 => \N__7192\,
            in2 => \N__7204\,
            in3 => \N__7400\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n2989_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_adj_20_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001111"
        )
    port map (
            in0 => \N__7250\,
            in1 => \N__7177\,
            in2 => \N__7201\,
            in3 => \N__7198\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7447\,
            in2 => \_gnd_net_\,
            in3 => \N__7249\,
            lcout => \receive_module.rx_counter.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_rep_2_2_lut_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7448\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7474\,
            lcout => \receive_module.rx_counter.n3166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__7424\,
            in1 => \N__7703\,
            in2 => \N__7737\,
            in3 => \N__7373\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n2978_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_4_lut_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__7229\,
            in1 => \N__7186\,
            in2 => \N__7180\,
            in3 => \N__7399\,
            lcout => \receive_module.rx_counter.n4_adj_571\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.Y__i0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7733\,
            in2 => \_gnd_net_\,
            in3 => \N__7171\,
            lcout => \Y_0\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \receive_module.rx_counter.n2758\,
            clk => \N__16092\,
            ce => \N__7539\,
            sr => \N__15979\
        );

    \receive_module.rx_counter.Y__i1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7704\,
            in2 => \_gnd_net_\,
            in3 => \N__7168\,
            lcout => \Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2758\,
            carryout => \receive_module.rx_counter.n2759\,
            clk => \N__16092\,
            ce => \N__7539\,
            sr => \N__15979\
        );

    \receive_module.rx_counter.Y__i2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7425\,
            in2 => \_gnd_net_\,
            in3 => \N__7276\,
            lcout => \receive_module.rx_counter.Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2759\,
            carryout => \receive_module.rx_counter.n2760\,
            clk => \N__16092\,
            ce => \N__7539\,
            sr => \N__15979\
        );

    \receive_module.rx_counter.Y__i3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7374\,
            in2 => \_gnd_net_\,
            in3 => \N__7273\,
            lcout => \receive_module.rx_counter.Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2760\,
            carryout => \receive_module.rx_counter.n2761\,
            clk => \N__16092\,
            ce => \N__7539\,
            sr => \N__15979\
        );

    \receive_module.rx_counter.Y__i4_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7230\,
            in2 => \_gnd_net_\,
            in3 => \N__7270\,
            lcout => \receive_module.rx_counter.Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2761\,
            carryout => \receive_module.rx_counter.n2762\,
            clk => \N__16092\,
            ce => \N__7539\,
            sr => \N__15979\
        );

    \receive_module.rx_counter.Y__i5_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7476\,
            in2 => \_gnd_net_\,
            in3 => \N__7267\,
            lcout => \receive_module.rx_counter.Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2762\,
            carryout => \receive_module.rx_counter.n2763\,
            clk => \N__16092\,
            ce => \N__7539\,
            sr => \N__15979\
        );

    \receive_module.rx_counter.Y__i6_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7449\,
            in2 => \_gnd_net_\,
            in3 => \N__7264\,
            lcout => \receive_module.rx_counter.Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2763\,
            carryout => \receive_module.rx_counter.n2764\,
            clk => \N__16092\,
            ce => \N__7539\,
            sr => \N__15979\
        );

    \receive_module.rx_counter.Y__i7_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7251\,
            in2 => \_gnd_net_\,
            in3 => \N__7261\,
            lcout => \receive_module.rx_counter.Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2764\,
            carryout => \receive_module.rx_counter.n2765\,
            clk => \N__16092\,
            ce => \N__7539\,
            sr => \N__15979\
        );

    \receive_module.rx_counter.Y__i8_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7401\,
            in2 => \_gnd_net_\,
            in3 => \N__7258\,
            lcout => \receive_module.rx_counter.Y_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16096\,
            ce => \N__7540\,
            sr => \N__15964\
        );

    \transmit_module.video_signal_controller.i1570_4_lut_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__8656\,
            in1 => \N__8691\,
            in2 => \N__7327\,
            in3 => \N__8026\,
            lcout => \transmit_module.video_signal_controller.n3014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_21_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7255\,
            in2 => \_gnd_net_\,
            in3 => \N__7231\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i4_4_lut_adj_22_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__7426\,
            in1 => \N__7402\,
            in2 => \N__7378\,
            in3 => \N__7375\,
            lcout => n3009,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i3_3_lut_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7641\,
            in1 => \N__7625\,
            in2 => \_gnd_net_\,
            in3 => \N__7603\,
            lcout => \transmit_module.video_signal_controller.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1596_3_lut_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18441\,
            in1 => \N__7351\,
            in2 => \_gnd_net_\,
            in3 => \N__7339\,
            lcout => \line_buffer.n3040\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__8050\,
            in1 => \N__7604\,
            in2 => \_gnd_net_\,
            in3 => \N__8081\,
            lcout => \transmit_module.video_signal_controller.n2972\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__8024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8083\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_HS_48_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__7291\,
            in1 => \N__7318\,
            in2 => \N__7312\,
            in3 => \N__8110\,
            lcout => \ADV_HSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i541_3_lut_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__7605\,
            in1 => \N__7627\,
            in2 => \_gnd_net_\,
            in3 => \N__8051\,
            lcout => \transmit_module.video_signal_controller.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_18_3_lut_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__8049\,
            in1 => \N__8080\,
            in2 => \_gnd_net_\,
            in3 => \N__8023\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3182_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1127_4_lut_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7671\,
            in1 => \N__7656\,
            in2 => \N__7285\,
            in3 => \N__7282\,
            lcout => \transmit_module.video_signal_controller.n2484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i9_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7762\,
            lcout => \transmit_module.X_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17424\,
            ce => \N__9961\,
            sr => \N__14404\
        );

    \transmit_module.X_DELTA_PATTERN_i8_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7576\,
            lcout => \transmit_module.X_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17424\,
            ce => \N__9961\,
            sr => \N__14404\
        );

    \transmit_module.X_DELTA_PATTERN_i7_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7570\,
            lcout => \transmit_module.X_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17424\,
            ce => \N__9961\,
            sr => \N__14404\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1661_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__18440\,
            in1 => \N__7564\,
            in2 => \N__15809\,
            in3 => \N__7552\,
            lcout => \line_buffer.n3101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i297_3_lut_3_lut_3_lut_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__7523\,
            in1 => \N__7489\,
            in2 => \_gnd_net_\,
            in3 => \N__16471\,
            lcout => \receive_module.n2152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_HS_48_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.old_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1145_4_lut_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__8655\,
            in1 => \N__7483\,
            in2 => \N__8692\,
            in3 => \N__8109\,
            lcout => n2147,
            ltout => \n2147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_3_lut_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7477\,
            in2 => \N__7453\,
            in3 => \N__7450\,
            lcout => OPEN,
            ltout => \n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1642_4_lut_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7738\,
            in1 => \N__7708\,
            in2 => \N__7681\,
            in3 => \N__7678\,
            lcout => \transmit_module.video_signal_controller.n2262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i1_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7672\,
            in2 => \_gnd_net_\,
            in3 => \N__7660\,
            lcout => \transmit_module.video_signal_controller.VGA_X_0\,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \transmit_module.video_signal_controller.n2766\,
            clk => \N__17516\,
            ce => 'H',
            sr => \N__8158\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i2_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7657\,
            in2 => \_gnd_net_\,
            in3 => \N__7645\,
            lcout => \transmit_module.video_signal_controller.VGA_X_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2766\,
            carryout => \transmit_module.video_signal_controller.n2767\,
            clk => \N__17516\,
            ce => 'H',
            sr => \N__8158\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i3_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7642\,
            in2 => \_gnd_net_\,
            in3 => \N__7630\,
            lcout => \transmit_module.video_signal_controller.VGA_X_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2767\,
            carryout => \transmit_module.video_signal_controller.n2768\,
            clk => \N__17516\,
            ce => 'H',
            sr => \N__8158\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i4_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7626\,
            in2 => \_gnd_net_\,
            in3 => \N__7609\,
            lcout => \transmit_module.video_signal_controller.VGA_X_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2768\,
            carryout => \transmit_module.video_signal_controller.n2769\,
            clk => \N__17516\,
            ce => 'H',
            sr => \N__8158\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i5_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7606\,
            in2 => \_gnd_net_\,
            in3 => \N__7588\,
            lcout => \transmit_module.video_signal_controller.VGA_X_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2769\,
            carryout => \transmit_module.video_signal_controller.n2770\,
            clk => \N__17516\,
            ce => 'H',
            sr => \N__8158\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i6_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8052\,
            in2 => \_gnd_net_\,
            in3 => \N__7585\,
            lcout => \transmit_module.video_signal_controller.VGA_X_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2770\,
            carryout => \transmit_module.video_signal_controller.n2771\,
            clk => \N__17516\,
            ce => 'H',
            sr => \N__8158\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i7_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8082\,
            in2 => \_gnd_net_\,
            in3 => \N__7582\,
            lcout => \transmit_module.video_signal_controller.VGA_X_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2771\,
            carryout => \transmit_module.video_signal_controller.n2772\,
            clk => \N__17516\,
            ce => 'H',
            sr => \N__8158\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i8_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8025\,
            in2 => \_gnd_net_\,
            in3 => \N__7579\,
            lcout => \transmit_module.video_signal_controller.VGA_X_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2772\,
            carryout => \transmit_module.video_signal_controller.n2773\,
            clk => \N__17516\,
            ce => 'H',
            sr => \N__8158\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i9_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8108\,
            in2 => \_gnd_net_\,
            in3 => \N__7777\,
            lcout => \transmit_module.video_signal_controller.VGA_X_8\,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \transmit_module.video_signal_controller.n2774\,
            clk => \N__17474\,
            ce => 'H',
            sr => \N__8157\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i10_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8686\,
            in2 => \_gnd_net_\,
            in3 => \N__7774\,
            lcout => \transmit_module.video_signal_controller.VGA_X_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2774\,
            carryout => \transmit_module.video_signal_controller.n2775\,
            clk => \N__17474\,
            ce => 'H',
            sr => \N__8157\
        );

    \transmit_module.video_signal_controller.VGA_X_288_289__i11_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8653\,
            in2 => \_gnd_net_\,
            in3 => \N__7771\,
            lcout => \transmit_module.video_signal_controller.VGA_X_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17474\,
            ce => 'H',
            sr => \N__8157\
        );

    \transmit_module.X_DELTA_PATTERN_i12_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7768\,
            lcout => \transmit_module.X_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17423\,
            ce => \N__9955\,
            sr => \N__14413\
        );

    \transmit_module.X_DELTA_PATTERN_i13_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7960\,
            lcout => \transmit_module.X_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17423\,
            ce => \N__9955\,
            sr => \N__14413\
        );

    \transmit_module.X_DELTA_PATTERN_i15_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8613\,
            lcout => \transmit_module.X_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17423\,
            ce => \N__9955\,
            sr => \N__14413\
        );

    \transmit_module.X_DELTA_PATTERN_i10_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7750\,
            lcout => \transmit_module.X_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17423\,
            ce => \N__9955\,
            sr => \N__14413\
        );

    \transmit_module.X_DELTA_PATTERN_i11_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7756\,
            lcout => \transmit_module.X_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17423\,
            ce => \N__9955\,
            sr => \N__14413\
        );

    \transmit_module.X_DELTA_PATTERN_i6_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7744\,
            lcout => \transmit_module.X_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17423\,
            ce => \N__9955\,
            sr => \N__14413\
        );

    \transmit_module.X_DELTA_PATTERN_i14_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7966\,
            lcout => \transmit_module.X_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17423\,
            ce => \N__9955\,
            sr => \N__14413\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1696_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__18393\,
            in1 => \N__7954\,
            in2 => \N__15781\,
            in3 => \N__7945\,
            lcout => OPEN,
            ltout => \line_buffer.n3143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3143_bdd_4_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__7930\,
            in1 => \N__15745\,
            in2 => \N__7915\,
            in3 => \N__7912\,
            lcout => \line_buffer.n3146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3101_bdd_4_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__7891\,
            in1 => \N__15772\,
            in2 => \N__7876\,
            in3 => \N__7855\,
            lcout => \line_buffer.n3104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1586_3_lut_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18471\,
            in1 => \N__7849\,
            in2 => \_gnd_net_\,
            in3 => \N__7831\,
            lcout => \line_buffer.n3030\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1656_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__18487\,
            in1 => \N__7819\,
            in2 => \N__15810\,
            in3 => \N__7804\,
            lcout => \line_buffer.n3089\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_Y_286_287__i1_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8124\,
            in2 => \_gnd_net_\,
            in3 => \N__7786\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_0\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \transmit_module.video_signal_controller.n2776\,
            clk => \N__17496\,
            ce => \N__8153\,
            sr => \N__8131\
        );

    \transmit_module.video_signal_controller.VGA_Y_286_287__i2_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7999\,
            in2 => \_gnd_net_\,
            in3 => \N__7783\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2776\,
            carryout => \transmit_module.video_signal_controller.n2777\,
            clk => \N__17496\,
            ce => \N__8153\,
            sr => \N__8131\
        );

    \transmit_module.video_signal_controller.VGA_Y_286_287__i3_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7983\,
            in2 => \_gnd_net_\,
            in3 => \N__7780\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2777\,
            carryout => \transmit_module.video_signal_controller.n2778\,
            clk => \N__17496\,
            ce => \N__8153\,
            sr => \N__8131\
        );

    \transmit_module.video_signal_controller.VGA_Y_286_287__i4_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8717\,
            in2 => \_gnd_net_\,
            in3 => \N__8170\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2778\,
            carryout => \transmit_module.video_signal_controller.n2779\,
            clk => \N__17496\,
            ce => \N__8153\,
            sr => \N__8131\
        );

    \transmit_module.video_signal_controller.VGA_Y_286_287__i5_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8751\,
            in2 => \_gnd_net_\,
            in3 => \N__8167\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2779\,
            carryout => \transmit_module.video_signal_controller.n2780\,
            clk => \N__17496\,
            ce => \N__8153\,
            sr => \N__8131\
        );

    \transmit_module.video_signal_controller.VGA_Y_286_287__i6_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8263\,
            in2 => \_gnd_net_\,
            in3 => \N__8164\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n2780\,
            carryout => \transmit_module.video_signal_controller.n2781\,
            clk => \N__17496\,
            ce => \N__8153\,
            sr => \N__8131\
        );

    \transmit_module.video_signal_controller.VGA_Y_286_287__i7_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8245\,
            in2 => \_gnd_net_\,
            in3 => \N__8161\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17496\,
            ce => \N__8153\,
            sr => \N__8131\
        );

    \transmit_module.video_signal_controller.i1578_3_lut_4_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8244\,
            in1 => \N__8750\,
            in2 => \N__8724\,
            in3 => \N__8262\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3022_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VS_49_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__7998\,
            in1 => \N__8125\,
            in2 => \N__8113\,
            in3 => \N__7984\,
            lcout => \ADV_VSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i511_2_lut_3_lut_4_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__8101\,
            in1 => \N__8079\,
            in2 => \N__8056\,
            in3 => \N__8022\,
            lcout => \transmit_module.video_signal_controller.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i508_2_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7997\,
            in2 => \_gnd_net_\,
            in3 => \N__7982\,
            lcout => \transmit_module.video_signal_controller.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8261\,
            in2 => \_gnd_net_\,
            in3 => \N__8243\,
            lcout => \transmit_module.video_signal_controller.n3183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8230\,
            lcout => \transmit_module.X_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17436\,
            ce => \N__9956\,
            sr => \N__14440\
        );

    \transmit_module.X_DELTA_PATTERN_i1_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8224\,
            lcout => \transmit_module.X_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17436\,
            ce => \N__9956\,
            sr => \N__14440\
        );

    \transmit_module.X_DELTA_PATTERN_i2_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8200\,
            lcout => \transmit_module.X_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17436\,
            ce => \N__9956\,
            sr => \N__14440\
        );

    \transmit_module.X_DELTA_PATTERN_i5_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8218\,
            lcout => \transmit_module.X_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17436\,
            ce => \N__9956\,
            sr => \N__14440\
        );

    \transmit_module.X_DELTA_PATTERN_i4_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8212\,
            lcout => \transmit_module.X_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17436\,
            ce => \N__9956\,
            sr => \N__14440\
        );

    \transmit_module.X_DELTA_PATTERN_i3_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8206\,
            lcout => \transmit_module.X_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17436\,
            ce => \N__9956\,
            sr => \N__14440\
        );

    \transmit_module.i1_2_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14348\,
            in2 => \_gnd_net_\,
            in3 => \N__14131\,
            lcout => \transmit_module.n2200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1587_3_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18386\,
            in1 => \N__8194\,
            in2 => \_gnd_net_\,
            in3 => \N__8185\,
            lcout => OPEN,
            ltout => \line_buffer.n3031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_1676_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__17635\,
            in1 => \N__15723\,
            in2 => \N__8389\,
            in3 => \N__8386\,
            lcout => OPEN,
            ltout => \line_buffer.n3095_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i3_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__17651\,
            in1 => \N__8275\,
            in2 => \N__8377\,
            in3 => \N__8374\,
            lcout => \TX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17446\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i7_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__14411\,
            in1 => \N__9897\,
            in2 => \N__9930\,
            in3 => \N__14172\,
            lcout => \DEBUG_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i11_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__14171\,
            in1 => \N__10634\,
            in2 => \N__10612\,
            in3 => \N__14412\,
            lcout => \transmit_module.TX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3089_bdd_4_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001100"
        )
    port map (
            in0 => \N__8362\,
            in1 => \N__8344\,
            in2 => \N__15768\,
            in3 => \N__8323\,
            lcout => OPEN,
            ltout => \line_buffer.n3092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i2_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17650\,
            in2 => \N__8314\,
            in3 => \N__8311\,
            lcout => \TX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1595_3_lut_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8305\,
            in1 => \N__8293\,
            in2 => \_gnd_net_\,
            in3 => \N__18439\,
            lcout => \line_buffer.n3039\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i4_4_lut_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__8538\,
            in1 => \N__8553\,
            in2 => \N__8587\,
            in3 => \N__8568\,
            lcout => \receive_module.rx_counter.n10_adj_570\,
            ltout => \receive_module.rx_counter.n10_adj_570_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i873_2_lut_4_lut_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8846\,
            in1 => \N__8819\,
            in2 => \N__8266\,
            in3 => \N__10334\,
            lcout => \receive_module.rx_counter.n2227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.FRAME_COUNTER_285__i0_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8820\,
            in2 => \_gnd_net_\,
            in3 => \N__8590\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_0\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \receive_module.rx_counter.n2753\,
            clk => \N__16084\,
            ce => \N__10341\,
            sr => \N__8521\
        );

    \receive_module.rx_counter.FRAME_COUNTER_285__i1_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8586\,
            in2 => \_gnd_net_\,
            in3 => \N__8572\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2753\,
            carryout => \receive_module.rx_counter.n2754\,
            clk => \N__16084\,
            ce => \N__10341\,
            sr => \N__8521\
        );

    \receive_module.rx_counter.FRAME_COUNTER_285__i2_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8569\,
            in2 => \_gnd_net_\,
            in3 => \N__8557\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2754\,
            carryout => \receive_module.rx_counter.n2755\,
            clk => \N__16084\,
            ce => \N__10341\,
            sr => \N__8521\
        );

    \receive_module.rx_counter.FRAME_COUNTER_285__i3_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8554\,
            in2 => \_gnd_net_\,
            in3 => \N__8542\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2755\,
            carryout => \receive_module.rx_counter.n2756\,
            clk => \N__16084\,
            ce => \N__10341\,
            sr => \N__8521\
        );

    \receive_module.rx_counter.FRAME_COUNTER_285__i4_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8539\,
            in2 => \_gnd_net_\,
            in3 => \N__8527\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n2756\,
            carryout => \receive_module.rx_counter.n2757\,
            clk => \N__16084\,
            ce => \N__10341\,
            sr => \N__8521\
        );

    \receive_module.rx_counter.FRAME_COUNTER_285__i5_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8848\,
            in2 => \_gnd_net_\,
            in3 => \N__8524\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16084\,
            ce => \N__10341\,
            sr => \N__8521\
        );

    \receive_module.i24_1_lut_rep_21_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16386\,
            lcout => \receive_module.n3185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADV_R__i1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12220\,
            lcout => n1955,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__14184\
        );

    \ADV_R__i3_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8452\,
            lcout => n1953,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i3C_net\,
            ce => 'H',
            sr => \N__14130\
        );

    \transmit_module.BRAM_ADDR__i5_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__9384\,
            in1 => \N__9362\,
            in2 => \N__14360\,
            in3 => \N__14140\,
            lcout => \DEBUG_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__8752\,
            in1 => \N__8731\,
            in2 => \N__8725\,
            in3 => \N__8698\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.VGA_VISIBLE_N_558_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1636_4_lut_4_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110011111"
        )
    port map (
            in0 => \N__8687\,
            in1 => \N__8654\,
            in2 => \N__8626\,
            in3 => \N__8623\,
            lcout => \VGA_VISIBLE\,
            ltout => \VGA_VISIBLE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i3_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__14296\,
            in1 => \N__9126\,
            in2 => \N__8617\,
            in3 => \N__9092\,
            lcout => \DEBUG_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i6_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__9657\,
            in1 => \N__9626\,
            in2 => \N__14361\,
            in3 => \N__14141\,
            lcout => \DEBUG_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_2_lut_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14206\,
            in2 => \N__8614\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n388\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \transmit_module.n2740\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_3_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12085\,
            in2 => \_gnd_net_\,
            in3 => \N__8599\,
            lcout => \transmit_module.n387\,
            ltout => OPEN,
            carryin => \transmit_module.n2740\,
            carryout => \transmit_module.n2741\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_4_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9088\,
            in2 => \_gnd_net_\,
            in3 => \N__8596\,
            lcout => \transmit_module.n386\,
            ltout => OPEN,
            carryin => \transmit_module.n2741\,
            carryout => \transmit_module.n2742\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_5_lut_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11530\,
            in2 => \_gnd_net_\,
            in3 => \N__8593\,
            lcout => \transmit_module.n385\,
            ltout => OPEN,
            carryin => \transmit_module.n2742\,
            carryout => \transmit_module.n2743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_6_lut_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9358\,
            in2 => \_gnd_net_\,
            in3 => \N__8779\,
            lcout => \transmit_module.n384\,
            ltout => OPEN,
            carryin => \transmit_module.n2743\,
            carryout => \transmit_module.n2744\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_7_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9622\,
            in2 => \_gnd_net_\,
            in3 => \N__8776\,
            lcout => \transmit_module.n383\,
            ltout => OPEN,
            carryin => \transmit_module.n2744\,
            carryout => \transmit_module.n2745\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_8_lut_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9929\,
            in3 => \N__8773\,
            lcout => \transmit_module.n382\,
            ltout => OPEN,
            carryin => \transmit_module.n2745\,
            carryout => \transmit_module.n2746\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_9_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11833\,
            in2 => \_gnd_net_\,
            in3 => \N__8770\,
            lcout => \transmit_module.n381\,
            ltout => OPEN,
            carryin => \transmit_module.n2746\,
            carryout => \transmit_module.n2747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_10_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10880\,
            in2 => \_gnd_net_\,
            in3 => \N__8767\,
            lcout => \transmit_module.n380\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \transmit_module.n2748\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_11_lut_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10902\,
            in3 => \N__8764\,
            lcout => \transmit_module.n379\,
            ltout => OPEN,
            carryin => \transmit_module.n2748\,
            carryout => \transmit_module.n2749\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_15_12_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10635\,
            in3 => \N__8761\,
            lcout => \transmit_module.n378\,
            ltout => OPEN,
            carryin => \transmit_module.n2749\,
            carryout => \transmit_module.n2750\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18385\,
            in2 => \_gnd_net_\,
            in3 => \N__8758\,
            lcout => \TX_ADDR_11\,
            ltout => OPEN,
            carryin => \transmit_module.n2750\,
            carryout => \transmit_module.n2751\,
            clk => \N__17330\,
            ce => \N__9960\,
            sr => \N__14445\
        );

    \transmit_module.BRAM_ADDR__rep_1_i1_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15719\,
            in2 => \_gnd_net_\,
            in3 => \N__8755\,
            lcout => \TX_ADDR_12\,
            ltout => OPEN,
            carryin => \transmit_module.n2751\,
            carryout => \transmit_module.n2752\,
            clk => \N__17330\,
            ce => \N__9960\,
            sr => \N__14445\
        );

    \transmit_module.BRAM_ADDR__rep_1_i2_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17649\,
            in2 => \_gnd_net_\,
            in3 => \N__9964\,
            lcout => \TX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17330\,
            ce => \N__9960\,
            sr => \N__14445\
        );

    \transmit_module.i1056_4_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__9922\,
            in1 => \N__9898\,
            in2 => \N__14425\,
            in3 => \N__14164\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1057_4_lut_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__9658\,
            in1 => \N__9630\,
            in2 => \N__14427\,
            in3 => \N__14166\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1058_4_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__9388\,
            in1 => \N__9366\,
            in2 => \N__14426\,
            in3 => \N__14165\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i9_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__14167\,
            in1 => \N__14384\,
            in2 => \N__10864\,
            in3 => \N__10882\,
            lcout => \transmit_module.TX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1060_4_lut_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__9127\,
            in1 => \N__9102\,
            in2 => \N__14444\,
            in3 => \N__14185\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.PULSE_1HZ_46_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100100000"
        )
    port map (
            in0 => \N__8847\,
            in1 => \N__8830\,
            in2 => \N__8824\,
            in3 => \N__8790\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16080\,
            ce => \N__10345\,
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_VS_49_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.old_VS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i141_2_lut_2_lut_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10351\,
            in2 => \_gnd_net_\,
            in3 => \N__16405\,
            lcout => \receive_module.n252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADV_R__i6_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14803\,
            lcout => n1950,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i6C_net\,
            ce => 'H',
            sr => \N__14101\
        );

    \transmit_module.BRAM_ADDR__i4_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__11571\,
            in1 => \N__14398\,
            in2 => \N__11541\,
            in3 => \N__14139\,
            lcout => \DEBUG_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADV_R__i2_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11194\,
            lcout => n1954,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14102\
        );

    \ADV_R__i4_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10207\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n1952,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14102\
        );

    \ADV_R__i5_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n1951,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14102\
        );

    \ADV_R__i7_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10375\,
            lcout => n1949,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14102\
        );

    \ADV_R__i8_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11284\,
            lcout => \ADV_B_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14102\
        );

    \transmit_module.BRAM_ADDR__i2_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__14173\,
            in1 => \N__12114\,
            in2 => \N__14436\,
            in3 => \N__12093\,
            lcout => \DEBUG_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i1_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__14466\,
            in1 => \N__14174\,
            in2 => \N__14219\,
            in3 => \N__14402\,
            lcout => \DEBUG_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i8_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__11835\,
            in1 => \N__14175\,
            in2 => \N__11811\,
            in3 => \N__14403\,
            lcout => \DEBUG_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1053_4_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__14180\,
            in1 => \N__10898\,
            in2 => \N__14434\,
            in3 => \N__10911\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i10_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__10912\,
            in1 => \N__14397\,
            in2 => \N__10903\,
            in3 => \N__14182\,
            lcout => \transmit_module.TX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1054_4_lut_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__14181\,
            in1 => \N__10881\,
            in2 => \N__14435\,
            in3 => \N__10860\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1052_4_lut_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__10639\,
            in1 => \N__10608\,
            in2 => \N__14424\,
            in3 => \N__14179\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i6_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17668\,
            in1 => \N__10384\,
            in2 => \_gnd_net_\,
            in3 => \N__12679\,
            lcout => \TX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16129\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_TVP_CLK_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i1632_2_lut_rep_17_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__17861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16432\,
            lcout => \receive_module.n3181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i9_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__17869\,
            in1 => \N__16445\,
            in2 => \N__14506\,
            in3 => \N__14530\,
            lcout => \RX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16087\,
            ce => 'H',
            sr => \N__15965\
        );

    \receive_module.BRAM_ADDR__i8_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__12775\,
            in1 => \N__12751\,
            in2 => \N__16470\,
            in3 => \N__17868\,
            lcout => \RX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16087\,
            ce => 'H',
            sr => \N__15965\
        );

    \receive_module.BRAM_ADDR__i7_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__17867\,
            in1 => \N__12997\,
            in2 => \N__16481\,
            in3 => \N__13021\,
            lcout => \RX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16087\,
            ce => 'H',
            sr => \N__15965\
        );

    \receive_module.BRAM_ADDR__i5_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__17866\,
            in1 => \N__16444\,
            in2 => \N__13274\,
            in3 => \N__13246\,
            lcout => \RX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16087\,
            ce => 'H',
            sr => \N__15965\
        );

    \receive_module.BRAM_ADDR__i0_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__16443\,
            in1 => \N__13507\,
            in2 => \N__13544\,
            in3 => \N__17865\,
            lcout => \RX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16087\,
            ce => 'H',
            sr => \N__15965\
        );

    \line_buffer.n3137_bdd_4_lut_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__11239\,
            in1 => \N__15777\,
            in2 => \N__11218\,
            in3 => \N__12172\,
            lcout => OPEN,
            ltout => \line_buffer.n3140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i1_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17684\,
            in2 => \N__11197\,
            in3 => \N__11134\,
            lcout => \TX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1666_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__18470\,
            in1 => \N__11188\,
            in2 => \N__15830\,
            in3 => \N__11179\,
            lcout => OPEN,
            ltout => \line_buffer.n3107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3107_bdd_4_lut_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__11161\,
            in1 => \N__11149\,
            in2 => \N__11137\,
            in3 => \N__15808\,
            lcout => \line_buffer.n3110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1691_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__18469\,
            in1 => \N__12208\,
            in2 => \N__12193\,
            in3 => \N__15807\,
            lcout => \line_buffer.n3137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__18137\,
            in1 => \N__18046\,
            in2 => \N__17979\,
            in3 => \N__17878\,
            lcout => \line_buffer.n761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1061_4_lut_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__12118\,
            in1 => \N__12086\,
            in2 => \N__14443\,
            in3 => \N__14178\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1055_4_lut_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__11834\,
            in1 => \N__11812\,
            in2 => \N__14441\,
            in3 => \N__14176\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1059_4_lut_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__11575\,
            in1 => \N__11540\,
            in2 => \N__14442\,
            in3 => \N__14177\,
            lcout => n25_adj_573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_1681_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__15776\,
            in1 => \N__11296\,
            in2 => \N__17685\,
            in3 => \N__13753\,
            lcout => OPEN,
            ltout => \line_buffer.n3125_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i7_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__12640\,
            in1 => \N__17672\,
            in2 => \N__11287\,
            in3 => \N__11245\,
            lcout => \TX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1599_3_lut_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11275\,
            in1 => \N__11260\,
            in2 => \_gnd_net_\,
            in3 => \N__18450\,
            lcout => \line_buffer.n3043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__18451\,
            in1 => \N__12742\,
            in2 => \N__15812\,
            in3 => \N__12727\,
            lcout => OPEN,
            ltout => \line_buffer.n3161_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3161_bdd_4_lut_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__12712\,
            in1 => \N__12700\,
            in2 => \N__12682\,
            in3 => \N__15785\,
            lcout => \line_buffer.n3164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1598_3_lut_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12673\,
            in1 => \N__12658\,
            in2 => \_gnd_net_\,
            in3 => \N__18475\,
            lcout => \line_buffer.n3042\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_18_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3113_bdd_4_lut_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__15825\,
            in1 => \N__12343\,
            in2 => \N__12325\,
            in3 => \N__12271\,
            lcout => \line_buffer.n3116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1671_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__18477\,
            in1 => \N__12304\,
            in2 => \N__15836\,
            in3 => \N__12289\,
            lcout => \line_buffer.n3113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3119_bdd_4_lut_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__12265\,
            in1 => \N__15826\,
            in2 => \N__12247\,
            in3 => \N__13795\,
            lcout => OPEN,
            ltout => \line_buffer.n3122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i0_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17694\,
            in1 => \_gnd_net_\,
            in2 => \N__12229\,
            in3 => \N__12226\,
            lcout => \TX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_2_lut_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13534\,
            in2 => \_gnd_net_\,
            in3 => \N__13501\,
            lcout => \receive_module.n136\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \receive_module.n2727\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_3_lut_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14873\,
            in2 => \_gnd_net_\,
            in3 => \N__13498\,
            lcout => \receive_module.n135\,
            ltout => OPEN,
            carryin => \receive_module.n2727\,
            carryout => \receive_module.n2728\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_4_lut_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15119\,
            in2 => \_gnd_net_\,
            in3 => \N__13495\,
            lcout => \receive_module.n134\,
            ltout => OPEN,
            carryin => \receive_module.n2728\,
            carryout => \receive_module.n2729\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_5_lut_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15356\,
            in2 => \_gnd_net_\,
            in3 => \N__13492\,
            lcout => \receive_module.n133\,
            ltout => OPEN,
            carryin => \receive_module.n2729\,
            carryout => \receive_module.n2730\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_6_lut_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16763\,
            in2 => \_gnd_net_\,
            in3 => \N__13489\,
            lcout => \receive_module.n132\,
            ltout => OPEN,
            carryin => \receive_module.n2730\,
            carryout => \receive_module.n2731\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_7_lut_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13265\,
            in2 => \_gnd_net_\,
            in3 => \N__13240\,
            lcout => \receive_module.n131\,
            ltout => OPEN,
            carryin => \receive_module.n2731\,
            carryout => \receive_module.n2732\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_8_lut_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16523\,
            in2 => \_gnd_net_\,
            in3 => \N__13237\,
            lcout => \receive_module.n130\,
            ltout => OPEN,
            carryin => \receive_module.n2732\,
            carryout => \receive_module.n2733\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_9_lut_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13022\,
            in2 => \_gnd_net_\,
            in3 => \N__12991\,
            lcout => \receive_module.n129\,
            ltout => OPEN,
            carryin => \receive_module.n2733\,
            carryout => \receive_module.n2734\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_10_lut_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12776\,
            in2 => \_gnd_net_\,
            in3 => \N__12745\,
            lcout => \receive_module.n128\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \receive_module.n2735\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_11_lut_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14531\,
            in2 => \_gnd_net_\,
            in3 => \N__14497\,
            lcout => \receive_module.n127\,
            ltout => OPEN,
            carryin => \receive_module.n2735\,
            carryout => \receive_module.n2736\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_12_lut_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16160\,
            in2 => \_gnd_net_\,
            in3 => \N__14494\,
            lcout => \receive_module.n126\,
            ltout => OPEN,
            carryin => \receive_module.n2736\,
            carryout => \receive_module.n2737\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i11_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18007\,
            in2 => \_gnd_net_\,
            in3 => \N__14491\,
            lcout => \RX_ADDR_11\,
            ltout => OPEN,
            carryin => \receive_module.n2737\,
            carryout => \receive_module.n2738\,
            clk => \N__16090\,
            ce => \N__14482\,
            sr => \N__15966\
        );

    \receive_module.BRAM_ADDR__i12_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18107\,
            in2 => \_gnd_net_\,
            in3 => \N__14488\,
            lcout => \RX_ADDR_12\,
            ltout => OPEN,
            carryin => \receive_module.n2738\,
            carryout => \receive_module.n2739\,
            clk => \N__16090\,
            ce => \N__14482\,
            sr => \N__15966\
        );

    \receive_module.BRAM_ADDR__i13_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17925\,
            in2 => \_gnd_net_\,
            in3 => \N__14485\,
            lcout => \RX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16090\,
            ce => \N__14482\,
            sr => \N__15966\
        );

    \transmit_module.i1096_4_lut_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__14470\,
            in1 => \N__14423\,
            in2 => \N__14229\,
            in3 => \N__14183\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1686_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__18448\,
            in1 => \N__15813\,
            in2 => \N__13834\,
            in3 => \N__13810\,
            lcout => \line_buffer.n3119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1583_3_lut_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18449\,
            in1 => \N__13783\,
            in2 => \_gnd_net_\,
            in3 => \N__13774\,
            lcout => \line_buffer.n3027\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1701_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__15598\,
            in1 => \N__18476\,
            in2 => \N__15811\,
            in3 => \N__15583\,
            lcout => \line_buffer.n3149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i3_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__15574\,
            in1 => \N__15355\,
            in2 => \N__16480\,
            in3 => \N__17872\,
            lcout => \RX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16093\,
            ce => 'H',
            sr => \N__15967\
        );

    \receive_module.BRAM_ADDR__i2_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__17871\,
            in1 => \N__15118\,
            in2 => \N__15334\,
            in3 => \N__16466\,
            lcout => \RX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16093\,
            ce => 'H',
            sr => \N__15967\
        );

    \receive_module.BRAM_ADDR__i1_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__15091\,
            in1 => \N__14872\,
            in2 => \N__16479\,
            in3 => \N__17870\,
            lcout => \RX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16093\,
            ce => 'H',
            sr => \N__15967\
        );

    \line_buffer.n3149_bdd_4_lut_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__14848\,
            in1 => \N__15835\,
            in2 => \N__14833\,
            in3 => \N__14815\,
            lcout => OPEN,
            ltout => \line_buffer.n3152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i5_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17686\,
            in2 => \N__14806\,
            in3 => \N__15643\,
            lcout => \TX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1580_3_lut_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18472\,
            in1 => \N__14791\,
            in2 => \_gnd_net_\,
            in3 => \N__14779\,
            lcout => \line_buffer.n3024\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__15837\,
            in1 => \N__18250\,
            in2 => \N__17695\,
            in3 => \N__14764\,
            lcout => OPEN,
            ltout => \line_buffer.n3131_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i4_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__16981\,
            in1 => \N__15610\,
            in2 => \N__14752\,
            in3 => \N__17693\,
            lcout => \TX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1602_3_lut_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18490\,
            in1 => \N__17014\,
            in2 => \_gnd_net_\,
            in3 => \N__16999\,
            lcout => \line_buffer.n3046\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i4_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__16753\,
            in1 => \N__16975\,
            in2 => \N__16482\,
            in3 => \N__17873\,
            lcout => \RX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16094\,
            ce => 'H',
            sr => \N__15978\
        );

    \receive_module.BRAM_ADDR__i6_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__17874\,
            in1 => \N__16513\,
            in2 => \N__16729\,
            in3 => \N__16475\,
            lcout => \RX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16094\,
            ce => 'H',
            sr => \N__15978\
        );

    \receive_module.BRAM_ADDR__i10_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__16150\,
            in1 => \N__16492\,
            in2 => \N__16483\,
            in3 => \N__17875\,
            lcout => \RX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16097\,
            ce => 'H',
            sr => \N__15968\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_1706_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__18488\,
            in1 => \N__15904\,
            in2 => \N__15838\,
            in3 => \N__15892\,
            lcout => OPEN,
            ltout => \line_buffer.n3155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3155_bdd_4_lut_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__15874\,
            in1 => \N__15856\,
            in2 => \N__15841\,
            in3 => \N__15834\,
            lcout => \line_buffer.n3158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1601_3_lut_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15637\,
            in1 => \N__15622\,
            in2 => \_gnd_net_\,
            in3 => \N__18473\,
            lcout => \line_buffer.n3045\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1581_3_lut_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18489\,
            in1 => \N__18286\,
            in2 => \_gnd_net_\,
            in3 => \N__18271\,
            lcout => \line_buffer.n3025\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18138\,
            in1 => \N__18047\,
            in2 => \N__17974\,
            in3 => \N__17857\,
            lcout => \line_buffer.n729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__18135\,
            in1 => \N__18054\,
            in2 => \N__17973\,
            in3 => \N__17877\,
            lcout => \line_buffer.n697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__18136\,
            in1 => \N__18055\,
            in2 => \N__17975\,
            in3 => \N__17876\,
            lcout => \line_buffer.n633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
