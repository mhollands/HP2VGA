-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Oct 7 2018 23:14:28

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    TVP_VIDEO : in std_logic_vector(9 downto 0);
    ADV_B : out std_logic_vector(7 downto 0);
    ADV_G : out std_logic_vector(7 downto 0);
    ADV_R : out std_logic_vector(7 downto 0);
    DEBUG : inout std_logic_vector(7 downto 0);
    TVP_CLK : in std_logic;
    ADV_CLK : out std_logic;
    TVP_HSYNC : in std_logic;
    ADV_HSYNC : out std_logic;
    TVP_VSYNC : in std_logic;
    ADV_VSYNC : out std_logic;
    ADV_BLANK_N : out std_logic;
    LED : out std_logic;
    ADV_SYNC_N : out std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__24834\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_38\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_55\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_46\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_58\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_59\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_57\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_56\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_39\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_45\ : std_logic;
signal \line_buffer.n599\ : std_logic;
signal \line_buffer.n591\ : std_logic;
signal \line_buffer.n600\ : std_logic;
signal \line_buffer.n592\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_28\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_27\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_48\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_47\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_50\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_49\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_54\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_67\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_77\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_69\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_68\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_76\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_66\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_44\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_43\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_42\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_41\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_40\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_60\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_4\ : std_logic;
signal \line_buffer.n466\ : std_logic;
signal \line_buffer.n458\ : std_logic;
signal \line_buffer.n531\ : std_logic;
signal \line_buffer.n523\ : std_logic;
signal \TVP_VIDEO_c_4\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_29\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_30\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_32\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_31\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_33\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_37\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_36\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_35\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_34\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_81\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_82\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_80\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_51\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_70\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_71\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_79\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_78\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_72\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_75\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_53\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_52\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_74\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_73\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_61\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_65\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_64\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_63\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_62\ : std_logic;
signal \line_buffer.n3569\ : std_logic;
signal \line_buffer.n3566\ : std_logic;
signal \line_buffer.n3599_cascade_\ : std_logic;
signal \line_buffer.n595\ : std_logic;
signal \line_buffer.n587\ : std_logic;
signal \line_buffer.n3570\ : std_logic;
signal \TVP_VIDEO_c_3\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_10\ : std_logic;
signal \sync_buffer.BUFFER_0_0\ : std_logic;
signal \sync_buffer.BUFFER_1_0\ : std_logic;
signal \RX_TX_SYNC_BUFF\ : std_logic;
signal \transmit_module.video_signal_controller.n3479_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3475_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n55\ : std_logic;
signal \line_buffer.n563\ : std_logic;
signal \line_buffer.n555\ : std_logic;
signal \line_buffer.n3567\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3180\ : std_logic;
signal \transmit_module.video_signal_controller.n3181\ : std_logic;
signal \transmit_module.video_signal_controller.n3182\ : std_logic;
signal \transmit_module.video_signal_controller.n3183\ : std_logic;
signal \transmit_module.video_signal_controller.n3184\ : std_logic;
signal \transmit_module.video_signal_controller.n3185\ : std_logic;
signal \transmit_module.video_signal_controller.n3186\ : std_logic;
signal \transmit_module.video_signal_controller.n3187\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3188\ : std_logic;
signal \transmit_module.video_signal_controller.n3189\ : std_logic;
signal \transmit_module.video_signal_controller.n3190\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_1\ : std_logic;
signal \line_buffer.n536\ : std_logic;
signal \line_buffer.n528\ : std_logic;
signal \line_buffer.n3528\ : std_logic;
signal \line_buffer.n3527\ : std_logic;
signal \TX_DATA_2\ : std_logic;
signal n1816 : std_logic;
signal \line_buffer.n471\ : std_logic;
signal \line_buffer.n463\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_3\ : std_logic;
signal \RX_DATA_1\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_7\ : std_logic;
signal \DEBUG_c_6_c\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_7\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_4\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_17\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_16\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_18\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_4\ : std_logic;
signal \RX_DATA_2\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3191\ : std_logic;
signal \transmit_module.video_signal_controller.n3192\ : std_logic;
signal \transmit_module.video_signal_controller.n3193\ : std_logic;
signal \transmit_module.video_signal_controller.n3194\ : std_logic;
signal \transmit_module.video_signal_controller.n3195\ : std_logic;
signal \transmit_module.video_signal_controller.n3196\ : std_logic;
signal \transmit_module.video_signal_controller.n3197\ : std_logic;
signal \transmit_module.video_signal_controller.n3198\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3199\ : std_logic;
signal \transmit_module.video_signal_controller.n3200\ : std_logic;
signal \transmit_module.video_signal_controller.n3201\ : std_logic;
signal \transmit_module.video_signal_controller.n2395\ : std_logic;
signal \transmit_module.video_signal_controller.n7\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_0\ : std_logic;
signal \transmit_module.n3680\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_4\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_3\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_5\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_6\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_7\ : std_logic;
signal \transmit_module.video_signal_controller.n2014_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_2\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_1\ : std_logic;
signal \transmit_module.video_signal_controller.n3676\ : std_logic;
signal \transmit_module.n146\ : std_logic;
signal \transmit_module.n146_cascade_\ : std_logic;
signal n27 : std_logic;
signal \transmit_module.n107_cascade_\ : std_logic;
signal \transmit_module.n145_cascade_\ : std_logic;
signal \transmit_module.n115\ : std_logic;
signal \transmit_module.n142\ : std_logic;
signal \transmit_module.n142_cascade_\ : std_logic;
signal n23 : std_logic;
signal \transmit_module.n111\ : std_logic;
signal \transmit_module.n138\ : std_logic;
signal \transmit_module.n138_cascade_\ : std_logic;
signal \transmit_module.n107\ : std_logic;
signal n19 : std_logic;
signal \transmit_module.n139\ : std_logic;
signal \transmit_module.n108\ : std_logic;
signal \transmit_module.n139_cascade_\ : std_logic;
signal n20 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_10\ : std_logic;
signal \transmit_module.n145\ : std_logic;
signal n26 : std_logic;
signal \transmit_module.n114\ : std_logic;
signal \transmit_module.n144\ : std_logic;
signal \transmit_module.n144_cascade_\ : std_logic;
signal n25 : std_logic;
signal \transmit_module.n113\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_2\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_3\ : std_logic;
signal \line_buffer.n568\ : std_logic;
signal \line_buffer.n560\ : std_logic;
signal \line_buffer.n3530\ : std_logic;
signal \line_buffer.n3531_cascade_\ : std_logic;
signal \line_buffer.n3617\ : std_logic;
signal \TX_DATA_7\ : std_logic;
signal \ADV_B_c\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_26\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_25\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_19\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_20\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_21\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_22\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_24\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_23\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.video_signal_controller.n6_adj_622_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_3\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_4\ : std_logic;
signal \transmit_module.video_signal_controller.n3482_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_6\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_5\ : std_logic;
signal \transmit_module.video_signal_controller.n6_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2016\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_8\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_7\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_2\ : std_logic;
signal \transmit_module.video_signal_controller.n3517\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_1\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_0\ : std_logic;
signal \transmit_module.video_signal_controller.n2955\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_8\ : std_logic;
signal \transmit_module.video_signal_controller.n3363\ : std_logic;
signal \transmit_module.video_signal_controller.n2014\ : std_logic;
signal \transmit_module.video_signal_controller.n2972_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2047\ : std_logic;
signal \transmit_module.VGA_VISIBLE_Y\ : std_logic;
signal \ADV_HSYNC_c\ : std_logic;
signal \transmit_module.old_VGA_HS\ : std_logic;
signal \transmit_module.n3675_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n6_adj_623_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_VISIBLE_N_588\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_11\ : std_logic;
signal \transmit_module.video_signal_controller.n7_adj_624_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3004\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_10\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_9\ : std_logic;
signal \transmit_module.video_signal_controller.n3014\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \transmit_module.n131\ : std_logic;
signal \transmit_module.n3159\ : std_logic;
signal \transmit_module.TX_ADDR_2\ : std_logic;
signal \transmit_module.n130\ : std_logic;
signal \transmit_module.n3160\ : std_logic;
signal \transmit_module.TX_ADDR_3\ : std_logic;
signal \transmit_module.n129\ : std_logic;
signal \transmit_module.n3161\ : std_logic;
signal \transmit_module.n3162\ : std_logic;
signal \transmit_module.n127\ : std_logic;
signal \transmit_module.n3163\ : std_logic;
signal \transmit_module.n3164\ : std_logic;
signal \transmit_module.n3165\ : std_logic;
signal \transmit_module.n3166\ : std_logic;
signal \transmit_module.n124\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \transmit_module.n123\ : std_logic;
signal \transmit_module.n3167\ : std_logic;
signal \transmit_module.n3168\ : std_logic;
signal \transmit_module.n3169\ : std_logic;
signal \transmit_module.n3170\ : std_logic;
signal \transmit_module.n3171\ : std_logic;
signal \transmit_module.TX_ADDR_9\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_9\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_0\ : std_logic;
signal \transmit_module.TX_ADDR_1\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_1\ : std_logic;
signal \transmit_module.TX_ADDR_8\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_8\ : std_logic;
signal \transmit_module.TX_ADDR_5\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_5\ : std_logic;
signal \transmit_module.TX_ADDR_10\ : std_logic;
signal \transmit_module.n122\ : std_logic;
signal n22 : std_logic;
signal \transmit_module.n112_cascade_\ : std_logic;
signal n24 : std_logic;
signal \transmit_module.n125\ : std_logic;
signal \transmit_module.n140\ : std_logic;
signal \transmit_module.n140_cascade_\ : std_logic;
signal \transmit_module.n109\ : std_logic;
signal n21 : std_logic;
signal \transmit_module.n106\ : std_logic;
signal \transmit_module.n137\ : std_logic;
signal n18 : std_logic;
signal \TVP_VIDEO_c_5\ : std_logic;
signal \DEBUG_c_1_c\ : std_logic;
signal \tvp_vs_buffer.BUFFER_0_0\ : std_logic;
signal \tvp_vs_buffer.BUFFER_1_0\ : std_logic;
signal \RX_DATA_5\ : std_logic;
signal \receive_module.sync_wd.n6_cascade_\ : std_logic;
signal \receive_module.sync_wd.n4_cascade_\ : std_logic;
signal \receive_module.sync_wd.old_visible\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \receive_module.rx_counter.n3207\ : std_logic;
signal \receive_module.rx_counter.n3208\ : std_logic;
signal \receive_module.rx_counter.n3209\ : std_logic;
signal \receive_module.rx_counter.n3210\ : std_logic;
signal \receive_module.rx_counter.n3211\ : std_logic;
signal \receive_module.rx_counter.n3212\ : std_logic;
signal \receive_module.rx_counter.n3213\ : std_logic;
signal \receive_module.rx_counter.n3214\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \receive_module.rx_counter.n3215\ : std_logic;
signal \tvp_vs_buffer.BUFFER_2_0\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_11\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_10\ : std_logic;
signal \transmit_module.video_signal_controller.n3461\ : std_logic;
signal \transmit_module.video_signal_controller.n3375\ : std_logic;
signal \transmit_module.video_signal_controller.n3673_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_9\ : std_logic;
signal \transmit_module.video_signal_controller.n3379\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.n126\ : std_logic;
signal \transmit_module.n141\ : std_logic;
signal \transmit_module.n141_cascade_\ : std_logic;
signal \transmit_module.n110\ : std_logic;
signal \transmit_module.n132\ : std_logic;
signal \transmit_module.n147_cascade_\ : std_logic;
signal n28 : std_logic;
signal \transmit_module.VGA_VISIBLE\ : std_logic;
signal \transmit_module.n128\ : std_logic;
signal \transmit_module.n143\ : std_logic;
signal \transmit_module.n112\ : std_logic;
signal \transmit_module.n143_cascade_\ : std_logic;
signal \transmit_module.n116\ : std_logic;
signal \transmit_module.n147\ : std_logic;
signal \transmit_module.TX_ADDR_0\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \receive_module.n3146\ : std_logic;
signal \receive_module.n3147\ : std_logic;
signal \receive_module.n3148\ : std_logic;
signal \receive_module.n3149\ : std_logic;
signal \receive_module.n3150\ : std_logic;
signal \receive_module.n3151\ : std_logic;
signal \receive_module.n3152\ : std_logic;
signal \receive_module.n3153\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \receive_module.n3154\ : std_logic;
signal \receive_module.n3155\ : std_logic;
signal \receive_module.n3156\ : std_logic;
signal \receive_module.n3157\ : std_logic;
signal \receive_module.n3158\ : std_logic;
signal \transmit_module.TX_ADDR_4\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_4\ : std_logic;
signal \transmit_module.TX_ADDR_7\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_7\ : std_logic;
signal \transmit_module.TX_ADDR_6\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_6\ : std_logic;
signal \transmit_module.n2310\ : std_logic;
signal \receive_module.n136\ : std_logic;
signal \RX_ADDR_1\ : std_logic;
signal \receive_module.n127\ : std_logic;
signal \RX_ADDR_10\ : std_logic;
signal \receive_module.n137\ : std_logic;
signal \RX_ADDR_0\ : std_logic;
signal n1818 : std_logic;
signal \receive_module.n135\ : std_logic;
signal \RX_ADDR_2\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_5\ : std_logic;
signal \receive_module.rx_counter.n3452_cascade_\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_5\ : std_logic;
signal \RX_DATA_3\ : std_logic;
signal \receive_module.rx_counter.n10\ : std_logic;
signal \receive_module.rx_counter.n14_cascade_\ : std_logic;
signal \RX_TX_SYNC\ : std_logic;
signal \receive_module.rx_counter.n4\ : std_logic;
signal \receive_module.rx_counter.n5_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3450\ : std_logic;
signal \receive_module.rx_counter.n3677\ : std_logic;
signal \receive_module.rx_counter.n3\ : std_logic;
signal \receive_module.rx_counter.X_1\ : std_logic;
signal \receive_module.rx_counter.X_2\ : std_logic;
signal \receive_module.rx_counter.X_0\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \receive_module.rx_counter.n3202\ : std_logic;
signal \receive_module.rx_counter.n3203\ : std_logic;
signal \receive_module.rx_counter.n3204\ : std_logic;
signal \receive_module.rx_counter.n3205\ : std_logic;
signal \receive_module.rx_counter.n3206\ : std_logic;
signal \receive_module.rx_counter.n6\ : std_logic;
signal \receive_module.rx_counter.n7\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_5\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_1\ : std_logic;
signal \receive_module.rx_counter.X_3\ : std_logic;
signal \receive_module.rx_counter.X_5\ : std_logic;
signal \receive_module.rx_counter.X_4\ : std_logic;
signal \receive_module.rx_counter.n3222\ : std_logic;
signal \receive_module.rx_counter.X_7\ : std_logic;
signal \receive_module.rx_counter.n3455_cascade_\ : std_logic;
signal \receive_module.rx_counter.X_6\ : std_logic;
signal \receive_module.rx_counter.X_8\ : std_logic;
signal \receive_module.rx_counter.X_9\ : std_logic;
signal \receive_module.rx_counter.n39_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3426\ : std_logic;
signal \receive_module.rx_counter.n3478\ : std_logic;
signal \receive_module.rx_counter.n54_cascade_\ : std_logic;
signal \receive_module.rx_counter.n4_adj_612\ : std_logic;
signal \line_buffer.n473\ : std_logic;
signal \line_buffer.n570\ : std_logic;
signal \line_buffer.n571\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_11\ : std_logic;
signal \transmit_module.n121\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_13\ : std_logic;
signal \transmit_module.n119\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_12\ : std_logic;
signal \transmit_module.n3675\ : std_logic;
signal \transmit_module.n120\ : std_logic;
signal \transmit_module.n2070\ : std_logic;
signal \receive_module.n3671\ : std_logic;
signal \line_buffer.n603\ : std_logic;
signal \line_buffer.n539\ : std_logic;
signal \line_buffer.n474\ : std_logic;
signal \receive_module.n128\ : std_logic;
signal \RX_ADDR_9\ : std_logic;
signal \receive_module.n134\ : std_logic;
signal \RX_ADDR_3\ : std_logic;
signal \receive_module.n133\ : std_logic;
signal \RX_ADDR_4\ : std_logic;
signal \receive_module.n129\ : std_logic;
signal \RX_ADDR_8\ : std_logic;
signal \receive_module.n131\ : std_logic;
signal \RX_ADDR_6\ : std_logic;
signal \receive_module.n130\ : std_logic;
signal \RX_ADDR_7\ : std_logic;
signal \line_buffer.n564\ : std_logic;
signal \line_buffer.n556\ : std_logic;
signal \line_buffer.n532\ : std_logic;
signal \line_buffer.n524\ : std_logic;
signal \line_buffer.n467\ : std_logic;
signal \line_buffer.n459\ : std_logic;
signal \line_buffer.n3587\ : std_logic;
signal \line_buffer.n3590_cascade_\ : std_logic;
signal \line_buffer.n3626\ : std_logic;
signal \TX_DATA_3\ : std_logic;
signal n1815 : std_logic;
signal \line_buffer.n602\ : std_logic;
signal \GB_BUFFER_DEBUG_c_3_c_THRU_CO\ : std_logic;
signal \DEBUG_c_0\ : std_logic;
signal \LED_c\ : std_logic;
signal \TVP_VIDEO_c_2\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_2\ : std_logic;
signal \receive_module.rx_counter.Y_0\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \receive_module.rx_counter.Y_1\ : std_logic;
signal \receive_module.rx_counter.n3172\ : std_logic;
signal \receive_module.rx_counter.Y_2\ : std_logic;
signal \receive_module.rx_counter.n3173\ : std_logic;
signal \receive_module.rx_counter.Y_3\ : std_logic;
signal \receive_module.rx_counter.n3174\ : std_logic;
signal \receive_module.rx_counter.Y_4\ : std_logic;
signal \receive_module.rx_counter.n3175\ : std_logic;
signal \receive_module.rx_counter.Y_5\ : std_logic;
signal \receive_module.rx_counter.n3176\ : std_logic;
signal \receive_module.rx_counter.Y_6\ : std_logic;
signal \receive_module.rx_counter.n3177\ : std_logic;
signal \receive_module.rx_counter.Y_7\ : std_logic;
signal \receive_module.rx_counter.n3178\ : std_logic;
signal \receive_module.rx_counter.n3179\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \receive_module.rx_counter.Y_8\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_2\ : std_logic;
signal \RX_DATA_0\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_4\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_2\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_0\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_3\ : std_logic;
signal \receive_module.rx_counter.n7_adj_619_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3519\ : std_logic;
signal \receive_module.rx_counter.old_VS\ : std_logic;
signal \receive_module.rx_counter.n11_cascade_\ : std_logic;
signal \receive_module.rx_counter.n2547\ : std_logic;
signal \receive_module.rx_counter.n11\ : std_logic;
signal \PULSE_1HZ\ : std_logic;
signal \receive_module.rx_counter.n3672\ : std_logic;
signal \RX_ADDR_12\ : std_logic;
signal \RX_ADDR_13\ : std_logic;
signal \RX_ADDR_11\ : std_logic;
signal \line_buffer.n538\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.n2084\ : std_logic;
signal \DEBUG_c_7_c\ : std_logic;
signal \RX_DATA_6\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_8\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_8\ : std_logic;
signal \line_buffer.n598\ : std_logic;
signal \line_buffer.n590\ : std_logic;
signal \line_buffer.n526\ : std_logic;
signal \line_buffer.n534\ : std_logic;
signal \line_buffer.n3593_cascade_\ : std_logic;
signal \line_buffer.n554\ : std_logic;
signal \line_buffer.n562\ : std_logic;
signal \receive_module.n132\ : std_logic;
signal \DEBUG_c_4\ : std_logic;
signal \RX_ADDR_5\ : std_logic;
signal \receive_module.n3674\ : std_logic;
signal \line_buffer.n596\ : std_logic;
signal \line_buffer.n588\ : std_logic;
signal \line_buffer.n3623\ : std_logic;
signal \DEBUG_c_2_c\ : std_logic;
signal \tvp_hs_buffer.BUFFER_0_0\ : std_logic;
signal \tvp_hs_buffer.BUFFER_1_0\ : std_logic;
signal \TVP_VSYNC_buff\ : std_logic;
signal \receive_module.rx_counter.n2078\ : std_logic;
signal \TVP_HSYNC_buff\ : std_logic;
signal \receive_module.rx_counter.old_HS\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_98\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_89\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_92\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_91\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_90\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_99\ : std_logic;
signal \transmit_module.n3679\ : std_logic;
signal \line_buffer.n566\ : std_logic;
signal \line_buffer.n558\ : std_logic;
signal \line_buffer.n465\ : std_logic;
signal \line_buffer.n457\ : std_logic;
signal \line_buffer.n3629\ : std_logic;
signal \line_buffer.n561\ : std_logic;
signal \line_buffer.n553\ : std_logic;
signal \line_buffer.n456\ : std_logic;
signal \line_buffer.n464\ : std_logic;
signal \line_buffer.n3635_cascade_\ : std_logic;
signal \line_buffer.n469\ : std_logic;
signal \line_buffer.n461\ : std_logic;
signal \line_buffer.n3653\ : std_logic;
signal \line_buffer.n3656_cascade_\ : std_logic;
signal \line_buffer.n3596\ : std_logic;
signal \line_buffer.n3638\ : std_logic;
signal \TX_DATA_0\ : std_logic;
signal \line_buffer.n530\ : std_logic;
signal \line_buffer.n522\ : std_logic;
signal \line_buffer.n3632\ : std_logic;
signal \line_buffer.n3650_cascade_\ : std_logic;
signal \line_buffer.n594\ : std_logic;
signal \line_buffer.n586\ : std_logic;
signal \line_buffer.n3647\ : std_logic;
signal \line_buffer.n521\ : std_logic;
signal \line_buffer.n529\ : std_logic;
signal \line_buffer.n3644\ : std_logic;
signal \TX_DATA_5\ : std_logic;
signal n1813 : std_logic;
signal \TX_DATA_1\ : std_logic;
signal n1817 : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_97\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_96\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_95\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_94\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_93\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_83\ : std_logic;
signal \line_buffer.n593\ : std_logic;
signal \line_buffer.n585\ : std_logic;
signal \line_buffer.n3641\ : std_logic;
signal \line_buffer.n533\ : std_logic;
signal \line_buffer.n525\ : std_logic;
signal \RX_DATA_7\ : std_logic;
signal \line_buffer.n565\ : std_logic;
signal \line_buffer.n557\ : std_logic;
signal \line_buffer.n3533\ : std_logic;
signal \line_buffer.n3549\ : std_logic;
signal \line_buffer.n3611_cascade_\ : std_logic;
signal \RX_DATA_4\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_6\ : std_logic;
signal \DEBUG_c_5_c\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_6\ : std_logic;
signal \line_buffer.n468\ : std_logic;
signal \line_buffer.n460\ : std_logic;
signal \line_buffer.n3548\ : std_logic;
signal \line_buffer.n567\ : std_logic;
signal \line_buffer.n559\ : std_logic;
signal \TX_ADDR_12\ : std_logic;
signal \line_buffer.n3540\ : std_logic;
signal \line_buffer.n3573\ : std_logic;
signal \TX_ADDR_13\ : std_logic;
signal \line_buffer.n3605\ : std_logic;
signal \TX_DATA_4\ : std_logic;
signal n1814 : std_logic;
signal \TX_DATA_6\ : std_logic;
signal n1812 : std_logic;
signal \transmit_module.n2385\ : std_logic;
signal \line_buffer.n470\ : std_logic;
signal \line_buffer.n462\ : std_logic;
signal \line_buffer.n3572\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \TVP_VIDEO_c_9\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_9\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_9\ : std_logic;
signal \DEBUG_c_3_c\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_88\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_84\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_85\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_87\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_86\ : std_logic;
signal \ADV_CLK_c\ : std_logic;
signal \transmit_module.n2206\ : std_logic;
signal \ADV_VSYNC_c\ : std_logic;
signal \line_buffer.n589\ : std_logic;
signal \line_buffer.n597\ : std_logic;
signal \line_buffer.n3534\ : std_logic;
signal \TX_ADDR_11\ : std_logic;
signal \line_buffer.n535\ : std_logic;
signal \line_buffer.n527\ : std_logic;
signal \line_buffer.n3539\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \TVP_CLK_wire\ : std_logic;
signal \ADV_CLK_wire\ : std_logic;
signal \TVP_HSYNC_wire\ : std_logic;
signal \TVP_VIDEO_wire\ : std_logic_vector(9 downto 0);
signal \ADV_G_wire\ : std_logic_vector(7 downto 0);
signal \ADV_R_wire\ : std_logic_vector(7 downto 0);
signal \ADV_B_wire\ : std_logic_vector(7 downto 0);
signal \ADV_SYNC_N_wire\ : std_logic;
signal \ADV_BLANK_N_wire\ : std_logic;
signal \TVP_VSYNC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \ADV_HSYNC_wire\ : std_logic;
signal \ADV_VSYNC_wire\ : std_logic;
signal \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \line_buffer.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \TVP_CLK_wire\ <= TVP_CLK;
    ADV_CLK <= \ADV_CLK_wire\;
    \TVP_HSYNC_wire\ <= TVP_HSYNC;
    \TVP_VIDEO_wire\ <= TVP_VIDEO;
    ADV_G <= \ADV_G_wire\;
    ADV_R <= \ADV_R_wire\;
    ADV_B <= \ADV_B_wire\;
    ADV_SYNC_N <= \ADV_SYNC_N_wire\;
    ADV_BLANK_N <= \ADV_BLANK_N_wire\;
    \TVP_VSYNC_wire\ <= TVP_VSYNC;
    LED <= \LED_wire\;
    ADV_HSYNC <= \ADV_HSYNC_wire\;
    ADV_VSYNC <= \ADV_VSYNC_wire\;
    \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.n471\ <= \line_buffer.mem2_physical_RDATA_wire\(11);
    \line_buffer.n470\ <= \line_buffer.mem2_physical_RDATA_wire\(3);
    \line_buffer.mem2_physical_RADDR_wire\ <= \N__12593\&\N__10277\&\N__11276\&\N__12845\&\N__13319\&\N__10532\&\N__13100\&\N__10796\&\N__11048\&\N__10028\&\N__14129\;
    \line_buffer.mem2_physical_WADDR_wire\ <= \N__14939\&\N__17918\&\N__17168\&\N__16664\&\N__16916\&\N__19397\&\N__17420\&\N__17669\&\N__14402\&\N__15176\&\N__14693\;
    \line_buffer.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21057\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19914\&'0'&'0'&'0';
    \line_buffer.n558\ <= \line_buffer.mem14_physical_RDATA_wire\(11);
    \line_buffer.n557\ <= \line_buffer.mem14_physical_RDATA_wire\(3);
    \line_buffer.mem14_physical_RADDR_wire\ <= \N__12665\&\N__10349\&\N__11348\&\N__12917\&\N__13391\&\N__10604\&\N__13172\&\N__10868\&\N__11120\&\N__10100\&\N__14201\;
    \line_buffer.mem14_physical_WADDR_wire\ <= \N__15011\&\N__17990\&\N__17240\&\N__16736\&\N__16988\&\N__19469\&\N__17492\&\N__17741\&\N__14474\&\N__15248\&\N__14765\;
    \line_buffer.mem14_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem14_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__13572\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21727\&'0'&'0'&'0';
    \line_buffer.n568\ <= \line_buffer.mem5_physical_RDATA_wire\(11);
    \line_buffer.n567\ <= \line_buffer.mem5_physical_RDATA_wire\(3);
    \line_buffer.mem5_physical_RADDR_wire\ <= \N__12596\&\N__10274\&\N__11297\&\N__12848\&\N__13328\&\N__10523\&\N__13103\&\N__10787\&\N__11039\&\N__10043\&\N__14126\;
    \line_buffer.mem5_physical_WADDR_wire\ <= \N__14948\&\N__17927\&\N__17177\&\N__16679\&\N__16931\&\N__19412\&\N__17429\&\N__17672\&\N__14405\&\N__15185\&\N__14702\;
    \line_buffer.mem5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21051\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19909\&'0'&'0'&'0';
    \line_buffer.n526\ <= \line_buffer.mem11_physical_RDATA_wire\(11);
    \line_buffer.n525\ <= \line_buffer.mem11_physical_RDATA_wire\(3);
    \line_buffer.mem11_physical_RADDR_wire\ <= \N__12701\&\N__10385\&\N__11384\&\N__12953\&\N__13427\&\N__10640\&\N__13208\&\N__10904\&\N__11156\&\N__10136\&\N__14237\;
    \line_buffer.mem11_physical_WADDR_wire\ <= \N__15047\&\N__18026\&\N__17276\&\N__16772\&\N__17024\&\N__19505\&\N__17528\&\N__17777\&\N__14510\&\N__15284\&\N__14801\;
    \line_buffer.mem11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem11_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__13571\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21738\&'0'&'0'&'0';
    \line_buffer.n588\ <= \line_buffer.mem21_physical_RDATA_wire\(11);
    \line_buffer.n587\ <= \line_buffer.mem21_physical_RDATA_wire\(3);
    \line_buffer.mem21_physical_RADDR_wire\ <= \N__12569\&\N__10253\&\N__11252\&\N__12821\&\N__13295\&\N__10508\&\N__13076\&\N__10772\&\N__11024\&\N__10004\&\N__14105\;
    \line_buffer.mem21_physical_WADDR_wire\ <= \N__14915\&\N__17894\&\N__17144\&\N__16640\&\N__16892\&\N__19373\&\N__17396\&\N__17645\&\N__14378\&\N__15152\&\N__14669\;
    \line_buffer.mem21_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem21_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__15653\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9524\&'0'&'0'&'0';
    \line_buffer.n524\ <= \line_buffer.mem12_physical_RDATA_wire\(11);
    \line_buffer.n523\ <= \line_buffer.mem12_physical_RDATA_wire\(3);
    \line_buffer.mem12_physical_RADDR_wire\ <= \N__12689\&\N__10373\&\N__11372\&\N__12941\&\N__13415\&\N__10628\&\N__13196\&\N__10892\&\N__11144\&\N__10124\&\N__14225\;
    \line_buffer.mem12_physical_WADDR_wire\ <= \N__15035\&\N__18014\&\N__17264\&\N__16760\&\N__17012\&\N__19493\&\N__17516\&\N__17765\&\N__14498\&\N__15272\&\N__14789\;
    \line_buffer.mem12_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem12_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__15593\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9513\&'0'&'0'&'0';
    \line_buffer.n532\ <= \line_buffer.mem24_physical_RDATA_wire\(11);
    \line_buffer.n531\ <= \line_buffer.mem24_physical_RDATA_wire\(3);
    \line_buffer.mem24_physical_RADDR_wire\ <= \N__12716\&\N__10394\&\N__11417\&\N__12968\&\N__13448\&\N__10643\&\N__13223\&\N__10907\&\N__11159\&\N__10163\&\N__14246\;
    \line_buffer.mem24_physical_WADDR_wire\ <= \N__15068\&\N__18047\&\N__17297\&\N__16799\&\N__17051\&\N__19532\&\N__17549\&\N__17792\&\N__14525\&\N__15305\&\N__14822\;
    \line_buffer.mem24_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem24_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__15635\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9519\&'0'&'0'&'0';
    \line_buffer.n560\ <= \line_buffer.mem1_physical_RDATA_wire\(11);
    \line_buffer.n559\ <= \line_buffer.mem1_physical_RDATA_wire\(3);
    \line_buffer.mem1_physical_RADDR_wire\ <= \N__12725\&\N__10407\&\N__11408\&\N__12977\&\N__13451\&\N__10659\&\N__13232\&\N__10923\&\N__11175\&\N__10160\&\N__14259\;
    \line_buffer.mem1_physical_WADDR_wire\ <= \N__15071\&\N__18050\&\N__17300\&\N__16796\&\N__17048\&\N__19529\&\N__17552\&\N__17801\&\N__14534\&\N__15308\&\N__14825\;
    \line_buffer.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21029\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19922\&'0'&'0'&'0';
    \line_buffer.n556\ <= \line_buffer.mem15_physical_RDATA_wire\(11);
    \line_buffer.n555\ <= \line_buffer.mem15_physical_RDATA_wire\(3);
    \line_buffer.mem15_physical_RADDR_wire\ <= \N__12653\&\N__10337\&\N__11336\&\N__12905\&\N__13379\&\N__10592\&\N__13160\&\N__10856\&\N__11108\&\N__10088\&\N__14189\;
    \line_buffer.mem15_physical_WADDR_wire\ <= \N__14999\&\N__17978\&\N__17228\&\N__16724\&\N__16976\&\N__19457\&\N__17480\&\N__17729\&\N__14462\&\N__15236\&\N__14753\;
    \line_buffer.mem15_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem15_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__15640\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9514\&'0'&'0'&'0';
    \line_buffer.n564\ <= \line_buffer.mem27_physical_RDATA_wire\(11);
    \line_buffer.n563\ <= \line_buffer.mem27_physical_RDATA_wire\(3);
    \line_buffer.mem27_physical_RADDR_wire\ <= \N__12680\&\N__10358\&\N__11381\&\N__12932\&\N__13412\&\N__10607\&\N__13187\&\N__10871\&\N__11123\&\N__10127\&\N__14210\;
    \line_buffer.mem27_physical_WADDR_wire\ <= \N__15032\&\N__18011\&\N__17261\&\N__16763\&\N__17015\&\N__19496\&\N__17513\&\N__17756\&\N__14489\&\N__15269\&\N__14786\;
    \line_buffer.mem27_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem27_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__15586\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9503\&'0'&'0'&'0';
    \line_buffer.n536\ <= \line_buffer.mem4_physical_RDATA_wire\(11);
    \line_buffer.n535\ <= \line_buffer.mem4_physical_RDATA_wire\(3);
    \line_buffer.mem4_physical_RADDR_wire\ <= \N__12608\&\N__10286\&\N__11309\&\N__12860\&\N__13340\&\N__10535\&\N__13115\&\N__10799\&\N__11051\&\N__10055\&\N__14138\;
    \line_buffer.mem4_physical_WADDR_wire\ <= \N__14960\&\N__17939\&\N__17189\&\N__16691\&\N__16943\&\N__19424\&\N__17441\&\N__17684\&\N__14417\&\N__15197\&\N__14714\;
    \line_buffer.mem4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21050\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19891\&'0'&'0'&'0';
    \line_buffer.n554\ <= \line_buffer.mem16_physical_RDATA_wire\(11);
    \line_buffer.n553\ <= \line_buffer.mem16_physical_RDATA_wire\(3);
    \line_buffer.mem16_physical_RADDR_wire\ <= \N__12641\&\N__10325\&\N__11324\&\N__12893\&\N__13367\&\N__10580\&\N__13148\&\N__10844\&\N__11096\&\N__10076\&\N__14177\;
    \line_buffer.mem16_physical_WADDR_wire\ <= \N__14987\&\N__17966\&\N__17216\&\N__16712\&\N__16964\&\N__19445\&\N__17468\&\N__17717\&\N__14450\&\N__15224\&\N__14741\;
    \line_buffer.mem16_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem16_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9312\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19134\&'0'&'0'&'0';
    \line_buffer.n596\ <= \line_buffer.mem30_physical_RDATA_wire\(11);
    \line_buffer.n595\ <= \line_buffer.mem30_physical_RDATA_wire\(3);
    \line_buffer.mem30_physical_RADDR_wire\ <= \N__12632\&\N__10310\&\N__11333\&\N__12884\&\N__13364\&\N__10559\&\N__13139\&\N__10823\&\N__11075\&\N__10079\&\N__14162\;
    \line_buffer.mem30_physical_WADDR_wire\ <= \N__14984\&\N__17963\&\N__17213\&\N__16715\&\N__16967\&\N__19448\&\N__17465\&\N__17708\&\N__14441\&\N__15221\&\N__14738\;
    \line_buffer.mem30_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem30_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__15636\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9520\&'0'&'0'&'0';
    \line_buffer.n463\ <= \line_buffer.mem7_physical_RDATA_wire\(11);
    \line_buffer.n462\ <= \line_buffer.mem7_physical_RDATA_wire\(3);
    \line_buffer.mem7_physical_RADDR_wire\ <= \N__12572\&\N__10250\&\N__11273\&\N__12824\&\N__13304\&\N__10499\&\N__13079\&\N__10763\&\N__11015\&\N__10019\&\N__14102\;
    \line_buffer.mem7_physical_WADDR_wire\ <= \N__14924\&\N__17903\&\N__17153\&\N__16655\&\N__16907\&\N__19388\&\N__17405\&\N__17648\&\N__14381\&\N__15161\&\N__14678\;
    \line_buffer.mem7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem7_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21053\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19921\&'0'&'0'&'0';
    \line_buffer.n590\ <= \line_buffer.mem20_physical_RDATA_wire\(11);
    \line_buffer.n589\ <= \line_buffer.mem20_physical_RDATA_wire\(3);
    \line_buffer.mem20_physical_RADDR_wire\ <= \N__12581\&\N__10265\&\N__11264\&\N__12833\&\N__13307\&\N__10520\&\N__13088\&\N__10784\&\N__11036\&\N__10016\&\N__14117\;
    \line_buffer.mem20_physical_WADDR_wire\ <= \N__14927\&\N__17906\&\N__17156\&\N__16652\&\N__16904\&\N__19385\&\N__17408\&\N__17657\&\N__14390\&\N__15164\&\N__14681\;
    \line_buffer.mem20_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem20_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__13580\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21737\&'0'&'0'&'0';
    \line_buffer.n522\ <= \line_buffer.mem13_physical_RDATA_wire\(11);
    \line_buffer.n521\ <= \line_buffer.mem13_physical_RDATA_wire\(3);
    \line_buffer.mem13_physical_RADDR_wire\ <= \N__12677\&\N__10361\&\N__11360\&\N__12929\&\N__13403\&\N__10616\&\N__13184\&\N__10880\&\N__11132\&\N__10112\&\N__14213\;
    \line_buffer.mem13_physical_WADDR_wire\ <= \N__15023\&\N__18002\&\N__17252\&\N__16748\&\N__17000\&\N__19481\&\N__17504\&\N__17753\&\N__14486\&\N__15260\&\N__14777\;
    \line_buffer.mem13_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem13_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9311\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19119\&'0'&'0'&'0';
    \line_buffer.n465\ <= \line_buffer.mem19_physical_RDATA_wire\(11);
    \line_buffer.n464\ <= \line_buffer.mem19_physical_RDATA_wire\(3);
    \line_buffer.mem19_physical_RADDR_wire\ <= \N__12605\&\N__10289\&\N__11288\&\N__12857\&\N__13331\&\N__10544\&\N__13112\&\N__10808\&\N__11060\&\N__10040\&\N__14141\;
    \line_buffer.mem19_physical_WADDR_wire\ <= \N__14951\&\N__17930\&\N__17180\&\N__16676\&\N__16928\&\N__19409\&\N__17432\&\N__17681\&\N__14414\&\N__15188\&\N__14705\;
    \line_buffer.mem19_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem19_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9331\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19148\&'0'&'0'&'0';
    \line_buffer.n534\ <= \line_buffer.mem23_physical_RDATA_wire\(11);
    \line_buffer.n533\ <= \line_buffer.mem23_physical_RDATA_wire\(3);
    \line_buffer.mem23_physical_RADDR_wire\ <= \N__12728\&\N__10406\&\N__11424\&\N__12980\&\N__13460\&\N__10655\&\N__13235\&\N__10919\&\N__11171\&\N__10173\&\N__14258\;
    \line_buffer.mem23_physical_WADDR_wire\ <= \N__15080\&\N__18059\&\N__17309\&\N__16809\&\N__17061\&\N__19542\&\N__17561\&\N__17804\&\N__14537\&\N__15317\&\N__14834\;
    \line_buffer.mem23_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem23_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__13553\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21726\&'0'&'0'&'0';
    \line_buffer.n528\ <= \line_buffer.mem0_physical_RDATA_wire\(11);
    \line_buffer.n527\ <= \line_buffer.mem0_physical_RDATA_wire\(3);
    \line_buffer.mem0_physical_RADDR_wire\ <= \N__12732\&\N__10413\&\N__11420\&\N__12984\&\N__13461\&\N__10665\&\N__13239\&\N__10929\&\N__11181\&\N__10172\&\N__14265\;
    \line_buffer.mem0_physical_WADDR_wire\ <= \N__15081\&\N__18060\&\N__17310\&\N__16808\&\N__17060\&\N__19541\&\N__17562\&\N__17808\&\N__14541\&\N__15318\&\N__14835\;
    \line_buffer.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21049\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19926\&'0'&'0'&'0';
    \line_buffer.n566\ <= \line_buffer.mem26_physical_RDATA_wire\(11);
    \line_buffer.n565\ <= \line_buffer.mem26_physical_RDATA_wire\(3);
    \line_buffer.mem26_physical_RADDR_wire\ <= \N__12692\&\N__10370\&\N__11393\&\N__12944\&\N__13424\&\N__10619\&\N__13199\&\N__10883\&\N__11135\&\N__10139\&\N__14222\;
    \line_buffer.mem26_physical_WADDR_wire\ <= \N__15044\&\N__18023\&\N__17273\&\N__16775\&\N__17027\&\N__19508\&\N__17525\&\N__17768\&\N__14501\&\N__15281\&\N__14798\;
    \line_buffer.mem26_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem26_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__13570\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21724\&'0'&'0'&'0';
    \line_buffer.n592\ <= \line_buffer.mem3_physical_RDATA_wire\(11);
    \line_buffer.n591\ <= \line_buffer.mem3_physical_RDATA_wire\(3);
    \line_buffer.mem3_physical_RADDR_wire\ <= \N__12644\&\N__10322\&\N__11345\&\N__12896\&\N__13376\&\N__10571\&\N__13151\&\N__10835\&\N__11087\&\N__10091\&\N__14174\;
    \line_buffer.mem3_physical_WADDR_wire\ <= \N__14996\&\N__17975\&\N__17225\&\N__16727\&\N__16979\&\N__19460\&\N__17477\&\N__17720\&\N__14453\&\N__15233\&\N__14750\;
    \line_buffer.mem3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21033\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19874\&'0'&'0'&'0';
    \line_buffer.n469\ <= \line_buffer.mem17_physical_RDATA_wire\(11);
    \line_buffer.n468\ <= \line_buffer.mem17_physical_RDATA_wire\(3);
    \line_buffer.mem17_physical_RADDR_wire\ <= \N__12629\&\N__10313\&\N__11312\&\N__12881\&\N__13355\&\N__10568\&\N__13136\&\N__10832\&\N__11084\&\N__10064\&\N__14165\;
    \line_buffer.mem17_physical_WADDR_wire\ <= \N__14975\&\N__17954\&\N__17204\&\N__16700\&\N__16952\&\N__19433\&\N__17456\&\N__17705\&\N__14438\&\N__15212\&\N__14729\;
    \line_buffer.mem17_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem17_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__13573\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21714\&'0'&'0'&'0';
    \line_buffer.n594\ <= \line_buffer.mem31_physical_RDATA_wire\(11);
    \line_buffer.n593\ <= \line_buffer.mem31_physical_RDATA_wire\(3);
    \line_buffer.mem31_physical_RADDR_wire\ <= \N__12620\&\N__10298\&\N__11321\&\N__12872\&\N__13352\&\N__10547\&\N__13127\&\N__10811\&\N__11063\&\N__10067\&\N__14150\;
    \line_buffer.mem31_physical_WADDR_wire\ <= \N__14972\&\N__17951\&\N__17201\&\N__16703\&\N__16955\&\N__19436\&\N__17453\&\N__17696\&\N__14429\&\N__15209\&\N__14726\;
    \line_buffer.mem31_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem31_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9335\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19133\&'0'&'0'&'0';
    \line_buffer.n459\ <= \line_buffer.mem9_physical_RDATA_wire\(11);
    \line_buffer.n458\ <= \line_buffer.mem9_physical_RDATA_wire\(3);
    \line_buffer.mem9_physical_RADDR_wire\ <= \N__12548\&\N__10226\&\N__11249\&\N__12800\&\N__13280\&\N__10475\&\N__13055\&\N__10739\&\N__10991\&\N__9995\&\N__14078\;
    \line_buffer.mem9_physical_WADDR_wire\ <= \N__14900\&\N__17879\&\N__17129\&\N__16631\&\N__16883\&\N__19364\&\N__17381\&\N__17624\&\N__14357\&\N__15137\&\N__14654\;
    \line_buffer.mem9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem9_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__15657\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9534\&'0'&'0'&'0';
    \line_buffer.n598\ <= \line_buffer.mem29_physical_RDATA_wire\(11);
    \line_buffer.n597\ <= \line_buffer.mem29_physical_RDATA_wire\(3);
    \line_buffer.mem29_physical_RADDR_wire\ <= \N__12656\&\N__10334\&\N__11357\&\N__12908\&\N__13388\&\N__10583\&\N__13163\&\N__10847\&\N__11099\&\N__10103\&\N__14186\;
    \line_buffer.mem29_physical_WADDR_wire\ <= \N__15008\&\N__17987\&\N__17237\&\N__16739\&\N__16991\&\N__19472\&\N__17489\&\N__17732\&\N__14465\&\N__15245\&\N__14762\;
    \line_buffer.mem29_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem29_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__13554\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21704\&'0'&'0'&'0';
    \line_buffer.n600\ <= \line_buffer.mem6_physical_RDATA_wire\(11);
    \line_buffer.n599\ <= \line_buffer.mem6_physical_RDATA_wire\(3);
    \line_buffer.mem6_physical_RADDR_wire\ <= \N__12584\&\N__10262\&\N__11285\&\N__12836\&\N__13316\&\N__10511\&\N__13091\&\N__10775\&\N__11027\&\N__10031\&\N__14114\;
    \line_buffer.mem6_physical_WADDR_wire\ <= \N__14936\&\N__17915\&\N__17165\&\N__16667\&\N__16919\&\N__19400\&\N__17417\&\N__17660\&\N__14393\&\N__15173\&\N__14690\;
    \line_buffer.mem6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__21052\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19910\&'0'&'0'&'0';
    \line_buffer.n457\ <= \line_buffer.mem10_physical_RDATA_wire\(11);
    \line_buffer.n456\ <= \line_buffer.mem10_physical_RDATA_wire\(3);
    \line_buffer.mem10_physical_RADDR_wire\ <= \N__12713\&\N__10397\&\N__11396\&\N__12965\&\N__13439\&\N__10652\&\N__13220\&\N__10916\&\N__11168\&\N__10148\&\N__14249\;
    \line_buffer.mem10_physical_WADDR_wire\ <= \N__15059\&\N__18038\&\N__17288\&\N__16784\&\N__17036\&\N__19517\&\N__17540\&\N__17789\&\N__14522\&\N__15296\&\N__14813\;
    \line_buffer.mem10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem10_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9310\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19140\&'0'&'0'&'0';
    \line_buffer.n586\ <= \line_buffer.mem22_physical_RDATA_wire\(11);
    \line_buffer.n585\ <= \line_buffer.mem22_physical_RDATA_wire\(3);
    \line_buffer.mem22_physical_RADDR_wire\ <= \N__12557\&\N__10241\&\N__11240\&\N__12809\&\N__13283\&\N__10496\&\N__13064\&\N__10760\&\N__11012\&\N__9992\&\N__14093\;
    \line_buffer.mem22_physical_WADDR_wire\ <= \N__14903\&\N__17882\&\N__17132\&\N__16628\&\N__16880\&\N__19361\&\N__17384\&\N__17633\&\N__14366\&\N__15140\&\N__14657\;
    \line_buffer.mem22_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem22_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9339\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19155\&'0'&'0'&'0';
    \line_buffer.n530\ <= \line_buffer.mem25_physical_RDATA_wire\(11);
    \line_buffer.n529\ <= \line_buffer.mem25_physical_RDATA_wire\(3);
    \line_buffer.mem25_physical_RADDR_wire\ <= \N__12704\&\N__10382\&\N__11405\&\N__12956\&\N__13436\&\N__10631\&\N__13211\&\N__10895\&\N__11147\&\N__10151\&\N__14234\;
    \line_buffer.mem25_physical_WADDR_wire\ <= \N__15056\&\N__18035\&\N__17285\&\N__16787\&\N__17039\&\N__19520\&\N__17537\&\N__17780\&\N__14513\&\N__15293\&\N__14810\;
    \line_buffer.mem25_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem25_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9303\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19141\&'0'&'0'&'0';
    \line_buffer.n461\ <= \line_buffer.mem8_physical_RDATA_wire\(11);
    \line_buffer.n460\ <= \line_buffer.mem8_physical_RDATA_wire\(3);
    \line_buffer.mem8_physical_RADDR_wire\ <= \N__12560\&\N__10238\&\N__11261\&\N__12812\&\N__13292\&\N__10487\&\N__13067\&\N__10751\&\N__11003\&\N__10007\&\N__14090\;
    \line_buffer.mem8_physical_WADDR_wire\ <= \N__14912\&\N__17891\&\N__17141\&\N__16643\&\N__16895\&\N__19376\&\N__17393\&\N__17636\&\N__14369\&\N__15149\&\N__14666\;
    \line_buffer.mem8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem8_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__13581\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21725\&'0'&'0'&'0';
    \line_buffer.n562\ <= \line_buffer.mem28_physical_RDATA_wire\(11);
    \line_buffer.n561\ <= \line_buffer.mem28_physical_RDATA_wire\(3);
    \line_buffer.mem28_physical_RADDR_wire\ <= \N__12668\&\N__10346\&\N__11369\&\N__12920\&\N__13400\&\N__10595\&\N__13175\&\N__10859\&\N__11111\&\N__10115\&\N__14198\;
    \line_buffer.mem28_physical_WADDR_wire\ <= \N__15020\&\N__17999\&\N__17249\&\N__16751\&\N__17003\&\N__19484\&\N__17501\&\N__17744\&\N__14477\&\N__15257\&\N__14774\;
    \line_buffer.mem28_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem28_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9318\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19129\&'0'&'0'&'0';
    \line_buffer.n467\ <= \line_buffer.mem18_physical_RDATA_wire\(11);
    \line_buffer.n466\ <= \line_buffer.mem18_physical_RDATA_wire\(3);
    \line_buffer.mem18_physical_RADDR_wire\ <= \N__12617\&\N__10301\&\N__11300\&\N__12869\&\N__13343\&\N__10556\&\N__13124\&\N__10820\&\N__11072\&\N__10052\&\N__14153\;
    \line_buffer.mem18_physical_WADDR_wire\ <= \N__14963\&\N__17942\&\N__17192\&\N__16688\&\N__16940\&\N__19421\&\N__17444\&\N__17693\&\N__14426\&\N__15200\&\N__14717\;
    \line_buffer.mem18_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem18_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__15631\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9515\&'0'&'0'&'0';

    \tx_pll.TX_PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0100110",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \ADV_CLK_c\,
            REFERENCECLK => \N__18215\,
            RESETB => \N__22064\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \line_buffer.mem2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem2_physical_RDATA_wire\,
            RADDR => \line_buffer.mem2_physical_RADDR_wire\,
            WADDR => \line_buffer.mem2_physical_WADDR_wire\,
            MASK => \line_buffer.mem2_physical_MASK_wire\,
            WDATA => \line_buffer.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23950\,
            RE => \N__22138\,
            WCLKE => 'H',
            WCLK => \N__21988\,
            WE => \N__18108\
        );

    \line_buffer.mem14_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem14_physical_RDATA_wire\,
            RADDR => \line_buffer.mem14_physical_RADDR_wire\,
            WADDR => \line_buffer.mem14_physical_WADDR_wire\,
            MASK => \line_buffer.mem14_physical_MASK_wire\,
            WDATA => \line_buffer.mem14_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24336\,
            RE => \N__22211\,
            WCLKE => 'H',
            WCLK => \N__21972\,
            WE => \N__16466\
        );

    \line_buffer.mem5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem5_physical_RDATA_wire\,
            RADDR => \line_buffer.mem5_physical_RADDR_wire\,
            WADDR => \line_buffer.mem5_physical_WADDR_wire\,
            MASK => \line_buffer.mem5_physical_MASK_wire\,
            WDATA => \line_buffer.mem5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23616\,
            RE => \N__22202\,
            WCLKE => 'H',
            WCLK => \N__21986\,
            WE => \N__16427\
        );

    \line_buffer.mem11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem11_physical_RDATA_wire\,
            RADDR => \line_buffer.mem11_physical_RADDR_wire\,
            WADDR => \line_buffer.mem11_physical_WADDR_wire\,
            MASK => \line_buffer.mem11_physical_MASK_wire\,
            WDATA => \line_buffer.mem11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24138\,
            RE => \N__22236\,
            WCLKE => 'H',
            WCLK => \N__21961\,
            WE => \N__18725\
        );

    \line_buffer.mem21_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem21_physical_RDATA_wire\,
            RADDR => \line_buffer.mem21_physical_RADDR_wire\,
            WADDR => \line_buffer.mem21_physical_WADDR_wire\,
            MASK => \line_buffer.mem21_physical_MASK_wire\,
            WDATA => \line_buffer.mem21_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23811\,
            RE => \N__22099\,
            WCLKE => 'H',
            WCLK => \N__21992\,
            WE => \N__18271\
        );

    \line_buffer.mem12_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem12_physical_RDATA_wire\,
            RADDR => \line_buffer.mem12_physical_RADDR_wire\,
            WADDR => \line_buffer.mem12_physical_WADDR_wire\,
            MASK => \line_buffer.mem12_physical_MASK_wire\,
            WDATA => \line_buffer.mem12_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24001\,
            RE => \N__22235\,
            WCLKE => 'H',
            WCLK => \N__21963\,
            WE => \N__18718\
        );

    \line_buffer.mem24_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem24_physical_RDATA_wire\,
            RADDR => \line_buffer.mem24_physical_RADDR_wire\,
            WADDR => \line_buffer.mem24_physical_WADDR_wire\,
            MASK => \line_buffer.mem24_physical_MASK_wire\,
            WDATA => \line_buffer.mem24_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24362\,
            RE => \N__22322\,
            WCLKE => 'H',
            WCLK => \N__21950\,
            WE => \N__16103\
        );

    \line_buffer.mem1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem1_physical_RDATA_wire\,
            RADDR => \line_buffer.mem1_physical_RADDR_wire\,
            WADDR => \line_buffer.mem1_physical_WADDR_wire\,
            MASK => \line_buffer.mem1_physical_MASK_wire\,
            WDATA => \line_buffer.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24248\,
            RE => \N__22256\,
            WCLKE => 'H',
            WCLK => \N__21945\,
            WE => \N__16473\
        );

    \line_buffer.mem15_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem15_physical_RDATA_wire\,
            RADDR => \line_buffer.mem15_physical_RADDR_wire\,
            WADDR => \line_buffer.mem15_physical_WADDR_wire\,
            MASK => \line_buffer.mem15_physical_MASK_wire\,
            WDATA => \line_buffer.mem15_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24114\,
            RE => \N__22188\,
            WCLKE => 'H',
            WCLK => \N__21974\,
            WE => \N__16464\
        );

    \line_buffer.mem27_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem27_physical_RDATA_wire\,
            RADDR => \line_buffer.mem27_physical_RADDR_wire\,
            WADDR => \line_buffer.mem27_physical_WADDR_wire\,
            MASK => \line_buffer.mem27_physical_MASK_wire\,
            WDATA => \line_buffer.mem27_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24337\,
            RE => \N__22297\,
            WCLKE => 'H',
            WCLK => \N__21964\,
            WE => \N__16423\
        );

    \line_buffer.mem4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem4_physical_RDATA_wire\,
            RADDR => \line_buffer.mem4_physical_RADDR_wire\,
            WADDR => \line_buffer.mem4_physical_WADDR_wire\,
            MASK => \line_buffer.mem4_physical_MASK_wire\,
            WDATA => \line_buffer.mem4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23948\,
            RE => \N__22226\,
            WCLKE => 'H',
            WCLK => \N__21984\,
            WE => \N__16087\
        );

    \line_buffer.mem16_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem16_physical_RDATA_wire\,
            RADDR => \line_buffer.mem16_physical_RADDR_wire\,
            WADDR => \line_buffer.mem16_physical_WADDR_wire\,
            MASK => \line_buffer.mem16_physical_MASK_wire\,
            WDATA => \line_buffer.mem16_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24294\,
            RE => \N__22187\,
            WCLKE => 'H',
            WCLK => \N__21976\,
            WE => \N__16465\
        );

    \line_buffer.mem30_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem30_physical_RDATA_wire\,
            RADDR => \line_buffer.mem30_physical_RADDR_wire\,
            WADDR => \line_buffer.mem30_physical_WADDR_wire\,
            MASK => \line_buffer.mem30_physical_MASK_wire\,
            WDATA => \line_buffer.mem30_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24204\,
            RE => \N__22260\,
            WCLKE => 'H',
            WCLK => \N__21977\,
            WE => \N__16141\
        );

    \line_buffer.mem7_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem7_physical_RDATA_wire\,
            RADDR => \line_buffer.mem7_physical_RADDR_wire\,
            WADDR => \line_buffer.mem7_physical_WADDR_wire\,
            MASK => \line_buffer.mem7_physical_MASK_wire\,
            WDATA => \line_buffer.mem7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23807\,
            RE => \N__22154\,
            WCLKE => 'H',
            WCLK => \N__21991\,
            WE => \N__16528\
        );

    \line_buffer.mem20_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem20_physical_RDATA_wire\,
            RADDR => \line_buffer.mem20_physical_RADDR_wire\,
            WADDR => \line_buffer.mem20_physical_WADDR_wire\,
            MASK => \line_buffer.mem20_physical_MASK_wire\,
            WDATA => \line_buffer.mem20_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23909\,
            RE => \N__22112\,
            WCLKE => 'H',
            WCLK => \N__21990\,
            WE => \N__18270\
        );

    \line_buffer.mem13_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem13_physical_RDATA_wire\,
            RADDR => \line_buffer.mem13_physical_RADDR_wire\,
            WADDR => \line_buffer.mem13_physical_WADDR_wire\,
            MASK => \line_buffer.mem13_physical_MASK_wire\,
            WDATA => \line_buffer.mem13_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23869\,
            RE => \N__22212\,
            WCLKE => 'H',
            WCLK => \N__21967\,
            WE => \N__18717\
        );

    \line_buffer.mem19_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem19_physical_RDATA_wire\,
            RADDR => \line_buffer.mem19_physical_RADDR_wire\,
            WADDR => \line_buffer.mem19_physical_WADDR_wire\,
            MASK => \line_buffer.mem19_physical_MASK_wire\,
            WDATA => \line_buffer.mem19_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23735\,
            RE => \N__22139\,
            WCLKE => 'H',
            WCLK => \N__21985\,
            WE => \N__18097\
        );

    \line_buffer.mem23_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem23_physical_RDATA_wire\,
            RADDR => \line_buffer.mem23_physical_RADDR_wire\,
            WADDR => \line_buffer.mem23_physical_WADDR_wire\,
            MASK => \line_buffer.mem23_physical_MASK_wire\,
            WDATA => \line_buffer.mem23_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24363\,
            RE => \N__22326\,
            WCLKE => 'H',
            WCLK => \N__21939\,
            WE => \N__16104\
        );

    \line_buffer.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem0_physical_RDATA_wire\,
            RADDR => \line_buffer.mem0_physical_RADDR_wire\,
            WADDR => \line_buffer.mem0_physical_WADDR_wire\,
            MASK => \line_buffer.mem0_physical_MASK_wire\,
            WDATA => \line_buffer.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24249\,
            RE => \N__22269\,
            WCLKE => 'H',
            WCLK => \N__21934\,
            WE => \N__18729\
        );

    \line_buffer.mem26_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem26_physical_RDATA_wire\,
            RADDR => \line_buffer.mem26_physical_RADDR_wire\,
            WADDR => \line_buffer.mem26_physical_WADDR_wire\,
            MASK => \line_buffer.mem26_physical_MASK_wire\,
            WDATA => \line_buffer.mem26_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24354\,
            RE => \N__22306\,
            WCLKE => 'H',
            WCLK => \N__21962\,
            WE => \N__16428\
        );

    \line_buffer.mem3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem3_physical_RDATA_wire\,
            RADDR => \line_buffer.mem3_physical_RADDR_wire\,
            WADDR => \line_buffer.mem3_physical_WADDR_wire\,
            MASK => \line_buffer.mem3_physical_MASK_wire\,
            WDATA => \line_buffer.mem3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24293\,
            RE => \N__22270\,
            WCLKE => 'H',
            WCLK => \N__21975\,
            WE => \N__18275\
        );

    \line_buffer.mem17_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem17_physical_RDATA_wire\,
            RADDR => \line_buffer.mem17_physical_RADDR_wire\,
            WADDR => \line_buffer.mem17_physical_WADDR_wire\,
            MASK => \line_buffer.mem17_physical_MASK_wire\,
            WDATA => \line_buffer.mem17_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23980\,
            RE => \N__22164\,
            WCLKE => 'H',
            WCLK => \N__21981\,
            WE => \N__18091\
        );

    \line_buffer.mem31_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem31_physical_RDATA_wire\,
            RADDR => \line_buffer.mem31_physical_RADDR_wire\,
            WADDR => \line_buffer.mem31_physical_WADDR_wire\,
            MASK => \line_buffer.mem31_physical_MASK_wire\,
            WDATA => \line_buffer.mem31_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23979\,
            RE => \N__22246\,
            WCLKE => 'H',
            WCLK => \N__21982\,
            WE => \N__16148\
        );

    \line_buffer.mem9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem9_physical_RDATA_wire\,
            RADDR => \line_buffer.mem9_physical_RADDR_wire\,
            WADDR => \line_buffer.mem9_physical_WADDR_wire\,
            MASK => \line_buffer.mem9_physical_MASK_wire\,
            WDATA => \line_buffer.mem9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23643\,
            RE => \N__22153\,
            WCLKE => 'H',
            WCLK => \N__21995\,
            WE => \N__16532\
        );

    \line_buffer.mem29_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem29_physical_RDATA_wire\,
            RADDR => \line_buffer.mem29_physical_RADDR_wire\,
            WADDR => \line_buffer.mem29_physical_WADDR_wire\,
            MASK => \line_buffer.mem29_physical_MASK_wire\,
            WDATA => \line_buffer.mem29_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24313\,
            RE => \N__22279\,
            WCLKE => 'H',
            WCLK => \N__21973\,
            WE => \N__16140\
        );

    \line_buffer.mem6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem6_physical_RDATA_wire\,
            RADDR => \line_buffer.mem6_physical_RADDR_wire\,
            WADDR => \line_buffer.mem6_physical_WADDR_wire\,
            MASK => \line_buffer.mem6_physical_MASK_wire\,
            WDATA => \line_buffer.mem6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23949\,
            RE => \N__22178\,
            WCLKE => 'H',
            WCLK => \N__21989\,
            WE => \N__16152\
        );

    \line_buffer.mem10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem10_physical_RDATA_wire\,
            RADDR => \line_buffer.mem10_physical_RADDR_wire\,
            WADDR => \line_buffer.mem10_physical_WADDR_wire\,
            MASK => \line_buffer.mem10_physical_MASK_wire\,
            WDATA => \line_buffer.mem10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24139\,
            RE => \N__22255\,
            WCLKE => 'H',
            WCLK => \N__21954\,
            WE => \N__16533\
        );

    \line_buffer.mem22_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem22_physical_RDATA_wire\,
            RADDR => \line_buffer.mem22_physical_RADDR_wire\,
            WADDR => \line_buffer.mem22_physical_WADDR_wire\,
            MASK => \line_buffer.mem22_physical_MASK_wire\,
            WDATA => \line_buffer.mem22_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23764\,
            RE => \N__22111\,
            WCLKE => 'H',
            WCLK => \N__21994\,
            WE => \N__18276\
        );

    \line_buffer.mem25_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem25_physical_RDATA_wire\,
            RADDR => \line_buffer.mem25_physical_RADDR_wire\,
            WADDR => \line_buffer.mem25_physical_WADDR_wire\,
            MASK => \line_buffer.mem25_physical_MASK_wire\,
            WDATA => \line_buffer.mem25_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24355\,
            RE => \N__22315\,
            WCLKE => 'H',
            WCLK => \N__21956\,
            WE => \N__16096\
        );

    \line_buffer.mem8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem8_physical_RDATA_wire\,
            RADDR => \line_buffer.mem8_physical_RADDR_wire\,
            WADDR => \line_buffer.mem8_physical_WADDR_wire\,
            MASK => \line_buffer.mem8_physical_MASK_wire\,
            WDATA => \line_buffer.mem8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23681\,
            RE => \N__22126\,
            WCLKE => 'H',
            WCLK => \N__21993\,
            WE => \N__16527\
        );

    \line_buffer.mem28_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem28_physical_RDATA_wire\,
            RADDR => \line_buffer.mem28_physical_RADDR_wire\,
            WADDR => \line_buffer.mem28_physical_WADDR_wire\,
            MASK => \line_buffer.mem28_physical_MASK_wire\,
            WDATA => \line_buffer.mem28_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23745\,
            RE => \N__22288\,
            WCLKE => 'H',
            WCLK => \N__21970\,
            WE => \N__16413\
        );

    \line_buffer.mem18_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem18_physical_RDATA_wire\,
            RADDR => \line_buffer.mem18_physical_RADDR_wire\,
            WADDR => \line_buffer.mem18_physical_WADDR_wire\,
            MASK => \line_buffer.mem18_physical_MASK_wire\,
            WDATA => \line_buffer.mem18_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24065\,
            RE => \N__22163\,
            WCLKE => 'H',
            WCLK => \N__21983\,
            WE => \N__18104\
        );

    \DEBUG_c_3_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__24832\,
            GLOBALBUFFEROUTPUT => \DEBUG_c_3_c\
        );

    \DEBUG_c_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24834\,
            DIN => \N__24833\,
            DOUT => \N__24832\,
            PACKAGEPIN => \TVP_CLK_wire\
        );

    \DEBUG_c_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24834\,
            PADOUT => \N__24833\,
            PADIN => \N__24832\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24823\,
            DIN => \N__24822\,
            DOUT => \N__24821\,
            PACKAGEPIN => \ADV_CLK_wire\
        );

    \ADV_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24823\,
            PADOUT => \N__24822\,
            PADIN => \N__24821\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24064\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24814\,
            DIN => \N__24813\,
            DOUT => \N__24812\,
            PACKAGEPIN => \TVP_HSYNC_wire\
        );

    \DEBUG_c_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24814\,
            PADOUT => \N__24813\,
            PADIN => \N__24812\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_2_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24805\,
            DIN => \N__24804\,
            DOUT => \N__24803\,
            PACKAGEPIN => DEBUG(3)
        );

    \DEBUG_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24805\,
            PADOUT => \N__24804\,
            PADIN => \N__24803\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18225\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24796\,
            DIN => \N__24795\,
            DOUT => \N__24794\,
            PACKAGEPIN => \TVP_VIDEO_wire\(2)
        );

    \TVP_VIDEO_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24796\,
            PADOUT => \N__24795\,
            PADIN => \N__24794\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24787\,
            DIN => \N__24786\,
            DOUT => \N__24785\,
            PACKAGEPIN => \ADV_G_wire\(5)
        );

    \ADV_G_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24787\,
            PADOUT => \N__24786\,
            PADIN => \N__24785\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20762\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24778\,
            DIN => \N__24777\,
            DOUT => \N__24776\,
            PACKAGEPIN => \ADV_R_wire\(3)
        );

    \ADV_R_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24778\,
            PADOUT => \N__24777\,
            PADIN => \N__24776\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18337\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24769\,
            DIN => \N__24768\,
            DOUT => \N__24767\,
            PACKAGEPIN => \ADV_R_wire\(0)
        );

    \ADV_R_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24769\,
            PADOUT => \N__24768\,
            PADIN => \N__24767\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14598\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24760\,
            DIN => \N__24759\,
            DOUT => \N__24758\,
            PACKAGEPIN => DEBUG(2)
        );

    \DEBUG_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24760\,
            PADOUT => \N__24759\,
            PADIN => \N__24758\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20181\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24751\,
            DIN => \N__24750\,
            DOUT => \N__24749\,
            PACKAGEPIN => \TVP_VIDEO_wire\(3)
        );

    \TVP_VIDEO_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24751\,
            PADOUT => \N__24750\,
            PADIN => \N__24749\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24742\,
            DIN => \N__24741\,
            DOUT => \N__24740\,
            PACKAGEPIN => \ADV_G_wire\(4)
        );

    \ADV_G_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24742\,
            PADOUT => \N__24741\,
            PADIN => \N__24740\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22548\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24733\,
            DIN => \N__24732\,
            DOUT => \N__24731\,
            PACKAGEPIN => \ADV_R_wire\(5)
        );

    \ADV_R_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24733\,
            PADOUT => \N__24732\,
            PADIN => \N__24731\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20766\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24724\,
            DIN => \N__24723\,
            DOUT => \N__24722\,
            PACKAGEPIN => \TVP_VIDEO_wire\(9)
        );

    \TVP_VIDEO_pad_9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24724\,
            PADOUT => \N__24723\,
            PADIN => \N__24722\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24715\,
            DIN => \N__24714\,
            DOUT => \N__24713\,
            PACKAGEPIN => DEBUG(1)
        );

    \DEBUG_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24715\,
            PADOUT => \N__24714\,
            PADIN => \N__24713\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13623\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24706\,
            DIN => \N__24705\,
            DOUT => \N__24704\,
            PACKAGEPIN => \TVP_VIDEO_wire\(7)
        );

    \DEBUG_c_6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24706\,
            PADOUT => \N__24705\,
            PADIN => \N__24704\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_6_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24697\,
            DIN => \N__24696\,
            DOUT => \N__24695\,
            PACKAGEPIN => \ADV_B_wire\(1)
        );

    \ADV_B_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24697\,
            PADOUT => \N__24696\,
            PADIN => \N__24695\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20678\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_SYNC_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24688\,
            DIN => \N__24687\,
            DOUT => \N__24686\,
            PACKAGEPIN => \ADV_SYNC_N_wire\
        );

    \ADV_SYNC_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24688\,
            PADOUT => \N__24687\,
            PADIN => \N__24686\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24679\,
            DIN => \N__24678\,
            DOUT => \N__24677\,
            PACKAGEPIN => \ADV_B_wire\(6)
        );

    \ADV_B_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24679\,
            PADOUT => \N__24678\,
            PADIN => \N__24677\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22481\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24670\,
            DIN => \N__24669\,
            DOUT => \N__24668\,
            PACKAGEPIN => DEBUG(6)
        );

    \DEBUG_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24670\,
            PADOUT => \N__24669\,
            PADIN => \N__24668\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9240\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24661\,
            DIN => \N__24660\,
            DOUT => \N__24659\,
            PACKAGEPIN => \ADV_G_wire\(0)
        );

    \ADV_G_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24661\,
            PADOUT => \N__24660\,
            PADIN => \N__24659\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24652\,
            DIN => \N__24651\,
            DOUT => \N__24650\,
            PACKAGEPIN => \ADV_R_wire\(1)
        );

    \ADV_R_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24652\,
            PADOUT => \N__24651\,
            PADIN => \N__24650\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20696\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24643\,
            DIN => \N__24642\,
            DOUT => \N__24641\,
            PACKAGEPIN => DEBUG(5)
        );

    \DEBUG_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24643\,
            PADOUT => \N__24642\,
            PADIN => \N__24641\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21627\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24634\,
            DIN => \N__24633\,
            DOUT => \N__24632\,
            PACKAGEPIN => \ADV_G_wire\(7)
        );

    \ADV_G_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24634\,
            PADOUT => \N__24633\,
            PADIN => \N__24632\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11519\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24625\,
            DIN => \N__24624\,
            DOUT => \N__24623\,
            PACKAGEPIN => \ADV_R_wire\(6)
        );

    \ADV_R_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24625\,
            PADOUT => \N__24624\,
            PADIN => \N__24623\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22488\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_BLANK_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24616\,
            DIN => \N__24615\,
            DOUT => \N__24614\,
            PACKAGEPIN => \ADV_BLANK_N_wire\
        );

    \ADV_BLANK_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24616\,
            PADOUT => \N__24615\,
            PADIN => \N__24614\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22060\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24607\,
            DIN => \N__24606\,
            DOUT => \N__24605\,
            PACKAGEPIN => DEBUG(0)
        );

    \DEBUG_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24607\,
            PADOUT => \N__24606\,
            PADIN => \N__24605\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18186\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24598\,
            DIN => \N__24597\,
            DOUT => \N__24596\,
            PACKAGEPIN => \ADV_B_wire\(2)
        );

    \ADV_B_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24598\,
            PADOUT => \N__24597\,
            PADIN => \N__24596\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9419\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24589\,
            DIN => \N__24588\,
            DOUT => \N__24587\,
            PACKAGEPIN => \TVP_VIDEO_wire\(8)
        );

    \DEBUG_c_7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24589\,
            PADOUT => \N__24588\,
            PADIN => \N__24587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_7_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24580\,
            DIN => \N__24579\,
            DOUT => \N__24578\,
            PACKAGEPIN => \TVP_VSYNC_wire\
        );

    \DEBUG_c_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24580\,
            PADOUT => \N__24579\,
            PADIN => \N__24578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24571\,
            DIN => \N__24570\,
            DOUT => \N__24569\,
            PACKAGEPIN => \TVP_VIDEO_wire\(6)
        );

    \DEBUG_c_5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24571\,
            PADOUT => \N__24570\,
            PADIN => \N__24569\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_5_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24562\,
            DIN => \N__24561\,
            DOUT => \N__24560\,
            PACKAGEPIN => \ADV_B_wire\(7)
        );

    \ADV_B_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24562\,
            PADOUT => \N__24561\,
            PADIN => \N__24560\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11518\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24553\,
            DIN => \N__24552\,
            DOUT => \N__24551\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24553\,
            PADOUT => \N__24552\,
            PADIN => \N__24551\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18147\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24544\,
            DIN => \N__24543\,
            DOUT => \N__24542\,
            PACKAGEPIN => \TVP_VIDEO_wire\(4)
        );

    \TVP_VIDEO_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24544\,
            PADOUT => \N__24543\,
            PADIN => \N__24542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24535\,
            DIN => \N__24534\,
            DOUT => \N__24533\,
            PACKAGEPIN => \ADV_G_wire\(3)
        );

    \ADV_G_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24535\,
            PADOUT => \N__24534\,
            PADIN => \N__24533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18339\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24526\,
            DIN => \N__24525\,
            DOUT => \N__24524\,
            PACKAGEPIN => \ADV_HSYNC_wire\
        );

    \ADV_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24526\,
            PADOUT => \N__24525\,
            PADIN => \N__24524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11832\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24517\,
            DIN => \N__24516\,
            DOUT => \N__24515\,
            PACKAGEPIN => \ADV_R_wire\(2)
        );

    \ADV_R_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24517\,
            PADOUT => \N__24516\,
            PADIN => \N__24515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24508\,
            DIN => \N__24507\,
            DOUT => \N__24506\,
            PACKAGEPIN => \ADV_B_wire\(4)
        );

    \ADV_B_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24508\,
            PADOUT => \N__24507\,
            PADIN => \N__24506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22531\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24499\,
            DIN => \N__24498\,
            DOUT => \N__24497\,
            PACKAGEPIN => DEBUG(4)
        );

    \DEBUG_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24499\,
            PADOUT => \N__24498\,
            PADIN => \N__24497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19701\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24490\,
            DIN => \N__24489\,
            DOUT => \N__24488\,
            PACKAGEPIN => \ADV_G_wire\(6)
        );

    \ADV_G_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24490\,
            PADOUT => \N__24489\,
            PADIN => \N__24488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22477\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24481\,
            DIN => \N__24480\,
            DOUT => \N__24479\,
            PACKAGEPIN => \ADV_R_wire\(7)
        );

    \ADV_R_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24481\,
            PADOUT => \N__24480\,
            PADIN => \N__24479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24472\,
            DIN => \N__24471\,
            DOUT => \N__24470\,
            PACKAGEPIN => \ADV_B_wire\(3)
        );

    \ADV_B_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24472\,
            PADOUT => \N__24471\,
            PADIN => \N__24470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18338\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24463\,
            DIN => \N__24462\,
            DOUT => \N__24461\,
            PACKAGEPIN => \ADV_R_wire\(4)
        );

    \ADV_R_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24463\,
            PADOUT => \N__24462\,
            PADIN => \N__24461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22538\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24454\,
            DIN => \N__24453\,
            DOUT => \N__24452\,
            PACKAGEPIN => \ADV_B_wire\(0)
        );

    \ADV_B_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24454\,
            PADOUT => \N__24453\,
            PADIN => \N__24452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24445\,
            DIN => \N__24444\,
            DOUT => \N__24443\,
            PACKAGEPIN => \TVP_VIDEO_wire\(5)
        );

    \TVP_VIDEO_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24445\,
            PADOUT => \N__24444\,
            PADIN => \N__24443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24436\,
            DIN => \N__24435\,
            DOUT => \N__24434\,
            PACKAGEPIN => \ADV_G_wire\(2)
        );

    \ADV_G_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24436\,
            PADOUT => \N__24435\,
            PADIN => \N__24434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9420\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24427\,
            DIN => \N__24426\,
            DOUT => \N__24425\,
            PACKAGEPIN => \ADV_VSYNC_wire\
        );

    \ADV_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24427\,
            PADOUT => \N__24426\,
            PADIN => \N__24425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23346\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24418\,
            DIN => \N__24417\,
            DOUT => \N__24416\,
            PACKAGEPIN => \ADV_B_wire\(5)
        );

    \ADV_B_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24418\,
            PADOUT => \N__24417\,
            PADIN => \N__24416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20743\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24409\,
            DIN => \N__24408\,
            DOUT => \N__24407\,
            PACKAGEPIN => DEBUG(7)
        );

    \DEBUG_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24409\,
            PADOUT => \N__24408\,
            PADIN => \N__24407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19965\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24400\,
            DIN => \N__24399\,
            DOUT => \N__24398\,
            PACKAGEPIN => \ADV_G_wire\(1)
        );

    \ADV_G_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24400\,
            PADOUT => \N__24399\,
            PADIN => \N__24398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20700\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5856\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24378\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__24378\,
            I => \transmit_module.Y_DELTA_PATTERN_85\
        );

    \I__5854\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24372\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__24372\,
            I => \transmit_module.Y_DELTA_PATTERN_87\
        );

    \I__5852\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24366\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__24366\,
            I => \transmit_module.Y_DELTA_PATTERN_86\
        );

    \I__5850\ : ClkMux
    port map (
            O => \N__24363\,
            I => \N__24359\
        );

    \I__5849\ : ClkMux
    port map (
            O => \N__24362\,
            I => \N__24356\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24344\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__24356\,
            I => \N__24344\
        );

    \I__5846\ : ClkMux
    port map (
            O => \N__24355\,
            I => \N__24341\
        );

    \I__5845\ : ClkMux
    port map (
            O => \N__24354\,
            I => \N__24338\
        );

    \I__5844\ : ClkMux
    port map (
            O => \N__24353\,
            I => \N__24328\
        );

    \I__5843\ : ClkMux
    port map (
            O => \N__24352\,
            I => \N__24325\
        );

    \I__5842\ : ClkMux
    port map (
            O => \N__24351\,
            I => \N__24322\
        );

    \I__5841\ : ClkMux
    port map (
            O => \N__24350\,
            I => \N__24319\
        );

    \I__5840\ : ClkMux
    port map (
            O => \N__24349\,
            I => \N__24316\
        );

    \I__5839\ : Span4Mux_s2_v
    port map (
            O => \N__24344\,
            I => \N__24305\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__24341\,
            I => \N__24305\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__24338\,
            I => \N__24305\
        );

    \I__5836\ : ClkMux
    port map (
            O => \N__24337\,
            I => \N__24302\
        );

    \I__5835\ : ClkMux
    port map (
            O => \N__24336\,
            I => \N__24296\
        );

    \I__5834\ : ClkMux
    port map (
            O => \N__24335\,
            I => \N__24288\
        );

    \I__5833\ : ClkMux
    port map (
            O => \N__24334\,
            I => \N__24284\
        );

    \I__5832\ : ClkMux
    port map (
            O => \N__24333\,
            I => \N__24280\
        );

    \I__5831\ : ClkMux
    port map (
            O => \N__24332\,
            I => \N__24277\
        );

    \I__5830\ : ClkMux
    port map (
            O => \N__24331\,
            I => \N__24274\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__24328\,
            I => \N__24267\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__24325\,
            I => \N__24258\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__24322\,
            I => \N__24258\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__24319\,
            I => \N__24258\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__24316\,
            I => \N__24258\
        );

    \I__5824\ : ClkMux
    port map (
            O => \N__24315\,
            I => \N__24255\
        );

    \I__5823\ : ClkMux
    port map (
            O => \N__24314\,
            I => \N__24252\
        );

    \I__5822\ : ClkMux
    port map (
            O => \N__24313\,
            I => \N__24245\
        );

    \I__5821\ : ClkMux
    port map (
            O => \N__24312\,
            I => \N__24242\
        );

    \I__5820\ : Span4Mux_v
    port map (
            O => \N__24305\,
            I => \N__24236\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24236\
        );

    \I__5818\ : ClkMux
    port map (
            O => \N__24301\,
            I => \N__24233\
        );

    \I__5817\ : ClkMux
    port map (
            O => \N__24300\,
            I => \N__24230\
        );

    \I__5816\ : ClkMux
    port map (
            O => \N__24299\,
            I => \N__24224\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__24296\,
            I => \N__24217\
        );

    \I__5814\ : ClkMux
    port map (
            O => \N__24295\,
            I => \N__24214\
        );

    \I__5813\ : ClkMux
    port map (
            O => \N__24294\,
            I => \N__24210\
        );

    \I__5812\ : ClkMux
    port map (
            O => \N__24293\,
            I => \N__24205\
        );

    \I__5811\ : ClkMux
    port map (
            O => \N__24292\,
            I => \N__24201\
        );

    \I__5810\ : ClkMux
    port map (
            O => \N__24291\,
            I => \N__24198\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__24288\,
            I => \N__24194\
        );

    \I__5808\ : ClkMux
    port map (
            O => \N__24287\,
            I => \N__24191\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__24284\,
            I => \N__24188\
        );

    \I__5806\ : ClkMux
    port map (
            O => \N__24283\,
            I => \N__24185\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__24280\,
            I => \N__24181\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__24277\,
            I => \N__24176\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__24274\,
            I => \N__24176\
        );

    \I__5802\ : ClkMux
    port map (
            O => \N__24273\,
            I => \N__24173\
        );

    \I__5801\ : ClkMux
    port map (
            O => \N__24272\,
            I => \N__24170\
        );

    \I__5800\ : ClkMux
    port map (
            O => \N__24271\,
            I => \N__24167\
        );

    \I__5799\ : ClkMux
    port map (
            O => \N__24270\,
            I => \N__24164\
        );

    \I__5798\ : Span4Mux_v
    port map (
            O => \N__24267\,
            I => \N__24159\
        );

    \I__5797\ : Span4Mux_v
    port map (
            O => \N__24258\,
            I => \N__24159\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__24255\,
            I => \N__24156\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__24252\,
            I => \N__24153\
        );

    \I__5794\ : ClkMux
    port map (
            O => \N__24251\,
            I => \N__24150\
        );

    \I__5793\ : ClkMux
    port map (
            O => \N__24250\,
            I => \N__24147\
        );

    \I__5792\ : ClkMux
    port map (
            O => \N__24249\,
            I => \N__24143\
        );

    \I__5791\ : ClkMux
    port map (
            O => \N__24248\,
            I => \N__24140\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__24245\,
            I => \N__24133\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__24242\,
            I => \N__24133\
        );

    \I__5788\ : ClkMux
    port map (
            O => \N__24241\,
            I => \N__24130\
        );

    \I__5787\ : Span4Mux_v
    port map (
            O => \N__24236\,
            I => \N__24125\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__24233\,
            I => \N__24125\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24122\
        );

    \I__5784\ : ClkMux
    port map (
            O => \N__24229\,
            I => \N__24119\
        );

    \I__5783\ : ClkMux
    port map (
            O => \N__24228\,
            I => \N__24116\
        );

    \I__5782\ : ClkMux
    port map (
            O => \N__24227\,
            I => \N__24109\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__24224\,
            I => \N__24106\
        );

    \I__5780\ : ClkMux
    port map (
            O => \N__24223\,
            I => \N__24103\
        );

    \I__5779\ : ClkMux
    port map (
            O => \N__24222\,
            I => \N__24099\
        );

    \I__5778\ : ClkMux
    port map (
            O => \N__24221\,
            I => \N__24096\
        );

    \I__5777\ : ClkMux
    port map (
            O => \N__24220\,
            I => \N__24093\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__24217\,
            I => \N__24087\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24087\
        );

    \I__5774\ : ClkMux
    port map (
            O => \N__24213\,
            I => \N__24084\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__24210\,
            I => \N__24081\
        );

    \I__5772\ : ClkMux
    port map (
            O => \N__24209\,
            I => \N__24078\
        );

    \I__5771\ : ClkMux
    port map (
            O => \N__24208\,
            I => \N__24075\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__24205\,
            I => \N__24071\
        );

    \I__5769\ : ClkMux
    port map (
            O => \N__24204\,
            I => \N__24068\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__24201\,
            I => \N__24061\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__24198\,
            I => \N__24058\
        );

    \I__5766\ : ClkMux
    port map (
            O => \N__24197\,
            I => \N__24055\
        );

    \I__5765\ : Span4Mux_v
    port map (
            O => \N__24194\,
            I => \N__24050\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__24191\,
            I => \N__24050\
        );

    \I__5763\ : Span4Mux_h
    port map (
            O => \N__24188\,
            I => \N__24045\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24045\
        );

    \I__5761\ : ClkMux
    port map (
            O => \N__24184\,
            I => \N__24042\
        );

    \I__5760\ : Span4Mux_v
    port map (
            O => \N__24181\,
            I => \N__24033\
        );

    \I__5759\ : Span4Mux_h
    port map (
            O => \N__24176\,
            I => \N__24033\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__24173\,
            I => \N__24033\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24033\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__24167\,
            I => \N__24028\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__24164\,
            I => \N__24028\
        );

    \I__5754\ : Span4Mux_h
    port map (
            O => \N__24159\,
            I => \N__24017\
        );

    \I__5753\ : Span4Mux_h
    port map (
            O => \N__24156\,
            I => \N__24017\
        );

    \I__5752\ : Span4Mux_v
    port map (
            O => \N__24153\,
            I => \N__24017\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__24150\,
            I => \N__24017\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__24147\,
            I => \N__24017\
        );

    \I__5749\ : ClkMux
    port map (
            O => \N__24146\,
            I => \N__24014\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__24143\,
            I => \N__24011\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__24140\,
            I => \N__24008\
        );

    \I__5746\ : ClkMux
    port map (
            O => \N__24139\,
            I => \N__24005\
        );

    \I__5745\ : ClkMux
    port map (
            O => \N__24138\,
            I => \N__24002\
        );

    \I__5744\ : Span4Mux_v
    port map (
            O => \N__24133\,
            I => \N__23996\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__23996\
        );

    \I__5742\ : Span4Mux_h
    port map (
            O => \N__24125\,
            I => \N__23987\
        );

    \I__5741\ : Span4Mux_v
    port map (
            O => \N__24122\,
            I => \N__23987\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__24119\,
            I => \N__23987\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__24116\,
            I => \N__23987\
        );

    \I__5738\ : ClkMux
    port map (
            O => \N__24115\,
            I => \N__23984\
        );

    \I__5737\ : ClkMux
    port map (
            O => \N__24114\,
            I => \N__23981\
        );

    \I__5736\ : ClkMux
    port map (
            O => \N__24113\,
            I => \N__23974\
        );

    \I__5735\ : ClkMux
    port map (
            O => \N__24112\,
            I => \N__23969\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__24109\,
            I => \N__23966\
        );

    \I__5733\ : Span4Mux_h
    port map (
            O => \N__24106\,
            I => \N__23961\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__24103\,
            I => \N__23961\
        );

    \I__5731\ : ClkMux
    port map (
            O => \N__24102\,
            I => \N__23958\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__24099\,
            I => \N__23952\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__24096\,
            I => \N__23952\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__24093\,
            I => \N__23945\
        );

    \I__5727\ : ClkMux
    port map (
            O => \N__24092\,
            I => \N__23942\
        );

    \I__5726\ : Span4Mux_h
    port map (
            O => \N__24087\,
            I => \N__23937\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__24084\,
            I => \N__23937\
        );

    \I__5724\ : Span4Mux_h
    port map (
            O => \N__24081\,
            I => \N__23934\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__23931\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__24075\,
            I => \N__23928\
        );

    \I__5721\ : ClkMux
    port map (
            O => \N__24074\,
            I => \N__23925\
        );

    \I__5720\ : Span4Mux_v
    port map (
            O => \N__24071\,
            I => \N__23920\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__23920\
        );

    \I__5718\ : ClkMux
    port map (
            O => \N__24067\,
            I => \N__23917\
        );

    \I__5717\ : ClkMux
    port map (
            O => \N__24066\,
            I => \N__23914\
        );

    \I__5716\ : ClkMux
    port map (
            O => \N__24065\,
            I => \N__23911\
        );

    \I__5715\ : IoInMux
    port map (
            O => \N__24064\,
            I => \N__23906\
        );

    \I__5714\ : Span4Mux_v
    port map (
            O => \N__24061\,
            I => \N__23899\
        );

    \I__5713\ : Span4Mux_v
    port map (
            O => \N__24058\,
            I => \N__23899\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__24055\,
            I => \N__23899\
        );

    \I__5711\ : Span4Mux_h
    port map (
            O => \N__24050\,
            I => \N__23892\
        );

    \I__5710\ : Span4Mux_v
    port map (
            O => \N__24045\,
            I => \N__23892\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__24042\,
            I => \N__23892\
        );

    \I__5708\ : Span4Mux_v
    port map (
            O => \N__24033\,
            I => \N__23883\
        );

    \I__5707\ : Span4Mux_h
    port map (
            O => \N__24028\,
            I => \N__23883\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__24017\,
            I => \N__23883\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__24014\,
            I => \N__23883\
        );

    \I__5704\ : Span4Mux_s2_v
    port map (
            O => \N__24011\,
            I => \N__23876\
        );

    \I__5703\ : Span4Mux_h
    port map (
            O => \N__24008\,
            I => \N__23876\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__24005\,
            I => \N__23876\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23873\
        );

    \I__5700\ : ClkMux
    port map (
            O => \N__24001\,
            I => \N__23870\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__23996\,
            I => \N__23862\
        );

    \I__5698\ : Span4Mux_v
    port map (
            O => \N__23987\,
            I => \N__23862\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__23984\,
            I => \N__23862\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__23981\,
            I => \N__23859\
        );

    \I__5695\ : ClkMux
    port map (
            O => \N__23980\,
            I => \N__23856\
        );

    \I__5694\ : ClkMux
    port map (
            O => \N__23979\,
            I => \N__23853\
        );

    \I__5693\ : ClkMux
    port map (
            O => \N__23978\,
            I => \N__23849\
        );

    \I__5692\ : ClkMux
    port map (
            O => \N__23977\,
            I => \N__23846\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__23974\,
            I => \N__23842\
        );

    \I__5690\ : ClkMux
    port map (
            O => \N__23973\,
            I => \N__23839\
        );

    \I__5689\ : ClkMux
    port map (
            O => \N__23972\,
            I => \N__23836\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__23969\,
            I => \N__23832\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__23966\,
            I => \N__23825\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__23961\,
            I => \N__23825\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__23958\,
            I => \N__23825\
        );

    \I__5684\ : ClkMux
    port map (
            O => \N__23957\,
            I => \N__23822\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__23952\,
            I => \N__23819\
        );

    \I__5682\ : ClkMux
    port map (
            O => \N__23951\,
            I => \N__23816\
        );

    \I__5681\ : ClkMux
    port map (
            O => \N__23950\,
            I => \N__23812\
        );

    \I__5680\ : ClkMux
    port map (
            O => \N__23949\,
            I => \N__23808\
        );

    \I__5679\ : ClkMux
    port map (
            O => \N__23948\,
            I => \N__23804\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__23945\,
            I => \N__23799\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__23942\,
            I => \N__23799\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__23937\,
            I => \N__23795\
        );

    \I__5675\ : Span4Mux_h
    port map (
            O => \N__23934\,
            I => \N__23786\
        );

    \I__5674\ : Span4Mux_v
    port map (
            O => \N__23931\,
            I => \N__23786\
        );

    \I__5673\ : Span4Mux_h
    port map (
            O => \N__23928\,
            I => \N__23786\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__23925\,
            I => \N__23786\
        );

    \I__5671\ : Span4Mux_h
    port map (
            O => \N__23920\,
            I => \N__23779\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__23917\,
            I => \N__23779\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__23914\,
            I => \N__23779\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__23911\,
            I => \N__23776\
        );

    \I__5667\ : ClkMux
    port map (
            O => \N__23910\,
            I => \N__23773\
        );

    \I__5666\ : ClkMux
    port map (
            O => \N__23909\,
            I => \N__23768\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__23906\,
            I => \N__23765\
        );

    \I__5664\ : Span4Mux_h
    port map (
            O => \N__23899\,
            I => \N__23759\
        );

    \I__5663\ : Span4Mux_v
    port map (
            O => \N__23892\,
            I => \N__23759\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__23883\,
            I => \N__23756\
        );

    \I__5661\ : Span4Mux_v
    port map (
            O => \N__23876\,
            I => \N__23749\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__23873\,
            I => \N__23749\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__23870\,
            I => \N__23749\
        );

    \I__5658\ : ClkMux
    port map (
            O => \N__23869\,
            I => \N__23746\
        );

    \I__5657\ : Span4Mux_h
    port map (
            O => \N__23862\,
            I => \N__23742\
        );

    \I__5656\ : Span4Mux_h
    port map (
            O => \N__23859\,
            I => \N__23739\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__23856\,
            I => \N__23736\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__23853\,
            I => \N__23732\
        );

    \I__5653\ : ClkMux
    port map (
            O => \N__23852\,
            I => \N__23729\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__23849\,
            I => \N__23726\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__23846\,
            I => \N__23723\
        );

    \I__5650\ : ClkMux
    port map (
            O => \N__23845\,
            I => \N__23720\
        );

    \I__5649\ : Span4Mux_v
    port map (
            O => \N__23842\,
            I => \N__23713\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23713\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__23836\,
            I => \N__23713\
        );

    \I__5646\ : ClkMux
    port map (
            O => \N__23835\,
            I => \N__23710\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__23832\,
            I => \N__23705\
        );

    \I__5644\ : Span4Mux_v
    port map (
            O => \N__23825\,
            I => \N__23705\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__23822\,
            I => \N__23702\
        );

    \I__5642\ : Span4Mux_v
    port map (
            O => \N__23819\,
            I => \N__23697\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__23816\,
            I => \N__23697\
        );

    \I__5640\ : ClkMux
    port map (
            O => \N__23815\,
            I => \N__23694\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__23812\,
            I => \N__23691\
        );

    \I__5638\ : ClkMux
    port map (
            O => \N__23811\,
            I => \N__23688\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__23808\,
            I => \N__23685\
        );

    \I__5636\ : ClkMux
    port map (
            O => \N__23807\,
            I => \N__23682\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__23804\,
            I => \N__23678\
        );

    \I__5634\ : Span4Mux_v
    port map (
            O => \N__23799\,
            I => \N__23675\
        );

    \I__5633\ : ClkMux
    port map (
            O => \N__23798\,
            I => \N__23672\
        );

    \I__5632\ : Span4Mux_v
    port map (
            O => \N__23795\,
            I => \N__23665\
        );

    \I__5631\ : Span4Mux_h
    port map (
            O => \N__23786\,
            I => \N__23665\
        );

    \I__5630\ : Span4Mux_h
    port map (
            O => \N__23779\,
            I => \N__23665\
        );

    \I__5629\ : Span4Mux_h
    port map (
            O => \N__23776\,
            I => \N__23660\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__23773\,
            I => \N__23660\
        );

    \I__5627\ : ClkMux
    port map (
            O => \N__23772\,
            I => \N__23657\
        );

    \I__5626\ : ClkMux
    port map (
            O => \N__23771\,
            I => \N__23654\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__23768\,
            I => \N__23650\
        );

    \I__5624\ : IoSpan4Mux
    port map (
            O => \N__23765\,
            I => \N__23647\
        );

    \I__5623\ : ClkMux
    port map (
            O => \N__23764\,
            I => \N__23644\
        );

    \I__5622\ : Span4Mux_v
    port map (
            O => \N__23759\,
            I => \N__23640\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__23756\,
            I => \N__23637\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__23749\,
            I => \N__23634\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__23746\,
            I => \N__23631\
        );

    \I__5618\ : ClkMux
    port map (
            O => \N__23745\,
            I => \N__23628\
        );

    \I__5617\ : Span4Mux_v
    port map (
            O => \N__23742\,
            I => \N__23625\
        );

    \I__5616\ : Span4Mux_v
    port map (
            O => \N__23739\,
            I => \N__23620\
        );

    \I__5615\ : Span4Mux_h
    port map (
            O => \N__23736\,
            I => \N__23620\
        );

    \I__5614\ : ClkMux
    port map (
            O => \N__23735\,
            I => \N__23617\
        );

    \I__5613\ : Span4Mux_h
    port map (
            O => \N__23732\,
            I => \N__23611\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__23729\,
            I => \N__23611\
        );

    \I__5611\ : Span4Mux_h
    port map (
            O => \N__23726\,
            I => \N__23604\
        );

    \I__5610\ : Span4Mux_v
    port map (
            O => \N__23723\,
            I => \N__23604\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23604\
        );

    \I__5608\ : Span4Mux_v
    port map (
            O => \N__23713\,
            I => \N__23599\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__23710\,
            I => \N__23599\
        );

    \I__5606\ : Span4Mux_v
    port map (
            O => \N__23705\,
            I => \N__23590\
        );

    \I__5605\ : Span4Mux_h
    port map (
            O => \N__23702\,
            I => \N__23590\
        );

    \I__5604\ : Span4Mux_h
    port map (
            O => \N__23697\,
            I => \N__23590\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__23694\,
            I => \N__23590\
        );

    \I__5602\ : Span4Mux_h
    port map (
            O => \N__23691\,
            I => \N__23587\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__23688\,
            I => \N__23584\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__23685\,
            I => \N__23579\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__23682\,
            I => \N__23579\
        );

    \I__5598\ : ClkMux
    port map (
            O => \N__23681\,
            I => \N__23576\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__23678\,
            I => \N__23573\
        );

    \I__5596\ : Span4Mux_v
    port map (
            O => \N__23675\,
            I => \N__23568\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__23672\,
            I => \N__23568\
        );

    \I__5594\ : Span4Mux_v
    port map (
            O => \N__23665\,
            I => \N__23559\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__23660\,
            I => \N__23559\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23559\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__23654\,
            I => \N__23559\
        );

    \I__5590\ : ClkMux
    port map (
            O => \N__23653\,
            I => \N__23556\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__23650\,
            I => \N__23553\
        );

    \I__5588\ : Span4Mux_s1_v
    port map (
            O => \N__23647\,
            I => \N__23550\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__23644\,
            I => \N__23547\
        );

    \I__5586\ : ClkMux
    port map (
            O => \N__23643\,
            I => \N__23544\
        );

    \I__5585\ : Span4Mux_v
    port map (
            O => \N__23640\,
            I => \N__23541\
        );

    \I__5584\ : Span4Mux_v
    port map (
            O => \N__23637\,
            I => \N__23538\
        );

    \I__5583\ : Sp12to4
    port map (
            O => \N__23634\,
            I => \N__23533\
        );

    \I__5582\ : Sp12to4
    port map (
            O => \N__23631\,
            I => \N__23533\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__23628\,
            I => \N__23530\
        );

    \I__5580\ : Span4Mux_v
    port map (
            O => \N__23625\,
            I => \N__23527\
        );

    \I__5579\ : Span4Mux_v
    port map (
            O => \N__23620\,
            I => \N__23522\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__23617\,
            I => \N__23522\
        );

    \I__5577\ : ClkMux
    port map (
            O => \N__23616\,
            I => \N__23519\
        );

    \I__5576\ : Span4Mux_h
    port map (
            O => \N__23611\,
            I => \N__23516\
        );

    \I__5575\ : Span4Mux_v
    port map (
            O => \N__23604\,
            I => \N__23509\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__23599\,
            I => \N__23509\
        );

    \I__5573\ : Span4Mux_h
    port map (
            O => \N__23590\,
            I => \N__23509\
        );

    \I__5572\ : Span4Mux_v
    port map (
            O => \N__23587\,
            I => \N__23504\
        );

    \I__5571\ : Span4Mux_h
    port map (
            O => \N__23584\,
            I => \N__23504\
        );

    \I__5570\ : Span4Mux_v
    port map (
            O => \N__23579\,
            I => \N__23499\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__23576\,
            I => \N__23499\
        );

    \I__5568\ : Span4Mux_h
    port map (
            O => \N__23573\,
            I => \N__23490\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__23568\,
            I => \N__23490\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__23559\,
            I => \N__23490\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__23556\,
            I => \N__23490\
        );

    \I__5564\ : Span4Mux_v
    port map (
            O => \N__23553\,
            I => \N__23483\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__23550\,
            I => \N__23483\
        );

    \I__5562\ : Span4Mux_h
    port map (
            O => \N__23547\,
            I => \N__23483\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__23544\,
            I => \N__23480\
        );

    \I__5560\ : Span4Mux_v
    port map (
            O => \N__23541\,
            I => \N__23477\
        );

    \I__5559\ : Span4Mux_v
    port map (
            O => \N__23538\,
            I => \N__23474\
        );

    \I__5558\ : Span12Mux_h
    port map (
            O => \N__23533\,
            I => \N__23469\
        );

    \I__5557\ : Span12Mux_h
    port map (
            O => \N__23530\,
            I => \N__23469\
        );

    \I__5556\ : Sp12to4
    port map (
            O => \N__23527\,
            I => \N__23464\
        );

    \I__5555\ : Sp12to4
    port map (
            O => \N__23522\,
            I => \N__23464\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__23519\,
            I => \N__23461\
        );

    \I__5553\ : Span4Mux_v
    port map (
            O => \N__23516\,
            I => \N__23458\
        );

    \I__5552\ : Span4Mux_v
    port map (
            O => \N__23509\,
            I => \N__23455\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__23504\,
            I => \N__23452\
        );

    \I__5550\ : Span4Mux_h
    port map (
            O => \N__23499\,
            I => \N__23449\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__23490\,
            I => \N__23446\
        );

    \I__5548\ : Span4Mux_h
    port map (
            O => \N__23483\,
            I => \N__23443\
        );

    \I__5547\ : Span4Mux_h
    port map (
            O => \N__23480\,
            I => \N__23440\
        );

    \I__5546\ : IoSpan4Mux
    port map (
            O => \N__23477\,
            I => \N__23437\
        );

    \I__5545\ : IoSpan4Mux
    port map (
            O => \N__23474\,
            I => \N__23434\
        );

    \I__5544\ : Span12Mux_v
    port map (
            O => \N__23469\,
            I => \N__23425\
        );

    \I__5543\ : Span12Mux_h
    port map (
            O => \N__23464\,
            I => \N__23425\
        );

    \I__5542\ : Span12Mux_h
    port map (
            O => \N__23461\,
            I => \N__23425\
        );

    \I__5541\ : Sp12to4
    port map (
            O => \N__23458\,
            I => \N__23425\
        );

    \I__5540\ : Span4Mux_v
    port map (
            O => \N__23455\,
            I => \N__23422\
        );

    \I__5539\ : Span4Mux_h
    port map (
            O => \N__23452\,
            I => \N__23415\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__23449\,
            I => \N__23415\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__23446\,
            I => \N__23415\
        );

    \I__5536\ : Span4Mux_h
    port map (
            O => \N__23443\,
            I => \N__23410\
        );

    \I__5535\ : Span4Mux_h
    port map (
            O => \N__23440\,
            I => \N__23410\
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__23437\,
            I => \ADV_CLK_c\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__23434\,
            I => \ADV_CLK_c\
        );

    \I__5532\ : Odrv12
    port map (
            O => \N__23425\,
            I => \ADV_CLK_c\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__23422\,
            I => \ADV_CLK_c\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__23415\,
            I => \ADV_CLK_c\
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__23410\,
            I => \ADV_CLK_c\
        );

    \I__5528\ : CEMux
    port map (
            O => \N__23397\,
            I => \N__23392\
        );

    \I__5527\ : CEMux
    port map (
            O => \N__23396\,
            I => \N__23388\
        );

    \I__5526\ : CEMux
    port map (
            O => \N__23395\,
            I => \N__23384\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__23392\,
            I => \N__23381\
        );

    \I__5524\ : CEMux
    port map (
            O => \N__23391\,
            I => \N__23378\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__23388\,
            I => \N__23375\
        );

    \I__5522\ : CEMux
    port map (
            O => \N__23387\,
            I => \N__23372\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__23384\,
            I => \N__23369\
        );

    \I__5520\ : Span4Mux_v
    port map (
            O => \N__23381\,
            I => \N__23364\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23364\
        );

    \I__5518\ : Span4Mux_h
    port map (
            O => \N__23375\,
            I => \N__23359\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__23372\,
            I => \N__23359\
        );

    \I__5516\ : Span4Mux_h
    port map (
            O => \N__23369\,
            I => \N__23356\
        );

    \I__5515\ : Span4Mux_h
    port map (
            O => \N__23364\,
            I => \N__23351\
        );

    \I__5514\ : Span4Mux_h
    port map (
            O => \N__23359\,
            I => \N__23351\
        );

    \I__5513\ : Odrv4
    port map (
            O => \N__23356\,
            I => \transmit_module.n2206\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__23351\,
            I => \transmit_module.n2206\
        );

    \I__5511\ : IoInMux
    port map (
            O => \N__23346\,
            I => \N__23343\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__23343\,
            I => \N__23340\
        );

    \I__5509\ : IoSpan4Mux
    port map (
            O => \N__23340\,
            I => \N__23337\
        );

    \I__5508\ : Span4Mux_s1_h
    port map (
            O => \N__23337\,
            I => \N__23328\
        );

    \I__5507\ : SRMux
    port map (
            O => \N__23336\,
            I => \N__23320\
        );

    \I__5506\ : SRMux
    port map (
            O => \N__23335\,
            I => \N__23317\
        );

    \I__5505\ : SRMux
    port map (
            O => \N__23334\,
            I => \N__23314\
        );

    \I__5504\ : SRMux
    port map (
            O => \N__23333\,
            I => \N__23311\
        );

    \I__5503\ : SRMux
    port map (
            O => \N__23332\,
            I => \N__23307\
        );

    \I__5502\ : SRMux
    port map (
            O => \N__23331\,
            I => \N__23304\
        );

    \I__5501\ : Span4Mux_h
    port map (
            O => \N__23328\,
            I => \N__23293\
        );

    \I__5500\ : SRMux
    port map (
            O => \N__23327\,
            I => \N__23290\
        );

    \I__5499\ : SRMux
    port map (
            O => \N__23326\,
            I => \N__23287\
        );

    \I__5498\ : SRMux
    port map (
            O => \N__23325\,
            I => \N__23277\
        );

    \I__5497\ : SRMux
    port map (
            O => \N__23324\,
            I => \N__23271\
        );

    \I__5496\ : SRMux
    port map (
            O => \N__23323\,
            I => \N__23268\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__23320\,
            I => \N__23265\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__23317\,
            I => \N__23262\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__23314\,
            I => \N__23257\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__23311\,
            I => \N__23257\
        );

    \I__5491\ : SRMux
    port map (
            O => \N__23310\,
            I => \N__23254\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__23307\,
            I => \N__23247\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__23304\,
            I => \N__23247\
        );

    \I__5488\ : SRMux
    port map (
            O => \N__23303\,
            I => \N__23244\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__23302\,
            I => \N__23235\
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__23301\,
            I => \N__23230\
        );

    \I__5485\ : SRMux
    port map (
            O => \N__23300\,
            I => \N__23225\
        );

    \I__5484\ : CascadeMux
    port map (
            O => \N__23299\,
            I => \N__23220\
        );

    \I__5483\ : CascadeMux
    port map (
            O => \N__23298\,
            I => \N__23217\
        );

    \I__5482\ : CascadeMux
    port map (
            O => \N__23297\,
            I => \N__23214\
        );

    \I__5481\ : SRMux
    port map (
            O => \N__23296\,
            I => \N__23209\
        );

    \I__5480\ : Span4Mux_h
    port map (
            O => \N__23293\,
            I => \N__23202\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__23290\,
            I => \N__23202\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__23287\,
            I => \N__23202\
        );

    \I__5477\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23199\
        );

    \I__5476\ : SRMux
    port map (
            O => \N__23285\,
            I => \N__23193\
        );

    \I__5475\ : SRMux
    port map (
            O => \N__23284\,
            I => \N__23190\
        );

    \I__5474\ : SRMux
    port map (
            O => \N__23283\,
            I => \N__23187\
        );

    \I__5473\ : SRMux
    port map (
            O => \N__23282\,
            I => \N__23184\
        );

    \I__5472\ : SRMux
    port map (
            O => \N__23281\,
            I => \N__23181\
        );

    \I__5471\ : SRMux
    port map (
            O => \N__23280\,
            I => \N__23178\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__23277\,
            I => \N__23175\
        );

    \I__5469\ : SRMux
    port map (
            O => \N__23276\,
            I => \N__23171\
        );

    \I__5468\ : SRMux
    port map (
            O => \N__23275\,
            I => \N__23168\
        );

    \I__5467\ : SRMux
    port map (
            O => \N__23274\,
            I => \N__23165\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__23271\,
            I => \N__23158\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__23268\,
            I => \N__23158\
        );

    \I__5464\ : Span4Mux_v
    port map (
            O => \N__23265\,
            I => \N__23158\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__23262\,
            I => \N__23151\
        );

    \I__5462\ : Span4Mux_v
    port map (
            O => \N__23257\,
            I => \N__23151\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__23254\,
            I => \N__23151\
        );

    \I__5460\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23148\
        );

    \I__5459\ : SRMux
    port map (
            O => \N__23252\,
            I => \N__23145\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__23247\,
            I => \N__23135\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__23244\,
            I => \N__23135\
        );

    \I__5456\ : SRMux
    port map (
            O => \N__23243\,
            I => \N__23132\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__23242\,
            I => \N__23129\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__23241\,
            I => \N__23126\
        );

    \I__5453\ : CascadeMux
    port map (
            O => \N__23240\,
            I => \N__23122\
        );

    \I__5452\ : SRMux
    port map (
            O => \N__23239\,
            I => \N__23116\
        );

    \I__5451\ : SRMux
    port map (
            O => \N__23238\,
            I => \N__23111\
        );

    \I__5450\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23111\
        );

    \I__5449\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23108\
        );

    \I__5448\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23101\
        );

    \I__5447\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23101\
        );

    \I__5446\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23101\
        );

    \I__5445\ : SRMux
    port map (
            O => \N__23228\,
            I => \N__23098\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__23225\,
            I => \N__23095\
        );

    \I__5443\ : SRMux
    port map (
            O => \N__23224\,
            I => \N__23092\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__23223\,
            I => \N__23088\
        );

    \I__5441\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23083\
        );

    \I__5440\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23083\
        );

    \I__5439\ : InMux
    port map (
            O => \N__23214\,
            I => \N__23080\
        );

    \I__5438\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23075\
        );

    \I__5437\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23075\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__23209\,
            I => \N__23068\
        );

    \I__5435\ : Span4Mux_v
    port map (
            O => \N__23202\,
            I => \N__23068\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__23199\,
            I => \N__23068\
        );

    \I__5433\ : SRMux
    port map (
            O => \N__23198\,
            I => \N__23065\
        );

    \I__5432\ : SRMux
    port map (
            O => \N__23197\,
            I => \N__23062\
        );

    \I__5431\ : SRMux
    port map (
            O => \N__23196\,
            I => \N__23059\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__23193\,
            I => \N__23056\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__23190\,
            I => \N__23053\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__23187\,
            I => \N__23050\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__23184\,
            I => \N__23047\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__23181\,
            I => \N__23040\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__23178\,
            I => \N__23040\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__23175\,
            I => \N__23040\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__23174\,
            I => \N__23037\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__23171\,
            I => \N__23034\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23031\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__23165\,
            I => \N__23026\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__23158\,
            I => \N__23026\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__23151\,
            I => \N__23019\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__23148\,
            I => \N__23019\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__23145\,
            I => \N__23016\
        );

    \I__5415\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23007\
        );

    \I__5414\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23007\
        );

    \I__5413\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23007\
        );

    \I__5412\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23007\
        );

    \I__5411\ : SRMux
    port map (
            O => \N__23140\,
            I => \N__23004\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__23135\,
            I => \N__23001\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__23132\,
            I => \N__22998\
        );

    \I__5408\ : InMux
    port map (
            O => \N__23129\,
            I => \N__22991\
        );

    \I__5407\ : InMux
    port map (
            O => \N__23126\,
            I => \N__22991\
        );

    \I__5406\ : InMux
    port map (
            O => \N__23125\,
            I => \N__22991\
        );

    \I__5405\ : InMux
    port map (
            O => \N__23122\,
            I => \N__22982\
        );

    \I__5404\ : InMux
    port map (
            O => \N__23121\,
            I => \N__22982\
        );

    \I__5403\ : InMux
    port map (
            O => \N__23120\,
            I => \N__22982\
        );

    \I__5402\ : InMux
    port map (
            O => \N__23119\,
            I => \N__22982\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__23116\,
            I => \N__22973\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__23111\,
            I => \N__22973\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__23108\,
            I => \N__22973\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__22973\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__23098\,
            I => \N__22970\
        );

    \I__5396\ : Span4Mux_h
    port map (
            O => \N__23095\,
            I => \N__22965\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__23092\,
            I => \N__22965\
        );

    \I__5394\ : InMux
    port map (
            O => \N__23091\,
            I => \N__22960\
        );

    \I__5393\ : InMux
    port map (
            O => \N__23088\,
            I => \N__22960\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__23083\,
            I => \N__22951\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N__22951\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__23075\,
            I => \N__22951\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__23068\,
            I => \N__22951\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__22946\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__23062\,
            I => \N__22946\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__23059\,
            I => \N__22941\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__23056\,
            I => \N__22941\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__23053\,
            I => \N__22932\
        );

    \I__5383\ : Span4Mux_v
    port map (
            O => \N__23050\,
            I => \N__22932\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__23047\,
            I => \N__22932\
        );

    \I__5381\ : Span4Mux_h
    port map (
            O => \N__23040\,
            I => \N__22932\
        );

    \I__5380\ : InMux
    port map (
            O => \N__23037\,
            I => \N__22929\
        );

    \I__5379\ : Span4Mux_v
    port map (
            O => \N__23034\,
            I => \N__22922\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__23031\,
            I => \N__22922\
        );

    \I__5377\ : Span4Mux_h
    port map (
            O => \N__23026\,
            I => \N__22922\
        );

    \I__5376\ : InMux
    port map (
            O => \N__23025\,
            I => \N__22917\
        );

    \I__5375\ : InMux
    port map (
            O => \N__23024\,
            I => \N__22917\
        );

    \I__5374\ : Span4Mux_h
    port map (
            O => \N__23019\,
            I => \N__22910\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__23016\,
            I => \N__22910\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__23007\,
            I => \N__22910\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__23004\,
            I => \N__22897\
        );

    \I__5370\ : Span4Mux_h
    port map (
            O => \N__23001\,
            I => \N__22897\
        );

    \I__5369\ : Span4Mux_h
    port map (
            O => \N__22998\,
            I => \N__22897\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22897\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__22982\,
            I => \N__22897\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__22973\,
            I => \N__22897\
        );

    \I__5365\ : Span4Mux_h
    port map (
            O => \N__22970\,
            I => \N__22888\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__22965\,
            I => \N__22888\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__22960\,
            I => \N__22888\
        );

    \I__5362\ : Span4Mux_v
    port map (
            O => \N__22951\,
            I => \N__22888\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__22946\,
            I => \ADV_VSYNC_c\
        );

    \I__5360\ : Odrv4
    port map (
            O => \N__22941\,
            I => \ADV_VSYNC_c\
        );

    \I__5359\ : Odrv4
    port map (
            O => \N__22932\,
            I => \ADV_VSYNC_c\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__22929\,
            I => \ADV_VSYNC_c\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__22922\,
            I => \ADV_VSYNC_c\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__22917\,
            I => \ADV_VSYNC_c\
        );

    \I__5355\ : Odrv4
    port map (
            O => \N__22910\,
            I => \ADV_VSYNC_c\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__22897\,
            I => \ADV_VSYNC_c\
        );

    \I__5353\ : Odrv4
    port map (
            O => \N__22888\,
            I => \ADV_VSYNC_c\
        );

    \I__5352\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22866\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__5350\ : Span12Mux_h
    port map (
            O => \N__22863\,
            I => \N__22860\
        );

    \I__5349\ : Span12Mux_v
    port map (
            O => \N__22860\,
            I => \N__22857\
        );

    \I__5348\ : Odrv12
    port map (
            O => \N__22857\,
            I => \line_buffer.n589\
        );

    \I__5347\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22851\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__22851\,
            I => \N__22848\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__22848\,
            I => \N__22845\
        );

    \I__5344\ : Sp12to4
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__5343\ : Odrv12
    port map (
            O => \N__22842\,
            I => \line_buffer.n597\
        );

    \I__5342\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__22836\,
            I => \line_buffer.n3534\
        );

    \I__5340\ : InMux
    port map (
            O => \N__22833\,
            I => \N__22822\
        );

    \I__5339\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22818\
        );

    \I__5338\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22815\
        );

    \I__5337\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22812\
        );

    \I__5336\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22809\
        );

    \I__5335\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22804\
        );

    \I__5334\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22799\
        );

    \I__5333\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22799\
        );

    \I__5332\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22795\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__22822\,
            I => \N__22792\
        );

    \I__5330\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22789\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__22818\,
            I => \N__22786\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__22815\,
            I => \N__22783\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__22812\,
            I => \N__22778\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__22809\,
            I => \N__22778\
        );

    \I__5325\ : InMux
    port map (
            O => \N__22808\,
            I => \N__22775\
        );

    \I__5324\ : InMux
    port map (
            O => \N__22807\,
            I => \N__22772\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__22804\,
            I => \N__22764\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__22799\,
            I => \N__22760\
        );

    \I__5321\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22756\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__22795\,
            I => \N__22748\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__22792\,
            I => \N__22748\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__22789\,
            I => \N__22745\
        );

    \I__5317\ : Span4Mux_h
    port map (
            O => \N__22786\,
            I => \N__22736\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__22783\,
            I => \N__22736\
        );

    \I__5315\ : Span4Mux_v
    port map (
            O => \N__22778\,
            I => \N__22736\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__22775\,
            I => \N__22736\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22733\
        );

    \I__5312\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22730\
        );

    \I__5311\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22727\
        );

    \I__5310\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22724\
        );

    \I__5309\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22720\
        );

    \I__5308\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22717\
        );

    \I__5307\ : Span4Mux_v
    port map (
            O => \N__22764\,
            I => \N__22714\
        );

    \I__5306\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22711\
        );

    \I__5305\ : Span4Mux_h
    port map (
            O => \N__22760\,
            I => \N__22708\
        );

    \I__5304\ : InMux
    port map (
            O => \N__22759\,
            I => \N__22704\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__22756\,
            I => \N__22701\
        );

    \I__5302\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22698\
        );

    \I__5301\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22695\
        );

    \I__5300\ : InMux
    port map (
            O => \N__22753\,
            I => \N__22692\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__22748\,
            I => \N__22689\
        );

    \I__5298\ : Span4Mux_v
    port map (
            O => \N__22745\,
            I => \N__22684\
        );

    \I__5297\ : Span4Mux_v
    port map (
            O => \N__22736\,
            I => \N__22684\
        );

    \I__5296\ : Span4Mux_v
    port map (
            O => \N__22733\,
            I => \N__22675\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22675\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__22727\,
            I => \N__22675\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__22724\,
            I => \N__22675\
        );

    \I__5292\ : InMux
    port map (
            O => \N__22723\,
            I => \N__22672\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__22720\,
            I => \N__22669\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__22717\,
            I => \N__22662\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__22714\,
            I => \N__22662\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__22711\,
            I => \N__22662\
        );

    \I__5287\ : Span4Mux_h
    port map (
            O => \N__22708\,
            I => \N__22659\
        );

    \I__5286\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22656\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22651\
        );

    \I__5284\ : Span4Mux_h
    port map (
            O => \N__22701\,
            I => \N__22651\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__22698\,
            I => \N__22648\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__22695\,
            I => \N__22643\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__22692\,
            I => \N__22643\
        );

    \I__5280\ : Span4Mux_v
    port map (
            O => \N__22689\,
            I => \N__22634\
        );

    \I__5279\ : Span4Mux_h
    port map (
            O => \N__22684\,
            I => \N__22634\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__22675\,
            I => \N__22634\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__22672\,
            I => \N__22634\
        );

    \I__5276\ : Span4Mux_h
    port map (
            O => \N__22669\,
            I => \N__22620\
        );

    \I__5275\ : Span4Mux_h
    port map (
            O => \N__22662\,
            I => \N__22620\
        );

    \I__5274\ : Span4Mux_v
    port map (
            O => \N__22659\,
            I => \N__22620\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22620\
        );

    \I__5272\ : Span4Mux_v
    port map (
            O => \N__22651\,
            I => \N__22620\
        );

    \I__5271\ : Span4Mux_v
    port map (
            O => \N__22648\,
            I => \N__22620\
        );

    \I__5270\ : Span4Mux_v
    port map (
            O => \N__22643\,
            I => \N__22617\
        );

    \I__5269\ : Span4Mux_h
    port map (
            O => \N__22634\,
            I => \N__22614\
        );

    \I__5268\ : InMux
    port map (
            O => \N__22633\,
            I => \N__22611\
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__22620\,
            I => \TX_ADDR_11\
        );

    \I__5266\ : Odrv4
    port map (
            O => \N__22617\,
            I => \TX_ADDR_11\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__22614\,
            I => \TX_ADDR_11\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__22611\,
            I => \TX_ADDR_11\
        );

    \I__5263\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22599\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__22599\,
            I => \N__22596\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__22596\,
            I => \N__22593\
        );

    \I__5260\ : Sp12to4
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__5259\ : Odrv12
    port map (
            O => \N__22590\,
            I => \line_buffer.n535\
        );

    \I__5258\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__22581\,
            I => \N__22578\
        );

    \I__5255\ : Span4Mux_v
    port map (
            O => \N__22578\,
            I => \N__22575\
        );

    \I__5254\ : Sp12to4
    port map (
            O => \N__22575\,
            I => \N__22572\
        );

    \I__5253\ : Span12Mux_v
    port map (
            O => \N__22572\,
            I => \N__22569\
        );

    \I__5252\ : Odrv12
    port map (
            O => \N__22569\,
            I => \line_buffer.n527\
        );

    \I__5251\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22563\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__22563\,
            I => \line_buffer.n3539\
        );

    \I__5249\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22557\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__22557\,
            I => \N__22554\
        );

    \I__5247\ : Span4Mux_v
    port map (
            O => \N__22554\,
            I => \N__22551\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__22551\,
            I => \TX_DATA_4\
        );

    \I__5245\ : IoInMux
    port map (
            O => \N__22548\,
            I => \N__22545\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__5243\ : IoSpan4Mux
    port map (
            O => \N__22542\,
            I => \N__22539\
        );

    \I__5242\ : IoSpan4Mux
    port map (
            O => \N__22539\,
            I => \N__22535\
        );

    \I__5241\ : IoInMux
    port map (
            O => \N__22538\,
            I => \N__22532\
        );

    \I__5240\ : IoSpan4Mux
    port map (
            O => \N__22535\,
            I => \N__22526\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__22532\,
            I => \N__22526\
        );

    \I__5238\ : IoInMux
    port map (
            O => \N__22531\,
            I => \N__22523\
        );

    \I__5237\ : IoSpan4Mux
    port map (
            O => \N__22526\,
            I => \N__22520\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__22523\,
            I => \N__22517\
        );

    \I__5235\ : Span4Mux_s2_h
    port map (
            O => \N__22520\,
            I => \N__22514\
        );

    \I__5234\ : Span4Mux_s1_v
    port map (
            O => \N__22517\,
            I => \N__22511\
        );

    \I__5233\ : Sp12to4
    port map (
            O => \N__22514\,
            I => \N__22508\
        );

    \I__5232\ : Sp12to4
    port map (
            O => \N__22511\,
            I => \N__22505\
        );

    \I__5231\ : Span12Mux_h
    port map (
            O => \N__22508\,
            I => \N__22502\
        );

    \I__5230\ : Span12Mux_h
    port map (
            O => \N__22505\,
            I => \N__22499\
        );

    \I__5229\ : Odrv12
    port map (
            O => \N__22502\,
            I => n1814
        );

    \I__5228\ : Odrv12
    port map (
            O => \N__22499\,
            I => n1814
        );

    \I__5227\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22491\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__22491\,
            I => \TX_DATA_6\
        );

    \I__5225\ : IoInMux
    port map (
            O => \N__22488\,
            I => \N__22485\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__22485\,
            I => \N__22482\
        );

    \I__5223\ : IoSpan4Mux
    port map (
            O => \N__22482\,
            I => \N__22478\
        );

    \I__5222\ : IoInMux
    port map (
            O => \N__22481\,
            I => \N__22474\
        );

    \I__5221\ : Span4Mux_s1_h
    port map (
            O => \N__22478\,
            I => \N__22471\
        );

    \I__5220\ : IoInMux
    port map (
            O => \N__22477\,
            I => \N__22468\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__22474\,
            I => \N__22465\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__22471\,
            I => \N__22462\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__22468\,
            I => \N__22459\
        );

    \I__5216\ : Span4Mux_s3_v
    port map (
            O => \N__22465\,
            I => \N__22456\
        );

    \I__5215\ : Span4Mux_h
    port map (
            O => \N__22462\,
            I => \N__22451\
        );

    \I__5214\ : Span4Mux_s3_v
    port map (
            O => \N__22459\,
            I => \N__22451\
        );

    \I__5213\ : Span4Mux_v
    port map (
            O => \N__22456\,
            I => \N__22448\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__22451\,
            I => \N__22445\
        );

    \I__5211\ : Sp12to4
    port map (
            O => \N__22448\,
            I => \N__22442\
        );

    \I__5210\ : Sp12to4
    port map (
            O => \N__22445\,
            I => \N__22439\
        );

    \I__5209\ : Span12Mux_h
    port map (
            O => \N__22442\,
            I => \N__22434\
        );

    \I__5208\ : Span12Mux_h
    port map (
            O => \N__22439\,
            I => \N__22434\
        );

    \I__5207\ : Odrv12
    port map (
            O => \N__22434\,
            I => n1812
        );

    \I__5206\ : SRMux
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__22428\,
            I => \N__22421\
        );

    \I__5204\ : SRMux
    port map (
            O => \N__22427\,
            I => \N__22418\
        );

    \I__5203\ : SRMux
    port map (
            O => \N__22426\,
            I => \N__22415\
        );

    \I__5202\ : SRMux
    port map (
            O => \N__22425\,
            I => \N__22411\
        );

    \I__5201\ : SRMux
    port map (
            O => \N__22424\,
            I => \N__22408\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__22421\,
            I => \N__22401\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__22418\,
            I => \N__22401\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__22415\,
            I => \N__22401\
        );

    \I__5197\ : SRMux
    port map (
            O => \N__22414\,
            I => \N__22398\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__22411\,
            I => \N__22394\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__22408\,
            I => \N__22391\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__22401\,
            I => \N__22386\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__22398\,
            I => \N__22386\
        );

    \I__5192\ : SRMux
    port map (
            O => \N__22397\,
            I => \N__22383\
        );

    \I__5191\ : Span4Mux_h
    port map (
            O => \N__22394\,
            I => \N__22380\
        );

    \I__5190\ : Span4Mux_v
    port map (
            O => \N__22391\,
            I => \N__22377\
        );

    \I__5189\ : Span4Mux_h
    port map (
            O => \N__22386\,
            I => \N__22374\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22371\
        );

    \I__5187\ : Odrv4
    port map (
            O => \N__22380\,
            I => \transmit_module.n2385\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__22377\,
            I => \transmit_module.n2385\
        );

    \I__5185\ : Odrv4
    port map (
            O => \N__22374\,
            I => \transmit_module.n2385\
        );

    \I__5184\ : Odrv12
    port map (
            O => \N__22371\,
            I => \transmit_module.n2385\
        );

    \I__5183\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22359\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__22359\,
            I => \N__22356\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__22356\,
            I => \N__22353\
        );

    \I__5180\ : Span4Mux_h
    port map (
            O => \N__22353\,
            I => \N__22350\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__22350\,
            I => \line_buffer.n470\
        );

    \I__5178\ : InMux
    port map (
            O => \N__22347\,
            I => \N__22344\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__5176\ : Span12Mux_v
    port map (
            O => \N__22341\,
            I => \N__22338\
        );

    \I__5175\ : Odrv12
    port map (
            O => \N__22338\,
            I => \line_buffer.n462\
        );

    \I__5174\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22332\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__22332\,
            I => \N__22329\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__22329\,
            I => \line_buffer.n3572\
        );

    \I__5171\ : SRMux
    port map (
            O => \N__22326\,
            I => \N__22323\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22319\
        );

    \I__5169\ : SRMux
    port map (
            O => \N__22322\,
            I => \N__22316\
        );

    \I__5168\ : Span4Mux_h
    port map (
            O => \N__22319\,
            I => \N__22310\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22310\
        );

    \I__5166\ : SRMux
    port map (
            O => \N__22315\,
            I => \N__22307\
        );

    \I__5165\ : Span4Mux_v
    port map (
            O => \N__22310\,
            I => \N__22301\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22301\
        );

    \I__5163\ : SRMux
    port map (
            O => \N__22306\,
            I => \N__22298\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__22301\,
            I => \N__22292\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22292\
        );

    \I__5160\ : SRMux
    port map (
            O => \N__22297\,
            I => \N__22289\
        );

    \I__5159\ : Span4Mux_v
    port map (
            O => \N__22292\,
            I => \N__22283\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__22289\,
            I => \N__22283\
        );

    \I__5157\ : SRMux
    port map (
            O => \N__22288\,
            I => \N__22280\
        );

    \I__5156\ : Span4Mux_h
    port map (
            O => \N__22283\,
            I => \N__22274\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__22280\,
            I => \N__22274\
        );

    \I__5154\ : SRMux
    port map (
            O => \N__22279\,
            I => \N__22271\
        );

    \I__5153\ : Span4Mux_v
    port map (
            O => \N__22274\,
            I => \N__22264\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__22271\,
            I => \N__22264\
        );

    \I__5151\ : SRMux
    port map (
            O => \N__22270\,
            I => \N__22261\
        );

    \I__5150\ : SRMux
    port map (
            O => \N__22269\,
            I => \N__22257\
        );

    \I__5149\ : Span4Mux_h
    port map (
            O => \N__22264\,
            I => \N__22250\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22250\
        );

    \I__5147\ : SRMux
    port map (
            O => \N__22260\,
            I => \N__22247\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__22257\,
            I => \N__22243\
        );

    \I__5145\ : SRMux
    port map (
            O => \N__22256\,
            I => \N__22240\
        );

    \I__5144\ : SRMux
    port map (
            O => \N__22255\,
            I => \N__22237\
        );

    \I__5143\ : Span4Mux_v
    port map (
            O => \N__22250\,
            I => \N__22230\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__22247\,
            I => \N__22230\
        );

    \I__5141\ : SRMux
    port map (
            O => \N__22246\,
            I => \N__22227\
        );

    \I__5140\ : Span4Mux_s1_v
    port map (
            O => \N__22243\,
            I => \N__22219\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__22240\,
            I => \N__22219\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22219\
        );

    \I__5137\ : SRMux
    port map (
            O => \N__22236\,
            I => \N__22216\
        );

    \I__5136\ : SRMux
    port map (
            O => \N__22235\,
            I => \N__22213\
        );

    \I__5135\ : Span4Mux_h
    port map (
            O => \N__22230\,
            I => \N__22206\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22206\
        );

    \I__5133\ : SRMux
    port map (
            O => \N__22226\,
            I => \N__22203\
        );

    \I__5132\ : Span4Mux_v
    port map (
            O => \N__22219\,
            I => \N__22195\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__22216\,
            I => \N__22195\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__22213\,
            I => \N__22195\
        );

    \I__5129\ : SRMux
    port map (
            O => \N__22212\,
            I => \N__22192\
        );

    \I__5128\ : SRMux
    port map (
            O => \N__22211\,
            I => \N__22189\
        );

    \I__5127\ : Span4Mux_v
    port map (
            O => \N__22206\,
            I => \N__22182\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22182\
        );

    \I__5125\ : SRMux
    port map (
            O => \N__22202\,
            I => \N__22179\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__22195\,
            I => \N__22171\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__22192\,
            I => \N__22171\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__22189\,
            I => \N__22171\
        );

    \I__5121\ : SRMux
    port map (
            O => \N__22188\,
            I => \N__22168\
        );

    \I__5120\ : SRMux
    port map (
            O => \N__22187\,
            I => \N__22165\
        );

    \I__5119\ : Span4Mux_h
    port map (
            O => \N__22182\,
            I => \N__22158\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__22179\,
            I => \N__22158\
        );

    \I__5117\ : SRMux
    port map (
            O => \N__22178\,
            I => \N__22155\
        );

    \I__5116\ : Span4Mux_v
    port map (
            O => \N__22171\,
            I => \N__22146\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__22146\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__22165\,
            I => \N__22146\
        );

    \I__5113\ : SRMux
    port map (
            O => \N__22164\,
            I => \N__22143\
        );

    \I__5112\ : SRMux
    port map (
            O => \N__22163\,
            I => \N__22140\
        );

    \I__5111\ : Span4Mux_v
    port map (
            O => \N__22158\,
            I => \N__22133\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__22155\,
            I => \N__22133\
        );

    \I__5109\ : SRMux
    port map (
            O => \N__22154\,
            I => \N__22130\
        );

    \I__5108\ : SRMux
    port map (
            O => \N__22153\,
            I => \N__22127\
        );

    \I__5107\ : Span4Mux_v
    port map (
            O => \N__22146\,
            I => \N__22119\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__22143\,
            I => \N__22119\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__22140\,
            I => \N__22119\
        );

    \I__5104\ : SRMux
    port map (
            O => \N__22139\,
            I => \N__22116\
        );

    \I__5103\ : SRMux
    port map (
            O => \N__22138\,
            I => \N__22113\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__22133\,
            I => \N__22106\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__22130\,
            I => \N__22106\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__22127\,
            I => \N__22103\
        );

    \I__5099\ : SRMux
    port map (
            O => \N__22126\,
            I => \N__22100\
        );

    \I__5098\ : Span4Mux_v
    port map (
            O => \N__22119\,
            I => \N__22092\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__22116\,
            I => \N__22092\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__22113\,
            I => \N__22092\
        );

    \I__5095\ : SRMux
    port map (
            O => \N__22112\,
            I => \N__22089\
        );

    \I__5094\ : SRMux
    port map (
            O => \N__22111\,
            I => \N__22086\
        );

    \I__5093\ : Span4Mux_v
    port map (
            O => \N__22106\,
            I => \N__22079\
        );

    \I__5092\ : Span4Mux_s3_v
    port map (
            O => \N__22103\,
            I => \N__22079\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__22100\,
            I => \N__22079\
        );

    \I__5090\ : SRMux
    port map (
            O => \N__22099\,
            I => \N__22076\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__22092\,
            I => \N__22071\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22071\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__22086\,
            I => \N__22068\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__22079\,
            I => \N__22065\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__22076\,
            I => \N__22061\
        );

    \I__5084\ : Span4Mux_v
    port map (
            O => \N__22071\,
            I => \N__22055\
        );

    \I__5083\ : Span4Mux_s2_v
    port map (
            O => \N__22068\,
            I => \N__22055\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__22065\,
            I => \N__22052\
        );

    \I__5081\ : IoInMux
    port map (
            O => \N__22064\,
            I => \N__22049\
        );

    \I__5080\ : Span4Mux_h
    port map (
            O => \N__22061\,
            I => \N__22046\
        );

    \I__5079\ : IoInMux
    port map (
            O => \N__22060\,
            I => \N__22043\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__22055\,
            I => \N__22040\
        );

    \I__5077\ : Span4Mux_h
    port map (
            O => \N__22052\,
            I => \N__22031\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__22049\,
            I => \N__22031\
        );

    \I__5075\ : Span4Mux_h
    port map (
            O => \N__22046\,
            I => \N__22031\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__22043\,
            I => \N__22031\
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__22040\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__22031\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5071\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22023\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22020\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__22020\,
            I => \N__22017\
        );

    \I__5068\ : Span4Mux_v
    port map (
            O => \N__22017\,
            I => \N__22014\
        );

    \I__5067\ : Odrv4
    port map (
            O => \N__22014\,
            I => \TVP_VIDEO_c_9\
        );

    \I__5066\ : InMux
    port map (
            O => \N__22011\,
            I => \N__22008\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__22008\,
            I => \tvp_video_buffer.BUFFER_0_9\
        );

    \I__5064\ : InMux
    port map (
            O => \N__22005\,
            I => \N__22002\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__22002\,
            I => \tvp_video_buffer.BUFFER_1_9\
        );

    \I__5062\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21996\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__21996\,
            I => \N__21978\
        );

    \I__5060\ : ClkMux
    port map (
            O => \N__21995\,
            I => \N__21789\
        );

    \I__5059\ : ClkMux
    port map (
            O => \N__21994\,
            I => \N__21789\
        );

    \I__5058\ : ClkMux
    port map (
            O => \N__21993\,
            I => \N__21789\
        );

    \I__5057\ : ClkMux
    port map (
            O => \N__21992\,
            I => \N__21789\
        );

    \I__5056\ : ClkMux
    port map (
            O => \N__21991\,
            I => \N__21789\
        );

    \I__5055\ : ClkMux
    port map (
            O => \N__21990\,
            I => \N__21789\
        );

    \I__5054\ : ClkMux
    port map (
            O => \N__21989\,
            I => \N__21789\
        );

    \I__5053\ : ClkMux
    port map (
            O => \N__21988\,
            I => \N__21789\
        );

    \I__5052\ : ClkMux
    port map (
            O => \N__21987\,
            I => \N__21789\
        );

    \I__5051\ : ClkMux
    port map (
            O => \N__21986\,
            I => \N__21789\
        );

    \I__5050\ : ClkMux
    port map (
            O => \N__21985\,
            I => \N__21789\
        );

    \I__5049\ : ClkMux
    port map (
            O => \N__21984\,
            I => \N__21789\
        );

    \I__5048\ : ClkMux
    port map (
            O => \N__21983\,
            I => \N__21789\
        );

    \I__5047\ : ClkMux
    port map (
            O => \N__21982\,
            I => \N__21789\
        );

    \I__5046\ : ClkMux
    port map (
            O => \N__21981\,
            I => \N__21789\
        );

    \I__5045\ : Glb2LocalMux
    port map (
            O => \N__21978\,
            I => \N__21789\
        );

    \I__5044\ : ClkMux
    port map (
            O => \N__21977\,
            I => \N__21789\
        );

    \I__5043\ : ClkMux
    port map (
            O => \N__21976\,
            I => \N__21789\
        );

    \I__5042\ : ClkMux
    port map (
            O => \N__21975\,
            I => \N__21789\
        );

    \I__5041\ : ClkMux
    port map (
            O => \N__21974\,
            I => \N__21789\
        );

    \I__5040\ : ClkMux
    port map (
            O => \N__21973\,
            I => \N__21789\
        );

    \I__5039\ : ClkMux
    port map (
            O => \N__21972\,
            I => \N__21789\
        );

    \I__5038\ : ClkMux
    port map (
            O => \N__21971\,
            I => \N__21789\
        );

    \I__5037\ : ClkMux
    port map (
            O => \N__21970\,
            I => \N__21789\
        );

    \I__5036\ : ClkMux
    port map (
            O => \N__21969\,
            I => \N__21789\
        );

    \I__5035\ : ClkMux
    port map (
            O => \N__21968\,
            I => \N__21789\
        );

    \I__5034\ : ClkMux
    port map (
            O => \N__21967\,
            I => \N__21789\
        );

    \I__5033\ : ClkMux
    port map (
            O => \N__21966\,
            I => \N__21789\
        );

    \I__5032\ : ClkMux
    port map (
            O => \N__21965\,
            I => \N__21789\
        );

    \I__5031\ : ClkMux
    port map (
            O => \N__21964\,
            I => \N__21789\
        );

    \I__5030\ : ClkMux
    port map (
            O => \N__21963\,
            I => \N__21789\
        );

    \I__5029\ : ClkMux
    port map (
            O => \N__21962\,
            I => \N__21789\
        );

    \I__5028\ : ClkMux
    port map (
            O => \N__21961\,
            I => \N__21789\
        );

    \I__5027\ : ClkMux
    port map (
            O => \N__21960\,
            I => \N__21789\
        );

    \I__5026\ : ClkMux
    port map (
            O => \N__21959\,
            I => \N__21789\
        );

    \I__5025\ : ClkMux
    port map (
            O => \N__21958\,
            I => \N__21789\
        );

    \I__5024\ : ClkMux
    port map (
            O => \N__21957\,
            I => \N__21789\
        );

    \I__5023\ : ClkMux
    port map (
            O => \N__21956\,
            I => \N__21789\
        );

    \I__5022\ : ClkMux
    port map (
            O => \N__21955\,
            I => \N__21789\
        );

    \I__5021\ : ClkMux
    port map (
            O => \N__21954\,
            I => \N__21789\
        );

    \I__5020\ : ClkMux
    port map (
            O => \N__21953\,
            I => \N__21789\
        );

    \I__5019\ : ClkMux
    port map (
            O => \N__21952\,
            I => \N__21789\
        );

    \I__5018\ : ClkMux
    port map (
            O => \N__21951\,
            I => \N__21789\
        );

    \I__5017\ : ClkMux
    port map (
            O => \N__21950\,
            I => \N__21789\
        );

    \I__5016\ : ClkMux
    port map (
            O => \N__21949\,
            I => \N__21789\
        );

    \I__5015\ : ClkMux
    port map (
            O => \N__21948\,
            I => \N__21789\
        );

    \I__5014\ : ClkMux
    port map (
            O => \N__21947\,
            I => \N__21789\
        );

    \I__5013\ : ClkMux
    port map (
            O => \N__21946\,
            I => \N__21789\
        );

    \I__5012\ : ClkMux
    port map (
            O => \N__21945\,
            I => \N__21789\
        );

    \I__5011\ : ClkMux
    port map (
            O => \N__21944\,
            I => \N__21789\
        );

    \I__5010\ : ClkMux
    port map (
            O => \N__21943\,
            I => \N__21789\
        );

    \I__5009\ : ClkMux
    port map (
            O => \N__21942\,
            I => \N__21789\
        );

    \I__5008\ : ClkMux
    port map (
            O => \N__21941\,
            I => \N__21789\
        );

    \I__5007\ : ClkMux
    port map (
            O => \N__21940\,
            I => \N__21789\
        );

    \I__5006\ : ClkMux
    port map (
            O => \N__21939\,
            I => \N__21789\
        );

    \I__5005\ : ClkMux
    port map (
            O => \N__21938\,
            I => \N__21789\
        );

    \I__5004\ : ClkMux
    port map (
            O => \N__21937\,
            I => \N__21789\
        );

    \I__5003\ : ClkMux
    port map (
            O => \N__21936\,
            I => \N__21789\
        );

    \I__5002\ : ClkMux
    port map (
            O => \N__21935\,
            I => \N__21789\
        );

    \I__5001\ : ClkMux
    port map (
            O => \N__21934\,
            I => \N__21789\
        );

    \I__5000\ : ClkMux
    port map (
            O => \N__21933\,
            I => \N__21789\
        );

    \I__4999\ : ClkMux
    port map (
            O => \N__21932\,
            I => \N__21789\
        );

    \I__4998\ : ClkMux
    port map (
            O => \N__21931\,
            I => \N__21789\
        );

    \I__4997\ : ClkMux
    port map (
            O => \N__21930\,
            I => \N__21789\
        );

    \I__4996\ : ClkMux
    port map (
            O => \N__21929\,
            I => \N__21789\
        );

    \I__4995\ : ClkMux
    port map (
            O => \N__21928\,
            I => \N__21789\
        );

    \I__4994\ : ClkMux
    port map (
            O => \N__21927\,
            I => \N__21789\
        );

    \I__4993\ : ClkMux
    port map (
            O => \N__21926\,
            I => \N__21789\
        );

    \I__4992\ : GlobalMux
    port map (
            O => \N__21789\,
            I => \N__21786\
        );

    \I__4991\ : gio2CtrlBuf
    port map (
            O => \N__21786\,
            I => \DEBUG_c_3_c\
        );

    \I__4990\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__21780\,
            I => \N__21777\
        );

    \I__4988\ : Odrv4
    port map (
            O => \N__21777\,
            I => \transmit_module.Y_DELTA_PATTERN_88\
        );

    \I__4987\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21771\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21771\,
            I => \N__21768\
        );

    \I__4985\ : Span4Mux_v
    port map (
            O => \N__21768\,
            I => \N__21765\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__21765\,
            I => \transmit_module.Y_DELTA_PATTERN_84\
        );

    \I__4983\ : InMux
    port map (
            O => \N__21762\,
            I => \N__21759\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__21759\,
            I => \N__21756\
        );

    \I__4981\ : Sp12to4
    port map (
            O => \N__21756\,
            I => \N__21753\
        );

    \I__4980\ : Odrv12
    port map (
            O => \N__21753\,
            I => \line_buffer.n3533\
        );

    \I__4979\ : InMux
    port map (
            O => \N__21750\,
            I => \N__21747\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__21747\,
            I => \N__21744\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__21744\,
            I => \line_buffer.n3549\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__21741\,
            I => \line_buffer.n3611_cascade_\
        );

    \I__4975\ : InMux
    port map (
            O => \N__21738\,
            I => \N__21734\
        );

    \I__4974\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21731\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__21734\,
            I => \N__21728\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__21731\,
            I => \N__21721\
        );

    \I__4971\ : Span4Mux_v
    port map (
            O => \N__21728\,
            I => \N__21718\
        );

    \I__4970\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21715\
        );

    \I__4969\ : InMux
    port map (
            O => \N__21726\,
            I => \N__21711\
        );

    \I__4968\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21708\
        );

    \I__4967\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21705\
        );

    \I__4966\ : Span4Mux_v
    port map (
            O => \N__21721\,
            I => \N__21701\
        );

    \I__4965\ : Span4Mux_v
    port map (
            O => \N__21718\,
            I => \N__21696\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__21715\,
            I => \N__21696\
        );

    \I__4963\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21693\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__21711\,
            I => \N__21689\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__21708\,
            I => \N__21686\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__21705\,
            I => \N__21683\
        );

    \I__4959\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21680\
        );

    \I__4958\ : Span4Mux_v
    port map (
            O => \N__21701\,
            I => \N__21673\
        );

    \I__4957\ : Span4Mux_v
    port map (
            O => \N__21696\,
            I => \N__21673\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__21693\,
            I => \N__21673\
        );

    \I__4955\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21670\
        );

    \I__4954\ : Span12Mux_s5_v
    port map (
            O => \N__21689\,
            I => \N__21667\
        );

    \I__4953\ : Span12Mux_s6_v
    port map (
            O => \N__21686\,
            I => \N__21664\
        );

    \I__4952\ : Span12Mux_v
    port map (
            O => \N__21683\,
            I => \N__21659\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__21680\,
            I => \N__21659\
        );

    \I__4950\ : Span4Mux_v
    port map (
            O => \N__21673\,
            I => \N__21656\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__21670\,
            I => \N__21653\
        );

    \I__4948\ : Span12Mux_h
    port map (
            O => \N__21667\,
            I => \N__21650\
        );

    \I__4947\ : Span12Mux_h
    port map (
            O => \N__21664\,
            I => \N__21645\
        );

    \I__4946\ : Span12Mux_h
    port map (
            O => \N__21659\,
            I => \N__21645\
        );

    \I__4945\ : Sp12to4
    port map (
            O => \N__21656\,
            I => \N__21640\
        );

    \I__4944\ : Span12Mux_v
    port map (
            O => \N__21653\,
            I => \N__21640\
        );

    \I__4943\ : Odrv12
    port map (
            O => \N__21650\,
            I => \RX_DATA_4\
        );

    \I__4942\ : Odrv12
    port map (
            O => \N__21645\,
            I => \RX_DATA_4\
        );

    \I__4941\ : Odrv12
    port map (
            O => \N__21640\,
            I => \RX_DATA_4\
        );

    \I__4940\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__21630\,
            I => \tvp_video_buffer.BUFFER_1_6\
        );

    \I__4938\ : IoInMux
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__21624\,
            I => \N__21620\
        );

    \I__4936\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21617\
        );

    \I__4935\ : IoSpan4Mux
    port map (
            O => \N__21620\,
            I => \N__21614\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__21617\,
            I => \N__21611\
        );

    \I__4933\ : Span4Mux_s0_h
    port map (
            O => \N__21614\,
            I => \N__21608\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__21611\,
            I => \N__21605\
        );

    \I__4931\ : Sp12to4
    port map (
            O => \N__21608\,
            I => \N__21602\
        );

    \I__4930\ : Sp12to4
    port map (
            O => \N__21605\,
            I => \N__21599\
        );

    \I__4929\ : Span12Mux_s11_h
    port map (
            O => \N__21602\,
            I => \N__21596\
        );

    \I__4928\ : Span12Mux_v
    port map (
            O => \N__21599\,
            I => \N__21593\
        );

    \I__4927\ : Span12Mux_v
    port map (
            O => \N__21596\,
            I => \N__21588\
        );

    \I__4926\ : Span12Mux_h
    port map (
            O => \N__21593\,
            I => \N__21588\
        );

    \I__4925\ : Odrv12
    port map (
            O => \N__21588\,
            I => \DEBUG_c_5_c\
        );

    \I__4924\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21582\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__21582\,
            I => \tvp_video_buffer.BUFFER_0_6\
        );

    \I__4922\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21576\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__21576\,
            I => \N__21573\
        );

    \I__4920\ : Span4Mux_h
    port map (
            O => \N__21573\,
            I => \N__21570\
        );

    \I__4919\ : Span4Mux_h
    port map (
            O => \N__21570\,
            I => \N__21567\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__21567\,
            I => \line_buffer.n468\
        );

    \I__4917\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21561\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21558\
        );

    \I__4915\ : Span12Mux_h
    port map (
            O => \N__21558\,
            I => \N__21555\
        );

    \I__4914\ : Span12Mux_v
    port map (
            O => \N__21555\,
            I => \N__21552\
        );

    \I__4913\ : Odrv12
    port map (
            O => \N__21552\,
            I => \line_buffer.n460\
        );

    \I__4912\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21546\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__21546\,
            I => \N__21543\
        );

    \I__4910\ : Odrv4
    port map (
            O => \N__21543\,
            I => \line_buffer.n3548\
        );

    \I__4909\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21537\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__21537\,
            I => \N__21534\
        );

    \I__4907\ : Span12Mux_v
    port map (
            O => \N__21534\,
            I => \N__21531\
        );

    \I__4906\ : Odrv12
    port map (
            O => \N__21531\,
            I => \line_buffer.n567\
        );

    \I__4905\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21525\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__21525\,
            I => \N__21522\
        );

    \I__4903\ : Span4Mux_h
    port map (
            O => \N__21522\,
            I => \N__21519\
        );

    \I__4902\ : Sp12to4
    port map (
            O => \N__21519\,
            I => \N__21516\
        );

    \I__4901\ : Span12Mux_s7_h
    port map (
            O => \N__21516\,
            I => \N__21513\
        );

    \I__4900\ : Span12Mux_v
    port map (
            O => \N__21513\,
            I => \N__21510\
        );

    \I__4899\ : Odrv12
    port map (
            O => \N__21510\,
            I => \line_buffer.n559\
        );

    \I__4898\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21494\
        );

    \I__4897\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21491\
        );

    \I__4896\ : CascadeMux
    port map (
            O => \N__21505\,
            I => \N__21488\
        );

    \I__4895\ : CascadeMux
    port map (
            O => \N__21504\,
            I => \N__21485\
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__21503\,
            I => \N__21480\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__21502\,
            I => \N__21475\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__21501\,
            I => \N__21471\
        );

    \I__4891\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21468\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__21499\,
            I => \N__21465\
        );

    \I__4889\ : InMux
    port map (
            O => \N__21498\,
            I => \N__21460\
        );

    \I__4888\ : CascadeMux
    port map (
            O => \N__21497\,
            I => \N__21455\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21452\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21449\
        );

    \I__4885\ : InMux
    port map (
            O => \N__21488\,
            I => \N__21446\
        );

    \I__4884\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21443\
        );

    \I__4883\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21440\
        );

    \I__4882\ : InMux
    port map (
            O => \N__21483\,
            I => \N__21436\
        );

    \I__4881\ : InMux
    port map (
            O => \N__21480\,
            I => \N__21433\
        );

    \I__4880\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21426\
        );

    \I__4879\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21426\
        );

    \I__4878\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21426\
        );

    \I__4877\ : InMux
    port map (
            O => \N__21474\,
            I => \N__21421\
        );

    \I__4876\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21421\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__21468\,
            I => \N__21418\
        );

    \I__4874\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21415\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__21464\,
            I => \N__21411\
        );

    \I__4872\ : CascadeMux
    port map (
            O => \N__21463\,
            I => \N__21408\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__21460\,
            I => \N__21405\
        );

    \I__4870\ : InMux
    port map (
            O => \N__21459\,
            I => \N__21402\
        );

    \I__4869\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21397\
        );

    \I__4868\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21397\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__21452\,
            I => \N__21394\
        );

    \I__4866\ : Span4Mux_h
    port map (
            O => \N__21449\,
            I => \N__21389\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__21446\,
            I => \N__21389\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__21443\,
            I => \N__21386\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__21440\,
            I => \N__21383\
        );

    \I__4862\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21380\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__21436\,
            I => \N__21367\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__21433\,
            I => \N__21367\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__21426\,
            I => \N__21367\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21367\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__21418\,
            I => \N__21367\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__21415\,
            I => \N__21367\
        );

    \I__4855\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21362\
        );

    \I__4854\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21362\
        );

    \I__4853\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21359\
        );

    \I__4852\ : Span4Mux_v
    port map (
            O => \N__21405\,
            I => \N__21356\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__21402\,
            I => \N__21351\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__21397\,
            I => \N__21351\
        );

    \I__4849\ : Span4Mux_h
    port map (
            O => \N__21394\,
            I => \N__21344\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__21389\,
            I => \N__21344\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__21386\,
            I => \N__21344\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__21383\,
            I => \N__21337\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21337\
        );

    \I__4844\ : Span4Mux_v
    port map (
            O => \N__21367\,
            I => \N__21337\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__21362\,
            I => \TX_ADDR_12\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__21359\,
            I => \TX_ADDR_12\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__21356\,
            I => \TX_ADDR_12\
        );

    \I__4840\ : Odrv12
    port map (
            O => \N__21351\,
            I => \TX_ADDR_12\
        );

    \I__4839\ : Odrv4
    port map (
            O => \N__21344\,
            I => \TX_ADDR_12\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__21337\,
            I => \TX_ADDR_12\
        );

    \I__4837\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21321\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__21321\,
            I => \N__21318\
        );

    \I__4835\ : Span12Mux_h
    port map (
            O => \N__21318\,
            I => \N__21315\
        );

    \I__4834\ : Odrv12
    port map (
            O => \N__21315\,
            I => \line_buffer.n3540\
        );

    \I__4833\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21309\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__21309\,
            I => \line_buffer.n3573\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__21306\,
            I => \N__21301\
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__21305\,
            I => \N__21296\
        );

    \I__4829\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21290\
        );

    \I__4828\ : InMux
    port map (
            O => \N__21301\,
            I => \N__21287\
        );

    \I__4827\ : CascadeMux
    port map (
            O => \N__21300\,
            I => \N__21284\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__21299\,
            I => \N__21280\
        );

    \I__4825\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21277\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__21295\,
            I => \N__21274\
        );

    \I__4823\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21271\
        );

    \I__4822\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21264\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__21290\,
            I => \N__21261\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__21287\,
            I => \N__21258\
        );

    \I__4819\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21255\
        );

    \I__4818\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21252\
        );

    \I__4817\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21249\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__21277\,
            I => \N__21246\
        );

    \I__4815\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21243\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__21271\,
            I => \N__21240\
        );

    \I__4813\ : InMux
    port map (
            O => \N__21270\,
            I => \N__21237\
        );

    \I__4812\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21232\
        );

    \I__4811\ : InMux
    port map (
            O => \N__21268\,
            I => \N__21232\
        );

    \I__4810\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21229\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__21264\,
            I => \N__21225\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__21261\,
            I => \N__21220\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__21258\,
            I => \N__21220\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__21255\,
            I => \N__21217\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21212\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__21249\,
            I => \N__21212\
        );

    \I__4803\ : Span4Mux_v
    port map (
            O => \N__21246\,
            I => \N__21207\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__21243\,
            I => \N__21207\
        );

    \I__4801\ : Span4Mux_v
    port map (
            O => \N__21240\,
            I => \N__21202\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__21237\,
            I => \N__21202\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21197\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21197\
        );

    \I__4797\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21194\
        );

    \I__4796\ : Span4Mux_v
    port map (
            O => \N__21225\,
            I => \N__21189\
        );

    \I__4795\ : Span4Mux_h
    port map (
            O => \N__21220\,
            I => \N__21189\
        );

    \I__4794\ : Span4Mux_v
    port map (
            O => \N__21217\,
            I => \N__21186\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__21212\,
            I => \N__21181\
        );

    \I__4792\ : Span4Mux_v
    port map (
            O => \N__21207\,
            I => \N__21181\
        );

    \I__4791\ : Span4Mux_v
    port map (
            O => \N__21202\,
            I => \N__21174\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__21197\,
            I => \N__21174\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__21194\,
            I => \N__21174\
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__21189\,
            I => \TX_ADDR_13\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__21186\,
            I => \TX_ADDR_13\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__21181\,
            I => \TX_ADDR_13\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__21174\,
            I => \TX_ADDR_13\
        );

    \I__4784\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21162\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__21162\,
            I => \line_buffer.n3605\
        );

    \I__4782\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__21156\,
            I => \transmit_module.Y_DELTA_PATTERN_96\
        );

    \I__4780\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21150\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__21150\,
            I => \transmit_module.Y_DELTA_PATTERN_95\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__21144\,
            I => \transmit_module.Y_DELTA_PATTERN_94\
        );

    \I__4776\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__21138\,
            I => \transmit_module.Y_DELTA_PATTERN_93\
        );

    \I__4774\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__21132\,
            I => \N__21129\
        );

    \I__4772\ : Odrv12
    port map (
            O => \N__21129\,
            I => \transmit_module.Y_DELTA_PATTERN_83\
        );

    \I__4771\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21123\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__21123\,
            I => \N__21120\
        );

    \I__4769\ : Span4Mux_v
    port map (
            O => \N__21120\,
            I => \N__21117\
        );

    \I__4768\ : Sp12to4
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__4767\ : Odrv12
    port map (
            O => \N__21114\,
            I => \line_buffer.n593\
        );

    \I__4766\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21108\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__21108\,
            I => \N__21105\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__21105\,
            I => \N__21102\
        );

    \I__4763\ : Sp12to4
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__4762\ : Span12Mux_h
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__4761\ : Span12Mux_v
    port map (
            O => \N__21096\,
            I => \N__21093\
        );

    \I__4760\ : Odrv12
    port map (
            O => \N__21093\,
            I => \line_buffer.n585\
        );

    \I__4759\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21087\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__21087\,
            I => \line_buffer.n3641\
        );

    \I__4757\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21081\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__21081\,
            I => \N__21078\
        );

    \I__4755\ : Span12Mux_v
    port map (
            O => \N__21078\,
            I => \N__21075\
        );

    \I__4754\ : Odrv12
    port map (
            O => \N__21075\,
            I => \line_buffer.n533\
        );

    \I__4753\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21069\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__21069\,
            I => \N__21066\
        );

    \I__4751\ : Span4Mux_h
    port map (
            O => \N__21066\,
            I => \N__21063\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__21063\,
            I => \N__21060\
        );

    \I__4749\ : Odrv4
    port map (
            O => \N__21060\,
            I => \line_buffer.n525\
        );

    \I__4748\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__21054\,
            I => \N__21046\
        );

    \I__4746\ : InMux
    port map (
            O => \N__21053\,
            I => \N__21043\
        );

    \I__4745\ : InMux
    port map (
            O => \N__21052\,
            I => \N__21040\
        );

    \I__4744\ : InMux
    port map (
            O => \N__21051\,
            I => \N__21037\
        );

    \I__4743\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21034\
        );

    \I__4742\ : InMux
    port map (
            O => \N__21049\,
            I => \N__21030\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__21046\,
            I => \N__21026\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__21043\,
            I => \N__21017\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__21040\,
            I => \N__21017\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__21037\,
            I => \N__21017\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__21034\,
            I => \N__21017\
        );

    \I__4736\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21014\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__21030\,
            I => \N__21011\
        );

    \I__4734\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21008\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__21026\,
            I => \N__21004\
        );

    \I__4732\ : Span12Mux_v
    port map (
            O => \N__21017\,
            I => \N__20999\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__21014\,
            I => \N__20999\
        );

    \I__4730\ : Span4Mux_s1_v
    port map (
            O => \N__21011\,
            I => \N__20994\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__21008\,
            I => \N__20994\
        );

    \I__4728\ : InMux
    port map (
            O => \N__21007\,
            I => \N__20991\
        );

    \I__4727\ : Sp12to4
    port map (
            O => \N__21004\,
            I => \N__20988\
        );

    \I__4726\ : Span12Mux_v
    port map (
            O => \N__20999\,
            I => \N__20985\
        );

    \I__4725\ : Span4Mux_v
    port map (
            O => \N__20994\,
            I => \N__20982\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__20991\,
            I => \N__20979\
        );

    \I__4723\ : Span12Mux_v
    port map (
            O => \N__20988\,
            I => \N__20974\
        );

    \I__4722\ : Span12Mux_h
    port map (
            O => \N__20985\,
            I => \N__20974\
        );

    \I__4721\ : Span4Mux_h
    port map (
            O => \N__20982\,
            I => \N__20971\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__20979\,
            I => \N__20968\
        );

    \I__4719\ : Odrv12
    port map (
            O => \N__20974\,
            I => \RX_DATA_7\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__20971\,
            I => \RX_DATA_7\
        );

    \I__4717\ : Odrv4
    port map (
            O => \N__20968\,
            I => \RX_DATA_7\
        );

    \I__4716\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20958\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__20958\,
            I => \N__20955\
        );

    \I__4714\ : Span12Mux_v
    port map (
            O => \N__20955\,
            I => \N__20952\
        );

    \I__4713\ : Odrv12
    port map (
            O => \N__20952\,
            I => \line_buffer.n565\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20946\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20943\
        );

    \I__4710\ : Span4Mux_h
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__4709\ : Span4Mux_h
    port map (
            O => \N__20940\,
            I => \N__20937\
        );

    \I__4708\ : Odrv4
    port map (
            O => \N__20937\,
            I => \line_buffer.n557\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__20934\,
            I => \line_buffer.n3656_cascade_\
        );

    \I__4706\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20928\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__20928\,
            I => \line_buffer.n3596\
        );

    \I__4704\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20922\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__20922\,
            I => \line_buffer.n3638\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20919\,
            I => \N__20916\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20913\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__20913\,
            I => \N__20910\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__20910\,
            I => \TX_DATA_0\
        );

    \I__4698\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20901\
        );

    \I__4696\ : Span4Mux_v
    port map (
            O => \N__20901\,
            I => \N__20898\
        );

    \I__4695\ : Sp12to4
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__4694\ : Span12Mux_h
    port map (
            O => \N__20895\,
            I => \N__20892\
        );

    \I__4693\ : Span12Mux_v
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__4692\ : Odrv12
    port map (
            O => \N__20889\,
            I => \line_buffer.n530\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__20886\,
            I => \N__20883\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20880\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20877\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__20877\,
            I => \N__20874\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__20874\,
            I => \N__20871\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__20871\,
            I => \N__20868\
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__20868\,
            I => \line_buffer.n522\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20862\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__20862\,
            I => \line_buffer.n3632\
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__20859\,
            I => \line_buffer.n3650_cascade_\
        );

    \I__4681\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20853\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__4679\ : Span12Mux_h
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__4678\ : Odrv12
    port map (
            O => \N__20847\,
            I => \line_buffer.n594\
        );

    \I__4677\ : InMux
    port map (
            O => \N__20844\,
            I => \N__20841\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__20841\,
            I => \N__20838\
        );

    \I__4675\ : Span12Mux_h
    port map (
            O => \N__20838\,
            I => \N__20835\
        );

    \I__4674\ : Span12Mux_v
    port map (
            O => \N__20835\,
            I => \N__20832\
        );

    \I__4673\ : Odrv12
    port map (
            O => \N__20832\,
            I => \line_buffer.n586\
        );

    \I__4672\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20826\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__20826\,
            I => \line_buffer.n3647\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20820\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__20820\,
            I => \N__20817\
        );

    \I__4668\ : Span4Mux_h
    port map (
            O => \N__20817\,
            I => \N__20814\
        );

    \I__4667\ : Span4Mux_h
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__20811\,
            I => \N__20808\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__20808\,
            I => \line_buffer.n521\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20799\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__20796\,
            I => \N__20793\
        );

    \I__4660\ : Sp12to4
    port map (
            O => \N__20793\,
            I => \N__20790\
        );

    \I__4659\ : Span12Mux_h
    port map (
            O => \N__20790\,
            I => \N__20787\
        );

    \I__4658\ : Span12Mux_v
    port map (
            O => \N__20787\,
            I => \N__20784\
        );

    \I__4657\ : Odrv12
    port map (
            O => \N__20784\,
            I => \line_buffer.n529\
        );

    \I__4656\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__20778\,
            I => \line_buffer.n3644\
        );

    \I__4654\ : InMux
    port map (
            O => \N__20775\,
            I => \N__20772\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__20772\,
            I => \N__20769\
        );

    \I__4652\ : Odrv12
    port map (
            O => \N__20769\,
            I => \TX_DATA_5\
        );

    \I__4651\ : IoInMux
    port map (
            O => \N__20766\,
            I => \N__20763\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__20763\,
            I => \N__20759\
        );

    \I__4649\ : IoInMux
    port map (
            O => \N__20762\,
            I => \N__20756\
        );

    \I__4648\ : Span4Mux_s0_h
    port map (
            O => \N__20759\,
            I => \N__20753\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__20756\,
            I => \N__20750\
        );

    \I__4646\ : Span4Mux_h
    port map (
            O => \N__20753\,
            I => \N__20747\
        );

    \I__4645\ : Span4Mux_s3_v
    port map (
            O => \N__20750\,
            I => \N__20744\
        );

    \I__4644\ : Span4Mux_h
    port map (
            O => \N__20747\,
            I => \N__20740\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__20744\,
            I => \N__20737\
        );

    \I__4642\ : IoInMux
    port map (
            O => \N__20743\,
            I => \N__20734\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__20740\,
            I => \N__20731\
        );

    \I__4640\ : Span4Mux_h
    port map (
            O => \N__20737\,
            I => \N__20728\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__20734\,
            I => \N__20725\
        );

    \I__4638\ : Span4Mux_h
    port map (
            O => \N__20731\,
            I => \N__20720\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__20728\,
            I => \N__20720\
        );

    \I__4636\ : Span12Mux_s11_v
    port map (
            O => \N__20725\,
            I => \N__20717\
        );

    \I__4635\ : Span4Mux_v
    port map (
            O => \N__20720\,
            I => \N__20714\
        );

    \I__4634\ : Odrv12
    port map (
            O => \N__20717\,
            I => n1813
        );

    \I__4633\ : Odrv4
    port map (
            O => \N__20714\,
            I => n1813
        );

    \I__4632\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20706\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__20706\,
            I => \N__20703\
        );

    \I__4630\ : Odrv12
    port map (
            O => \N__20703\,
            I => \TX_DATA_1\
        );

    \I__4629\ : IoInMux
    port map (
            O => \N__20700\,
            I => \N__20697\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__20697\,
            I => \N__20693\
        );

    \I__4627\ : IoInMux
    port map (
            O => \N__20696\,
            I => \N__20690\
        );

    \I__4626\ : Span4Mux_s1_v
    port map (
            O => \N__20693\,
            I => \N__20687\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__20690\,
            I => \N__20684\
        );

    \I__4624\ : Span4Mux_v
    port map (
            O => \N__20687\,
            I => \N__20679\
        );

    \I__4623\ : Span4Mux_s2_h
    port map (
            O => \N__20684\,
            I => \N__20679\
        );

    \I__4622\ : Span4Mux_h
    port map (
            O => \N__20679\,
            I => \N__20675\
        );

    \I__4621\ : IoInMux
    port map (
            O => \N__20678\,
            I => \N__20672\
        );

    \I__4620\ : Sp12to4
    port map (
            O => \N__20675\,
            I => \N__20669\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__20672\,
            I => \N__20666\
        );

    \I__4618\ : Span12Mux_s10_v
    port map (
            O => \N__20669\,
            I => \N__20661\
        );

    \I__4617\ : Span12Mux_s10_v
    port map (
            O => \N__20666\,
            I => \N__20661\
        );

    \I__4616\ : Odrv12
    port map (
            O => \N__20661\,
            I => n1817
        );

    \I__4615\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20655\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__20655\,
            I => \transmit_module.Y_DELTA_PATTERN_97\
        );

    \I__4613\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20649\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__20649\,
            I => \transmit_module.Y_DELTA_PATTERN_92\
        );

    \I__4611\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__20643\,
            I => \transmit_module.Y_DELTA_PATTERN_91\
        );

    \I__4609\ : InMux
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__20637\,
            I => \transmit_module.Y_DELTA_PATTERN_90\
        );

    \I__4607\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20630\
        );

    \I__4606\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20622\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__20630\,
            I => \N__20619\
        );

    \I__4604\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20614\
        );

    \I__4603\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20614\
        );

    \I__4602\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20609\
        );

    \I__4601\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20609\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20606\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20601\
        );

    \I__4598\ : Span4Mux_h
    port map (
            O => \N__20619\,
            I => \N__20596\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__20614\,
            I => \N__20596\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20593\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__20606\,
            I => \N__20587\
        );

    \I__4594\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20584\
        );

    \I__4593\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20581\
        );

    \I__4592\ : Span4Mux_h
    port map (
            O => \N__20601\,
            I => \N__20576\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__20596\,
            I => \N__20573\
        );

    \I__4590\ : Span4Mux_h
    port map (
            O => \N__20593\,
            I => \N__20570\
        );

    \I__4589\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20567\
        );

    \I__4588\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20564\
        );

    \I__4587\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20561\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__20587\,
            I => \N__20554\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__20584\,
            I => \N__20554\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__20581\,
            I => \N__20554\
        );

    \I__4583\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20549\
        );

    \I__4582\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20549\
        );

    \I__4581\ : Odrv4
    port map (
            O => \N__20576\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__20573\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__20570\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__20567\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__20564\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__20561\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__20554\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__20549\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4573\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20529\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__20529\,
            I => \transmit_module.Y_DELTA_PATTERN_99\
        );

    \I__4571\ : CEMux
    port map (
            O => \N__20526\,
            I => \N__20522\
        );

    \I__4570\ : CEMux
    port map (
            O => \N__20525\,
            I => \N__20519\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__20522\,
            I => \N__20511\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20507\
        );

    \I__4567\ : CEMux
    port map (
            O => \N__20518\,
            I => \N__20504\
        );

    \I__4566\ : CEMux
    port map (
            O => \N__20517\,
            I => \N__20500\
        );

    \I__4565\ : CEMux
    port map (
            O => \N__20516\,
            I => \N__20496\
        );

    \I__4564\ : SRMux
    port map (
            O => \N__20515\,
            I => \N__20493\
        );

    \I__4563\ : CEMux
    port map (
            O => \N__20514\,
            I => \N__20489\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__20511\,
            I => \N__20483\
        );

    \I__4561\ : CEMux
    port map (
            O => \N__20510\,
            I => \N__20480\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__20507\,
            I => \N__20475\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__20504\,
            I => \N__20475\
        );

    \I__4558\ : CEMux
    port map (
            O => \N__20503\,
            I => \N__20472\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__20500\,
            I => \N__20469\
        );

    \I__4556\ : CEMux
    port map (
            O => \N__20499\,
            I => \N__20466\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__20496\,
            I => \N__20463\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__20493\,
            I => \N__20460\
        );

    \I__4553\ : SRMux
    port map (
            O => \N__20492\,
            I => \N__20457\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__20489\,
            I => \N__20454\
        );

    \I__4551\ : CEMux
    port map (
            O => \N__20488\,
            I => \N__20451\
        );

    \I__4550\ : CEMux
    port map (
            O => \N__20487\,
            I => \N__20448\
        );

    \I__4549\ : SRMux
    port map (
            O => \N__20486\,
            I => \N__20445\
        );

    \I__4548\ : Span4Mux_v
    port map (
            O => \N__20483\,
            I => \N__20440\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__20480\,
            I => \N__20440\
        );

    \I__4546\ : Span4Mux_h
    port map (
            O => \N__20475\,
            I => \N__20437\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__20472\,
            I => \N__20434\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__20469\,
            I => \N__20429\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__20466\,
            I => \N__20429\
        );

    \I__4542\ : Span4Mux_v
    port map (
            O => \N__20463\,
            I => \N__20426\
        );

    \I__4541\ : Span4Mux_v
    port map (
            O => \N__20460\,
            I => \N__20423\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__20457\,
            I => \N__20420\
        );

    \I__4539\ : Span4Mux_h
    port map (
            O => \N__20454\,
            I => \N__20414\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__20451\,
            I => \N__20414\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__20448\,
            I => \N__20411\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__20445\,
            I => \N__20408\
        );

    \I__4535\ : Span4Mux_v
    port map (
            O => \N__20440\,
            I => \N__20405\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__20437\,
            I => \N__20400\
        );

    \I__4533\ : Span4Mux_v
    port map (
            O => \N__20434\,
            I => \N__20400\
        );

    \I__4532\ : Span4Mux_h
    port map (
            O => \N__20429\,
            I => \N__20391\
        );

    \I__4531\ : Span4Mux_h
    port map (
            O => \N__20426\,
            I => \N__20391\
        );

    \I__4530\ : Span4Mux_h
    port map (
            O => \N__20423\,
            I => \N__20391\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__20420\,
            I => \N__20391\
        );

    \I__4528\ : SRMux
    port map (
            O => \N__20419\,
            I => \N__20388\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__20414\,
            I => \N__20381\
        );

    \I__4526\ : Span4Mux_v
    port map (
            O => \N__20411\,
            I => \N__20381\
        );

    \I__4525\ : Span4Mux_h
    port map (
            O => \N__20408\,
            I => \N__20381\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__20405\,
            I => \transmit_module.n3679\
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__20400\,
            I => \transmit_module.n3679\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__20391\,
            I => \transmit_module.n3679\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__20388\,
            I => \transmit_module.n3679\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__20381\,
            I => \transmit_module.n3679\
        );

    \I__4519\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20367\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__20367\,
            I => \N__20364\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__20364\,
            I => \N__20361\
        );

    \I__4516\ : Span4Mux_v
    port map (
            O => \N__20361\,
            I => \N__20358\
        );

    \I__4515\ : Sp12to4
    port map (
            O => \N__20358\,
            I => \N__20355\
        );

    \I__4514\ : Odrv12
    port map (
            O => \N__20355\,
            I => \line_buffer.n566\
        );

    \I__4513\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20349\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__20349\,
            I => \N__20346\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__20346\,
            I => \N__20343\
        );

    \I__4510\ : Span4Mux_h
    port map (
            O => \N__20343\,
            I => \N__20340\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__20340\,
            I => \line_buffer.n558\
        );

    \I__4508\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20334\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__20334\,
            I => \N__20331\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__20331\,
            I => \N__20328\
        );

    \I__4505\ : Span4Mux_v
    port map (
            O => \N__20328\,
            I => \N__20325\
        );

    \I__4504\ : Span4Mux_h
    port map (
            O => \N__20325\,
            I => \N__20322\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__20322\,
            I => \line_buffer.n465\
        );

    \I__4502\ : CascadeMux
    port map (
            O => \N__20319\,
            I => \N__20316\
        );

    \I__4501\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20313\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__20313\,
            I => \N__20310\
        );

    \I__4499\ : Span12Mux_h
    port map (
            O => \N__20310\,
            I => \N__20307\
        );

    \I__4498\ : Span12Mux_v
    port map (
            O => \N__20307\,
            I => \N__20304\
        );

    \I__4497\ : Odrv12
    port map (
            O => \N__20304\,
            I => \line_buffer.n457\
        );

    \I__4496\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__20298\,
            I => \line_buffer.n3629\
        );

    \I__4494\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20292\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__20292\,
            I => \N__20289\
        );

    \I__4492\ : Span4Mux_v
    port map (
            O => \N__20289\,
            I => \N__20286\
        );

    \I__4491\ : Span4Mux_v
    port map (
            O => \N__20286\,
            I => \N__20283\
        );

    \I__4490\ : Sp12to4
    port map (
            O => \N__20283\,
            I => \N__20280\
        );

    \I__4489\ : Odrv12
    port map (
            O => \N__20280\,
            I => \line_buffer.n561\
        );

    \I__4488\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20274\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__20274\,
            I => \N__20271\
        );

    \I__4486\ : Span4Mux_h
    port map (
            O => \N__20271\,
            I => \N__20268\
        );

    \I__4485\ : Span4Mux_h
    port map (
            O => \N__20268\,
            I => \N__20265\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__20265\,
            I => \line_buffer.n553\
        );

    \I__4483\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20259\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__20259\,
            I => \N__20256\
        );

    \I__4481\ : Span4Mux_h
    port map (
            O => \N__20256\,
            I => \N__20253\
        );

    \I__4480\ : Span4Mux_h
    port map (
            O => \N__20253\,
            I => \N__20250\
        );

    \I__4479\ : Span4Mux_v
    port map (
            O => \N__20250\,
            I => \N__20247\
        );

    \I__4478\ : Span4Mux_v
    port map (
            O => \N__20247\,
            I => \N__20244\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__20244\,
            I => \line_buffer.n456\
        );

    \I__4476\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__20238\,
            I => \N__20235\
        );

    \I__4474\ : Span4Mux_v
    port map (
            O => \N__20235\,
            I => \N__20232\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__20232\,
            I => \N__20229\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__20229\,
            I => \N__20226\
        );

    \I__4471\ : Odrv4
    port map (
            O => \N__20226\,
            I => \line_buffer.n464\
        );

    \I__4470\ : CascadeMux
    port map (
            O => \N__20223\,
            I => \line_buffer.n3635_cascade_\
        );

    \I__4469\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20217\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__20217\,
            I => \N__20214\
        );

    \I__4467\ : Span4Mux_h
    port map (
            O => \N__20214\,
            I => \N__20211\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__20211\,
            I => \N__20208\
        );

    \I__4465\ : Odrv4
    port map (
            O => \N__20208\,
            I => \line_buffer.n469\
        );

    \I__4464\ : InMux
    port map (
            O => \N__20205\,
            I => \N__20202\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__20202\,
            I => \N__20199\
        );

    \I__4462\ : Span12Mux_h
    port map (
            O => \N__20199\,
            I => \N__20196\
        );

    \I__4461\ : Span12Mux_v
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__4460\ : Odrv12
    port map (
            O => \N__20193\,
            I => \line_buffer.n461\
        );

    \I__4459\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20187\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__20187\,
            I => \N__20184\
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__20184\,
            I => \line_buffer.n3653\
        );

    \I__4456\ : IoInMux
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20175\
        );

    \I__4454\ : IoSpan4Mux
    port map (
            O => \N__20175\,
            I => \N__20172\
        );

    \I__4453\ : Span4Mux_s2_h
    port map (
            O => \N__20172\,
            I => \N__20169\
        );

    \I__4452\ : Span4Mux_h
    port map (
            O => \N__20169\,
            I => \N__20165\
        );

    \I__4451\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20162\
        );

    \I__4450\ : Sp12to4
    port map (
            O => \N__20165\,
            I => \N__20157\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__20162\,
            I => \N__20157\
        );

    \I__4448\ : Span12Mux_h
    port map (
            O => \N__20157\,
            I => \N__20154\
        );

    \I__4447\ : Odrv12
    port map (
            O => \N__20154\,
            I => \DEBUG_c_2_c\
        );

    \I__4446\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20148\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__20148\,
            I => \tvp_hs_buffer.BUFFER_0_0\
        );

    \I__4444\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20142\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__20142\,
            I => \tvp_hs_buffer.BUFFER_1_0\
        );

    \I__4442\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20126\
        );

    \I__4441\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20119\
        );

    \I__4440\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20119\
        );

    \I__4439\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20119\
        );

    \I__4438\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20112\
        );

    \I__4437\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20112\
        );

    \I__4436\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20112\
        );

    \I__4435\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20105\
        );

    \I__4434\ : InMux
    port map (
            O => \N__20131\,
            I => \N__20105\
        );

    \I__4433\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20105\
        );

    \I__4432\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20101\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__20126\,
            I => \N__20097\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__20119\,
            I => \N__20089\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__20112\,
            I => \N__20089\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__20105\,
            I => \N__20089\
        );

    \I__4427\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20086\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__20101\,
            I => \N__20083\
        );

    \I__4425\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20080\
        );

    \I__4424\ : Span12Mux_s2_v
    port map (
            O => \N__20097\,
            I => \N__20076\
        );

    \I__4423\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20073\
        );

    \I__4422\ : Span4Mux_v
    port map (
            O => \N__20089\,
            I => \N__20068\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__20086\,
            I => \N__20068\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__20083\,
            I => \N__20063\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__20080\,
            I => \N__20060\
        );

    \I__4418\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20057\
        );

    \I__4417\ : Span12Mux_v
    port map (
            O => \N__20076\,
            I => \N__20051\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__20073\,
            I => \N__20051\
        );

    \I__4415\ : Span4Mux_v
    port map (
            O => \N__20068\,
            I => \N__20048\
        );

    \I__4414\ : InMux
    port map (
            O => \N__20067\,
            I => \N__20043\
        );

    \I__4413\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20043\
        );

    \I__4412\ : Span4Mux_v
    port map (
            O => \N__20063\,
            I => \N__20036\
        );

    \I__4411\ : Span4Mux_v
    port map (
            O => \N__20060\,
            I => \N__20036\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__20057\,
            I => \N__20036\
        );

    \I__4409\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20033\
        );

    \I__4408\ : Odrv12
    port map (
            O => \N__20051\,
            I => \TVP_VSYNC_buff\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__20048\,
            I => \TVP_VSYNC_buff\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__20043\,
            I => \TVP_VSYNC_buff\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__20036\,
            I => \TVP_VSYNC_buff\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__20033\,
            I => \TVP_VSYNC_buff\
        );

    \I__4403\ : CEMux
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__20019\,
            I => \N__20015\
        );

    \I__4401\ : CEMux
    port map (
            O => \N__20018\,
            I => \N__20012\
        );

    \I__4400\ : Span4Mux_h
    port map (
            O => \N__20015\,
            I => \N__20009\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__20012\,
            I => \N__20006\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__20009\,
            I => \receive_module.rx_counter.n2078\
        );

    \I__4397\ : Odrv12
    port map (
            O => \N__20006\,
            I => \receive_module.rx_counter.n2078\
        );

    \I__4396\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19996\
        );

    \I__4395\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19991\
        );

    \I__4394\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19991\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__19996\,
            I => \N__19988\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__19991\,
            I => \TVP_HSYNC_buff\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__19988\,
            I => \TVP_HSYNC_buff\
        );

    \I__4390\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19980\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__19980\,
            I => \receive_module.rx_counter.old_HS\
        );

    \I__4388\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__19974\,
            I => \transmit_module.Y_DELTA_PATTERN_98\
        );

    \I__4386\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19968\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19968\,
            I => \transmit_module.Y_DELTA_PATTERN_89\
        );

    \I__4384\ : IoInMux
    port map (
            O => \N__19965\,
            I => \N__19962\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__19962\,
            I => \N__19959\
        );

    \I__4382\ : IoSpan4Mux
    port map (
            O => \N__19959\,
            I => \N__19956\
        );

    \I__4381\ : Span4Mux_s3_h
    port map (
            O => \N__19956\,
            I => \N__19952\
        );

    \I__4380\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19949\
        );

    \I__4379\ : Sp12to4
    port map (
            O => \N__19952\,
            I => \N__19946\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__19949\,
            I => \N__19943\
        );

    \I__4377\ : Span12Mux_v
    port map (
            O => \N__19946\,
            I => \N__19940\
        );

    \I__4376\ : Span12Mux_h
    port map (
            O => \N__19943\,
            I => \N__19937\
        );

    \I__4375\ : Span12Mux_h
    port map (
            O => \N__19940\,
            I => \N__19934\
        );

    \I__4374\ : Span12Mux_v
    port map (
            O => \N__19937\,
            I => \N__19931\
        );

    \I__4373\ : Odrv12
    port map (
            O => \N__19934\,
            I => \DEBUG_c_7_c\
        );

    \I__4372\ : Odrv12
    port map (
            O => \N__19931\,
            I => \DEBUG_c_7_c\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__19923\,
            I => \N__19918\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19915\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19921\,
            I => \N__19911\
        );

    \I__4367\ : Span4Mux_s2_v
    port map (
            O => \N__19918\,
            I => \N__19904\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__19915\,
            I => \N__19904\
        );

    \I__4365\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19901\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19898\
        );

    \I__4363\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19895\
        );

    \I__4362\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19892\
        );

    \I__4361\ : Span4Mux_v
    port map (
            O => \N__19904\,
            I => \N__19888\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19885\
        );

    \I__4359\ : Span4Mux_v
    port map (
            O => \N__19898\,
            I => \N__19878\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__19895\,
            I => \N__19878\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19878\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19875\
        );

    \I__4355\ : Span4Mux_h
    port map (
            O => \N__19888\,
            I => \N__19870\
        );

    \I__4354\ : Span4Mux_v
    port map (
            O => \N__19885\,
            I => \N__19867\
        );

    \I__4353\ : Span4Mux_v
    port map (
            O => \N__19878\,
            I => \N__19862\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__19875\,
            I => \N__19862\
        );

    \I__4351\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19859\
        );

    \I__4350\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19856\
        );

    \I__4349\ : Sp12to4
    port map (
            O => \N__19870\,
            I => \N__19853\
        );

    \I__4348\ : Span4Mux_h
    port map (
            O => \N__19867\,
            I => \N__19850\
        );

    \I__4347\ : Span4Mux_v
    port map (
            O => \N__19862\,
            I => \N__19845\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__19859\,
            I => \N__19845\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__19856\,
            I => \N__19842\
        );

    \I__4344\ : Span12Mux_v
    port map (
            O => \N__19853\,
            I => \N__19837\
        );

    \I__4343\ : Sp12to4
    port map (
            O => \N__19850\,
            I => \N__19837\
        );

    \I__4342\ : Span4Mux_v
    port map (
            O => \N__19845\,
            I => \N__19834\
        );

    \I__4341\ : Span4Mux_h
    port map (
            O => \N__19842\,
            I => \N__19831\
        );

    \I__4340\ : Span12Mux_v
    port map (
            O => \N__19837\,
            I => \N__19826\
        );

    \I__4339\ : Sp12to4
    port map (
            O => \N__19834\,
            I => \N__19826\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__19831\,
            I => \N__19823\
        );

    \I__4337\ : Odrv12
    port map (
            O => \N__19826\,
            I => \RX_DATA_6\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__19823\,
            I => \RX_DATA_6\
        );

    \I__4335\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19815\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__19815\,
            I => \tvp_video_buffer.BUFFER_0_8\
        );

    \I__4333\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19809\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__19809\,
            I => \tvp_video_buffer.BUFFER_1_8\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19803\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__4329\ : Span4Mux_v
    port map (
            O => \N__19800\,
            I => \N__19797\
        );

    \I__4328\ : Sp12to4
    port map (
            O => \N__19797\,
            I => \N__19794\
        );

    \I__4327\ : Odrv12
    port map (
            O => \N__19794\,
            I => \line_buffer.n598\
        );

    \I__4326\ : InMux
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__19788\,
            I => \N__19785\
        );

    \I__4324\ : Span12Mux_v
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__4323\ : Odrv12
    port map (
            O => \N__19782\,
            I => \line_buffer.n590\
        );

    \I__4322\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19776\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19776\,
            I => \N__19773\
        );

    \I__4320\ : Sp12to4
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__4319\ : Span12Mux_v
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__4318\ : Odrv12
    port map (
            O => \N__19767\,
            I => \line_buffer.n526\
        );

    \I__4317\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19761\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__19761\,
            I => \N__19758\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__4314\ : Sp12to4
    port map (
            O => \N__19755\,
            I => \N__19752\
        );

    \I__4313\ : Span12Mux_h
    port map (
            O => \N__19752\,
            I => \N__19749\
        );

    \I__4312\ : Span12Mux_v
    port map (
            O => \N__19749\,
            I => \N__19746\
        );

    \I__4311\ : Odrv12
    port map (
            O => \N__19746\,
            I => \line_buffer.n534\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__19743\,
            I => \line_buffer.n3593_cascade_\
        );

    \I__4309\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19737\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__19737\,
            I => \N__19734\
        );

    \I__4307\ : Odrv12
    port map (
            O => \N__19734\,
            I => \line_buffer.n554\
        );

    \I__4306\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19728\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__4304\ : Span4Mux_v
    port map (
            O => \N__19725\,
            I => \N__19722\
        );

    \I__4303\ : Span4Mux_h
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__4302\ : Span4Mux_h
    port map (
            O => \N__19719\,
            I => \N__19716\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__19716\,
            I => \line_buffer.n562\
        );

    \I__4300\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19710\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19710\,
            I => \N__19707\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__19707\,
            I => \N__19704\
        );

    \I__4297\ : Odrv4
    port map (
            O => \N__19704\,
            I => \receive_module.n132\
        );

    \I__4296\ : IoInMux
    port map (
            O => \N__19701\,
            I => \N__19698\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19694\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__19697\,
            I => \N__19691\
        );

    \I__4293\ : Span4Mux_s3_h
    port map (
            O => \N__19694\,
            I => \N__19687\
        );

    \I__4292\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19681\
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__19690\,
            I => \N__19677\
        );

    \I__4290\ : Span4Mux_h
    port map (
            O => \N__19687\,
            I => \N__19673\
        );

    \I__4289\ : CascadeMux
    port map (
            O => \N__19686\,
            I => \N__19664\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__19685\,
            I => \N__19661\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__19684\,
            I => \N__19656\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__19681\,
            I => \N__19653\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19650\
        );

    \I__4284\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19646\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__19676\,
            I => \N__19642\
        );

    \I__4282\ : Span4Mux_h
    port map (
            O => \N__19673\,
            I => \N__19638\
        );

    \I__4281\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19631\
        );

    \I__4280\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19631\
        );

    \I__4279\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19631\
        );

    \I__4278\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19626\
        );

    \I__4277\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19626\
        );

    \I__4276\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19613\
        );

    \I__4275\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19613\
        );

    \I__4274\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19613\
        );

    \I__4273\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19613\
        );

    \I__4272\ : InMux
    port map (
            O => \N__19659\,
            I => \N__19613\
        );

    \I__4271\ : InMux
    port map (
            O => \N__19656\,
            I => \N__19613\
        );

    \I__4270\ : Sp12to4
    port map (
            O => \N__19653\,
            I => \N__19608\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__19650\,
            I => \N__19608\
        );

    \I__4268\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19605\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19602\
        );

    \I__4266\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19595\
        );

    \I__4265\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19595\
        );

    \I__4264\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19595\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__19638\,
            I => \N__19586\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__19631\,
            I => \N__19586\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__19626\,
            I => \N__19583\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__19613\,
            I => \N__19576\
        );

    \I__4259\ : Span12Mux_v
    port map (
            O => \N__19608\,
            I => \N__19576\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__19605\,
            I => \N__19576\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__19602\,
            I => \N__19571\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__19595\,
            I => \N__19571\
        );

    \I__4255\ : InMux
    port map (
            O => \N__19594\,
            I => \N__19568\
        );

    \I__4254\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19565\
        );

    \I__4253\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19560\
        );

    \I__4252\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19560\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__19586\,
            I => \N__19555\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__19583\,
            I => \N__19555\
        );

    \I__4249\ : Odrv12
    port map (
            O => \N__19576\,
            I => \DEBUG_c_4\
        );

    \I__4248\ : Odrv4
    port map (
            O => \N__19571\,
            I => \DEBUG_c_4\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__19568\,
            I => \DEBUG_c_4\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__19565\,
            I => \DEBUG_c_4\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__19560\,
            I => \DEBUG_c_4\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__19555\,
            I => \DEBUG_c_4\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__19542\,
            I => \N__19538\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__19541\,
            I => \N__19535\
        );

    \I__4241\ : CascadeBuf
    port map (
            O => \N__19538\,
            I => \N__19532\
        );

    \I__4240\ : CascadeBuf
    port map (
            O => \N__19535\,
            I => \N__19529\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__19532\,
            I => \N__19526\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__19529\,
            I => \N__19523\
        );

    \I__4237\ : CascadeBuf
    port map (
            O => \N__19526\,
            I => \N__19520\
        );

    \I__4236\ : CascadeBuf
    port map (
            O => \N__19523\,
            I => \N__19517\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__19520\,
            I => \N__19514\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__19517\,
            I => \N__19511\
        );

    \I__4233\ : CascadeBuf
    port map (
            O => \N__19514\,
            I => \N__19508\
        );

    \I__4232\ : CascadeBuf
    port map (
            O => \N__19511\,
            I => \N__19505\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__19508\,
            I => \N__19502\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__19505\,
            I => \N__19499\
        );

    \I__4229\ : CascadeBuf
    port map (
            O => \N__19502\,
            I => \N__19496\
        );

    \I__4228\ : CascadeBuf
    port map (
            O => \N__19499\,
            I => \N__19493\
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__19496\,
            I => \N__19490\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__19493\,
            I => \N__19487\
        );

    \I__4225\ : CascadeBuf
    port map (
            O => \N__19490\,
            I => \N__19484\
        );

    \I__4224\ : CascadeBuf
    port map (
            O => \N__19487\,
            I => \N__19481\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \N__19478\
        );

    \I__4222\ : CascadeMux
    port map (
            O => \N__19481\,
            I => \N__19475\
        );

    \I__4221\ : CascadeBuf
    port map (
            O => \N__19478\,
            I => \N__19472\
        );

    \I__4220\ : CascadeBuf
    port map (
            O => \N__19475\,
            I => \N__19469\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__19472\,
            I => \N__19466\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__19469\,
            I => \N__19463\
        );

    \I__4217\ : CascadeBuf
    port map (
            O => \N__19466\,
            I => \N__19460\
        );

    \I__4216\ : CascadeBuf
    port map (
            O => \N__19463\,
            I => \N__19457\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__19460\,
            I => \N__19454\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__19457\,
            I => \N__19451\
        );

    \I__4213\ : CascadeBuf
    port map (
            O => \N__19454\,
            I => \N__19448\
        );

    \I__4212\ : CascadeBuf
    port map (
            O => \N__19451\,
            I => \N__19445\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__19448\,
            I => \N__19442\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__19445\,
            I => \N__19439\
        );

    \I__4209\ : CascadeBuf
    port map (
            O => \N__19442\,
            I => \N__19436\
        );

    \I__4208\ : CascadeBuf
    port map (
            O => \N__19439\,
            I => \N__19433\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__19436\,
            I => \N__19430\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__19433\,
            I => \N__19427\
        );

    \I__4205\ : CascadeBuf
    port map (
            O => \N__19430\,
            I => \N__19424\
        );

    \I__4204\ : CascadeBuf
    port map (
            O => \N__19427\,
            I => \N__19421\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__19424\,
            I => \N__19418\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__19421\,
            I => \N__19415\
        );

    \I__4201\ : CascadeBuf
    port map (
            O => \N__19418\,
            I => \N__19412\
        );

    \I__4200\ : CascadeBuf
    port map (
            O => \N__19415\,
            I => \N__19409\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__19412\,
            I => \N__19406\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__19409\,
            I => \N__19403\
        );

    \I__4197\ : CascadeBuf
    port map (
            O => \N__19406\,
            I => \N__19400\
        );

    \I__4196\ : CascadeBuf
    port map (
            O => \N__19403\,
            I => \N__19397\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__19400\,
            I => \N__19394\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__19397\,
            I => \N__19391\
        );

    \I__4193\ : CascadeBuf
    port map (
            O => \N__19394\,
            I => \N__19388\
        );

    \I__4192\ : CascadeBuf
    port map (
            O => \N__19391\,
            I => \N__19385\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__19388\,
            I => \N__19382\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__19385\,
            I => \N__19379\
        );

    \I__4189\ : CascadeBuf
    port map (
            O => \N__19382\,
            I => \N__19376\
        );

    \I__4188\ : CascadeBuf
    port map (
            O => \N__19379\,
            I => \N__19373\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__19376\,
            I => \N__19370\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__19373\,
            I => \N__19367\
        );

    \I__4185\ : CascadeBuf
    port map (
            O => \N__19370\,
            I => \N__19364\
        );

    \I__4184\ : CascadeBuf
    port map (
            O => \N__19367\,
            I => \N__19361\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__19364\,
            I => \N__19358\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__19361\,
            I => \N__19355\
        );

    \I__4181\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19352\
        );

    \I__4180\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19349\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N__19345\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__19349\,
            I => \N__19342\
        );

    \I__4177\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19339\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__19345\,
            I => \N__19336\
        );

    \I__4175\ : Span4Mux_s2_v
    port map (
            O => \N__19342\,
            I => \N__19333\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__19339\,
            I => \N__19330\
        );

    \I__4173\ : Sp12to4
    port map (
            O => \N__19336\,
            I => \N__19326\
        );

    \I__4172\ : Sp12to4
    port map (
            O => \N__19333\,
            I => \N__19323\
        );

    \I__4171\ : Span4Mux_h
    port map (
            O => \N__19330\,
            I => \N__19320\
        );

    \I__4170\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19317\
        );

    \I__4169\ : Span12Mux_v
    port map (
            O => \N__19326\,
            I => \N__19314\
        );

    \I__4168\ : Span12Mux_h
    port map (
            O => \N__19323\,
            I => \N__19311\
        );

    \I__4167\ : Odrv4
    port map (
            O => \N__19320\,
            I => \RX_ADDR_5\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__19317\,
            I => \RX_ADDR_5\
        );

    \I__4165\ : Odrv12
    port map (
            O => \N__19314\,
            I => \RX_ADDR_5\
        );

    \I__4164\ : Odrv12
    port map (
            O => \N__19311\,
            I => \RX_ADDR_5\
        );

    \I__4163\ : SRMux
    port map (
            O => \N__19302\,
            I => \N__19295\
        );

    \I__4162\ : SRMux
    port map (
            O => \N__19301\,
            I => \N__19292\
        );

    \I__4161\ : SRMux
    port map (
            O => \N__19300\,
            I => \N__19288\
        );

    \I__4160\ : SRMux
    port map (
            O => \N__19299\,
            I => \N__19285\
        );

    \I__4159\ : SRMux
    port map (
            O => \N__19298\,
            I => \N__19282\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__19295\,
            I => \N__19279\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19276\
        );

    \I__4156\ : SRMux
    port map (
            O => \N__19291\,
            I => \N__19273\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__19288\,
            I => \N__19269\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__19285\,
            I => \N__19266\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__19282\,
            I => \N__19263\
        );

    \I__4152\ : Sp12to4
    port map (
            O => \N__19279\,
            I => \N__19260\
        );

    \I__4151\ : Span4Mux_h
    port map (
            O => \N__19276\,
            I => \N__19255\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__19273\,
            I => \N__19255\
        );

    \I__4149\ : SRMux
    port map (
            O => \N__19272\,
            I => \N__19252\
        );

    \I__4148\ : Span4Mux_v
    port map (
            O => \N__19269\,
            I => \N__19249\
        );

    \I__4147\ : Span4Mux_h
    port map (
            O => \N__19266\,
            I => \N__19246\
        );

    \I__4146\ : Span4Mux_h
    port map (
            O => \N__19263\,
            I => \N__19243\
        );

    \I__4145\ : Span12Mux_s9_v
    port map (
            O => \N__19260\,
            I => \N__19236\
        );

    \I__4144\ : Sp12to4
    port map (
            O => \N__19255\,
            I => \N__19236\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__19252\,
            I => \N__19236\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__19249\,
            I => \receive_module.n3674\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__19246\,
            I => \receive_module.n3674\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__19243\,
            I => \receive_module.n3674\
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__19236\,
            I => \receive_module.n3674\
        );

    \I__4138\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__19224\,
            I => \N__19221\
        );

    \I__4136\ : Span4Mux_v
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__4135\ : Sp12to4
    port map (
            O => \N__19218\,
            I => \N__19215\
        );

    \I__4134\ : Odrv12
    port map (
            O => \N__19215\,
            I => \line_buffer.n596\
        );

    \I__4133\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19209\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__19209\,
            I => \N__19206\
        );

    \I__4131\ : Span12Mux_v
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__4130\ : Odrv12
    port map (
            O => \N__19203\,
            I => \line_buffer.n588\
        );

    \I__4129\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__19197\,
            I => \line_buffer.n3623\
        );

    \I__4127\ : InMux
    port map (
            O => \N__19194\,
            I => \bfn_17_10_0_\
        );

    \I__4126\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19187\
        );

    \I__4125\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19184\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__19187\,
            I => \N__19181\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__19184\,
            I => \N__19174\
        );

    \I__4122\ : Span4Mux_v
    port map (
            O => \N__19181\,
            I => \N__19174\
        );

    \I__4121\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19169\
        );

    \I__4120\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19169\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__19174\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__19169\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__4117\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19161\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__19158\,
            I => \tvp_video_buffer.BUFFER_1_2\
        );

    \I__4114\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19152\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__4112\ : Span4Mux_s1_v
    port map (
            O => \N__19149\,
            I => \N__19145\
        );

    \I__4111\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19142\
        );

    \I__4110\ : Span4Mux_v
    port map (
            O => \N__19145\,
            I => \N__19135\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19135\
        );

    \I__4108\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19130\
        );

    \I__4107\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19126\
        );

    \I__4106\ : Span4Mux_v
    port map (
            O => \N__19135\,
            I => \N__19123\
        );

    \I__4105\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19120\
        );

    \I__4104\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19116\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__19130\,
            I => \N__19113\
        );

    \I__4102\ : InMux
    port map (
            O => \N__19129\,
            I => \N__19110\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__19126\,
            I => \N__19107\
        );

    \I__4100\ : Span4Mux_v
    port map (
            O => \N__19123\,
            I => \N__19102\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19102\
        );

    \I__4098\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19099\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__19116\,
            I => \N__19096\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__19113\,
            I => \N__19093\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__19110\,
            I => \N__19090\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__19107\,
            I => \N__19087\
        );

    \I__4093\ : Span4Mux_v
    port map (
            O => \N__19102\,
            I => \N__19082\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__19099\,
            I => \N__19082\
        );

    \I__4091\ : Sp12to4
    port map (
            O => \N__19096\,
            I => \N__19079\
        );

    \I__4090\ : Span4Mux_v
    port map (
            O => \N__19093\,
            I => \N__19074\
        );

    \I__4089\ : Span4Mux_v
    port map (
            O => \N__19090\,
            I => \N__19074\
        );

    \I__4088\ : Span4Mux_v
    port map (
            O => \N__19087\,
            I => \N__19069\
        );

    \I__4087\ : Span4Mux_v
    port map (
            O => \N__19082\,
            I => \N__19069\
        );

    \I__4086\ : Span12Mux_v
    port map (
            O => \N__19079\,
            I => \N__19064\
        );

    \I__4085\ : Sp12to4
    port map (
            O => \N__19074\,
            I => \N__19064\
        );

    \I__4084\ : Span4Mux_h
    port map (
            O => \N__19069\,
            I => \N__19061\
        );

    \I__4083\ : Odrv12
    port map (
            O => \N__19064\,
            I => \RX_DATA_0\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__19061\,
            I => \RX_DATA_0\
        );

    \I__4081\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19052\
        );

    \I__4080\ : InMux
    port map (
            O => \N__19055\,
            I => \N__19049\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__19052\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__19049\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__4077\ : InMux
    port map (
            O => \N__19044\,
            I => \N__19040\
        );

    \I__4076\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19037\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__19040\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__19037\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__4073\ : InMux
    port map (
            O => \N__19032\,
            I => \N__19028\
        );

    \I__4072\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19025\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__19028\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__19025\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__4069\ : InMux
    port map (
            O => \N__19020\,
            I => \N__19016\
        );

    \I__4068\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19013\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__19016\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__19013\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__19008\,
            I => \receive_module.rx_counter.n7_adj_619_cascade_\
        );

    \I__4064\ : InMux
    port map (
            O => \N__19005\,
            I => \N__19002\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__19002\,
            I => \receive_module.rx_counter.n3519\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18999\,
            I => \N__18995\
        );

    \I__4061\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18992\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__18995\,
            I => \N__18989\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__18992\,
            I => \receive_module.rx_counter.old_VS\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__18989\,
            I => \receive_module.rx_counter.old_VS\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__18984\,
            I => \receive_module.rx_counter.n11_cascade_\
        );

    \I__4056\ : SRMux
    port map (
            O => \N__18981\,
            I => \N__18978\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__18978\,
            I => \N__18975\
        );

    \I__4054\ : Odrv12
    port map (
            O => \N__18975\,
            I => \receive_module.rx_counter.n2547\
        );

    \I__4053\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18969\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__18969\,
            I => \receive_module.rx_counter.n11\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18963\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__18963\,
            I => \N__18960\
        );

    \I__4049\ : Span12Mux_s6_v
    port map (
            O => \N__18960\,
            I => \N__18956\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18953\
        );

    \I__4047\ : Odrv12
    port map (
            O => \N__18956\,
            I => \PULSE_1HZ\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__18953\,
            I => \PULSE_1HZ\
        );

    \I__4045\ : CEMux
    port map (
            O => \N__18948\,
            I => \N__18944\
        );

    \I__4044\ : CEMux
    port map (
            O => \N__18947\,
            I => \N__18941\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18944\,
            I => \N__18938\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__18941\,
            I => \N__18935\
        );

    \I__4041\ : Odrv4
    port map (
            O => \N__18938\,
            I => \receive_module.rx_counter.n3672\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__18935\,
            I => \receive_module.rx_counter.n3672\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18930\,
            I => \N__18926\
        );

    \I__4038\ : InMux
    port map (
            O => \N__18929\,
            I => \N__18923\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18926\,
            I => \N__18913\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__18923\,
            I => \N__18910\
        );

    \I__4035\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18903\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18903\
        );

    \I__4033\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18903\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18919\,
            I => \N__18900\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18895\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18895\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18916\,
            I => \N__18892\
        );

    \I__4028\ : Span4Mux_v
    port map (
            O => \N__18913\,
            I => \N__18889\
        );

    \I__4027\ : Span4Mux_h
    port map (
            O => \N__18910\,
            I => \N__18884\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__18903\,
            I => \N__18884\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__18900\,
            I => \RX_ADDR_12\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__18895\,
            I => \RX_ADDR_12\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__18892\,
            I => \RX_ADDR_12\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__18889\,
            I => \RX_ADDR_12\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__18884\,
            I => \RX_ADDR_12\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__18873\,
            I => \N__18868\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__18872\,
            I => \N__18863\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__18871\,
            I => \N__18860\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18868\,
            I => \N__18857\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__18867\,
            I => \N__18854\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__18866\,
            I => \N__18851\
        );

    \I__4014\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18846\
        );

    \I__4013\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18843\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__18857\,
            I => \N__18840\
        );

    \I__4011\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18835\
        );

    \I__4010\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18835\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__18850\,
            I => \N__18830\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__18849\,
            I => \N__18827\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__18846\,
            I => \N__18824\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__18843\,
            I => \N__18817\
        );

    \I__4005\ : Span4Mux_h
    port map (
            O => \N__18840\,
            I => \N__18817\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__18835\,
            I => \N__18817\
        );

    \I__4003\ : InMux
    port map (
            O => \N__18834\,
            I => \N__18814\
        );

    \I__4002\ : InMux
    port map (
            O => \N__18833\,
            I => \N__18809\
        );

    \I__4001\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18809\
        );

    \I__4000\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18806\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__18824\,
            I => \N__18803\
        );

    \I__3998\ : Span4Mux_v
    port map (
            O => \N__18817\,
            I => \N__18800\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__18814\,
            I => \RX_ADDR_13\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__18809\,
            I => \RX_ADDR_13\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__18806\,
            I => \RX_ADDR_13\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__18803\,
            I => \RX_ADDR_13\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__18800\,
            I => \RX_ADDR_13\
        );

    \I__3992\ : InMux
    port map (
            O => \N__18789\,
            I => \N__18785\
        );

    \I__3991\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18782\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__18785\,
            I => \N__18773\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__18782\,
            I => \N__18770\
        );

    \I__3988\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18763\
        );

    \I__3987\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18763\
        );

    \I__3986\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18763\
        );

    \I__3985\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18759\
        );

    \I__3984\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18754\
        );

    \I__3983\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18754\
        );

    \I__3982\ : Span4Mux_v
    port map (
            O => \N__18773\,
            I => \N__18751\
        );

    \I__3981\ : Span4Mux_h
    port map (
            O => \N__18770\,
            I => \N__18748\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__18763\,
            I => \N__18745\
        );

    \I__3979\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18742\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__18759\,
            I => \RX_ADDR_11\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__18754\,
            I => \RX_ADDR_11\
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__18751\,
            I => \RX_ADDR_11\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__18748\,
            I => \RX_ADDR_11\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__18745\,
            I => \RX_ADDR_11\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__18742\,
            I => \RX_ADDR_11\
        );

    \I__3972\ : SRMux
    port map (
            O => \N__18729\,
            I => \N__18726\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18722\
        );

    \I__3970\ : SRMux
    port map (
            O => \N__18725\,
            I => \N__18719\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__18722\,
            I => \N__18712\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18712\
        );

    \I__3967\ : SRMux
    port map (
            O => \N__18718\,
            I => \N__18709\
        );

    \I__3966\ : SRMux
    port map (
            O => \N__18717\,
            I => \N__18706\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__18712\,
            I => \N__18699\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__18709\,
            I => \N__18699\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18699\
        );

    \I__3962\ : Span4Mux_v
    port map (
            O => \N__18699\,
            I => \N__18696\
        );

    \I__3961\ : Span4Mux_h
    port map (
            O => \N__18696\,
            I => \N__18693\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__18693\,
            I => \line_buffer.n538\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18690\,
            I => \N__18687\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__18687\,
            I => \N__18683\
        );

    \I__3957\ : InMux
    port map (
            O => \N__18686\,
            I => \N__18680\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__18683\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__18680\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__3954\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18672\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__18672\,
            I => \N__18669\
        );

    \I__3952\ : Span4Mux_h
    port map (
            O => \N__18669\,
            I => \N__18666\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__18666\,
            I => \transmit_module.X_DELTA_PATTERN_15\
        );

    \I__3950\ : CEMux
    port map (
            O => \N__18663\,
            I => \N__18659\
        );

    \I__3949\ : CEMux
    port map (
            O => \N__18662\,
            I => \N__18656\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__18659\,
            I => \N__18652\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__18656\,
            I => \N__18649\
        );

    \I__3946\ : CEMux
    port map (
            O => \N__18655\,
            I => \N__18646\
        );

    \I__3945\ : Span4Mux_v
    port map (
            O => \N__18652\,
            I => \N__18642\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__18649\,
            I => \N__18639\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__18646\,
            I => \N__18636\
        );

    \I__3942\ : CEMux
    port map (
            O => \N__18645\,
            I => \N__18633\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__18642\,
            I => \transmit_module.n2084\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__18639\,
            I => \transmit_module.n2084\
        );

    \I__3939\ : Odrv12
    port map (
            O => \N__18636\,
            I => \transmit_module.n2084\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__18633\,
            I => \transmit_module.n2084\
        );

    \I__3937\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18618\
        );

    \I__3936\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18613\
        );

    \I__3935\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18613\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18610\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__18618\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__18613\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__18610\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18603\,
            I => \bfn_17_9_0_\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__18600\,
            I => \N__18596\
        );

    \I__3928\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18591\
        );

    \I__3927\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18588\
        );

    \I__3926\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18583\
        );

    \I__3925\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18583\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__18591\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__18588\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__18583\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__3921\ : InMux
    port map (
            O => \N__18576\,
            I => \receive_module.rx_counter.n3172\
        );

    \I__3920\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18567\
        );

    \I__3919\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18562\
        );

    \I__3918\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18562\
        );

    \I__3917\ : InMux
    port map (
            O => \N__18570\,
            I => \N__18559\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__18567\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__18562\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__18559\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__3913\ : InMux
    port map (
            O => \N__18552\,
            I => \receive_module.rx_counter.n3173\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__18549\,
            I => \N__18546\
        );

    \I__3911\ : InMux
    port map (
            O => \N__18546\,
            I => \N__18540\
        );

    \I__3910\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18537\
        );

    \I__3909\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18532\
        );

    \I__3908\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18532\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__18540\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__18537\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__18532\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__3904\ : InMux
    port map (
            O => \N__18525\,
            I => \receive_module.rx_counter.n3174\
        );

    \I__3903\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18516\
        );

    \I__3902\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18509\
        );

    \I__3901\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18509\
        );

    \I__3900\ : InMux
    port map (
            O => \N__18519\,
            I => \N__18509\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__18516\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__18509\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__3897\ : InMux
    port map (
            O => \N__18504\,
            I => \receive_module.rx_counter.n3175\
        );

    \I__3896\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18496\
        );

    \I__3895\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18491\
        );

    \I__3894\ : InMux
    port map (
            O => \N__18499\,
            I => \N__18491\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__18496\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__18491\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__3891\ : InMux
    port map (
            O => \N__18486\,
            I => \receive_module.rx_counter.n3176\
        );

    \I__3890\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18478\
        );

    \I__3889\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18475\
        );

    \I__3888\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18472\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__18478\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__18475\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__18472\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__3884\ : InMux
    port map (
            O => \N__18465\,
            I => \receive_module.rx_counter.n3177\
        );

    \I__3883\ : InMux
    port map (
            O => \N__18462\,
            I => \N__18456\
        );

    \I__3882\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18451\
        );

    \I__3881\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18451\
        );

    \I__3880\ : InMux
    port map (
            O => \N__18459\,
            I => \N__18448\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__18456\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__18451\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__18448\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__3876\ : InMux
    port map (
            O => \N__18441\,
            I => \receive_module.rx_counter.n3178\
        );

    \I__3875\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18435\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__18435\,
            I => \N__18432\
        );

    \I__3873\ : Span4Mux_v
    port map (
            O => \N__18432\,
            I => \N__18429\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__18429\,
            I => \N__18426\
        );

    \I__3871\ : Span4Mux_h
    port map (
            O => \N__18426\,
            I => \N__18423\
        );

    \I__3870\ : Sp12to4
    port map (
            O => \N__18423\,
            I => \N__18420\
        );

    \I__3869\ : Span12Mux_v
    port map (
            O => \N__18420\,
            I => \N__18417\
        );

    \I__3868\ : Odrv12
    port map (
            O => \N__18417\,
            I => \line_buffer.n532\
        );

    \I__3867\ : CascadeMux
    port map (
            O => \N__18414\,
            I => \N__18411\
        );

    \I__3866\ : InMux
    port map (
            O => \N__18411\,
            I => \N__18408\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__18408\,
            I => \N__18405\
        );

    \I__3864\ : Span4Mux_v
    port map (
            O => \N__18405\,
            I => \N__18402\
        );

    \I__3863\ : Sp12to4
    port map (
            O => \N__18402\,
            I => \N__18399\
        );

    \I__3862\ : Span12Mux_v
    port map (
            O => \N__18399\,
            I => \N__18396\
        );

    \I__3861\ : Odrv12
    port map (
            O => \N__18396\,
            I => \line_buffer.n524\
        );

    \I__3860\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18390\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__18390\,
            I => \N__18387\
        );

    \I__3858\ : Sp12to4
    port map (
            O => \N__18387\,
            I => \N__18384\
        );

    \I__3857\ : Odrv12
    port map (
            O => \N__18384\,
            I => \line_buffer.n467\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__18381\,
            I => \N__18378\
        );

    \I__3855\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18375\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__18375\,
            I => \N__18372\
        );

    \I__3853\ : Span4Mux_v
    port map (
            O => \N__18372\,
            I => \N__18369\
        );

    \I__3852\ : Sp12to4
    port map (
            O => \N__18369\,
            I => \N__18366\
        );

    \I__3851\ : Span12Mux_h
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__3850\ : Odrv12
    port map (
            O => \N__18363\,
            I => \line_buffer.n459\
        );

    \I__3849\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18357\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__18357\,
            I => \line_buffer.n3587\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__18354\,
            I => \line_buffer.n3590_cascade_\
        );

    \I__3846\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18348\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__18348\,
            I => \line_buffer.n3626\
        );

    \I__3844\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18342\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__18342\,
            I => \TX_DATA_3\
        );

    \I__3842\ : IoInMux
    port map (
            O => \N__18339\,
            I => \N__18334\
        );

    \I__3841\ : IoInMux
    port map (
            O => \N__18338\,
            I => \N__18331\
        );

    \I__3840\ : IoInMux
    port map (
            O => \N__18337\,
            I => \N__18328\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__18334\,
            I => \N__18325\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__18331\,
            I => \N__18322\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__18328\,
            I => \N__18319\
        );

    \I__3836\ : IoSpan4Mux
    port map (
            O => \N__18325\,
            I => \N__18316\
        );

    \I__3835\ : IoSpan4Mux
    port map (
            O => \N__18322\,
            I => \N__18313\
        );

    \I__3834\ : Span4Mux_s3_h
    port map (
            O => \N__18319\,
            I => \N__18310\
        );

    \I__3833\ : Span4Mux_s3_v
    port map (
            O => \N__18316\,
            I => \N__18307\
        );

    \I__3832\ : Span4Mux_s3_v
    port map (
            O => \N__18313\,
            I => \N__18304\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__18310\,
            I => \N__18301\
        );

    \I__3830\ : Sp12to4
    port map (
            O => \N__18307\,
            I => \N__18298\
        );

    \I__3829\ : Sp12to4
    port map (
            O => \N__18304\,
            I => \N__18295\
        );

    \I__3828\ : Span4Mux_h
    port map (
            O => \N__18301\,
            I => \N__18292\
        );

    \I__3827\ : Span12Mux_s10_v
    port map (
            O => \N__18298\,
            I => \N__18289\
        );

    \I__3826\ : Span12Mux_h
    port map (
            O => \N__18295\,
            I => \N__18286\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__18292\,
            I => \N__18283\
        );

    \I__3824\ : Odrv12
    port map (
            O => \N__18289\,
            I => n1815
        );

    \I__3823\ : Odrv12
    port map (
            O => \N__18286\,
            I => n1815
        );

    \I__3822\ : Odrv4
    port map (
            O => \N__18283\,
            I => n1815
        );

    \I__3821\ : SRMux
    port map (
            O => \N__18276\,
            I => \N__18272\
        );

    \I__3820\ : SRMux
    port map (
            O => \N__18275\,
            I => \N__18267\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__18272\,
            I => \N__18264\
        );

    \I__3818\ : SRMux
    port map (
            O => \N__18271\,
            I => \N__18261\
        );

    \I__3817\ : SRMux
    port map (
            O => \N__18270\,
            I => \N__18258\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__18267\,
            I => \N__18255\
        );

    \I__3815\ : Span4Mux_s2_v
    port map (
            O => \N__18264\,
            I => \N__18248\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__18261\,
            I => \N__18248\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__18258\,
            I => \N__18248\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__18255\,
            I => \N__18245\
        );

    \I__3811\ : Span4Mux_v
    port map (
            O => \N__18248\,
            I => \N__18242\
        );

    \I__3810\ : Span4Mux_v
    port map (
            O => \N__18245\,
            I => \N__18239\
        );

    \I__3809\ : Span4Mux_h
    port map (
            O => \N__18242\,
            I => \N__18236\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__18239\,
            I => \N__18233\
        );

    \I__3807\ : Span4Mux_h
    port map (
            O => \N__18236\,
            I => \N__18230\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__18233\,
            I => \line_buffer.n602\
        );

    \I__3805\ : Odrv4
    port map (
            O => \N__18230\,
            I => \line_buffer.n602\
        );

    \I__3804\ : IoInMux
    port map (
            O => \N__18225\,
            I => \N__18222\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__18222\,
            I => \N__18219\
        );

    \I__3802\ : IoSpan4Mux
    port map (
            O => \N__18219\,
            I => \N__18216\
        );

    \I__3801\ : Span4Mux_s2_h
    port map (
            O => \N__18216\,
            I => \N__18212\
        );

    \I__3800\ : IoInMux
    port map (
            O => \N__18215\,
            I => \N__18209\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__18212\,
            I => \N__18206\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18203\
        );

    \I__3797\ : Sp12to4
    port map (
            O => \N__18206\,
            I => \N__18200\
        );

    \I__3796\ : IoSpan4Mux
    port map (
            O => \N__18203\,
            I => \N__18197\
        );

    \I__3795\ : Span12Mux_h
    port map (
            O => \N__18200\,
            I => \N__18194\
        );

    \I__3794\ : Span4Mux_s3_v
    port map (
            O => \N__18197\,
            I => \N__18191\
        );

    \I__3793\ : Odrv12
    port map (
            O => \N__18194\,
            I => \GB_BUFFER_DEBUG_c_3_c_THRU_CO\
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__18191\,
            I => \GB_BUFFER_DEBUG_c_3_c_THRU_CO\
        );

    \I__3791\ : IoInMux
    port map (
            O => \N__18186\,
            I => \N__18183\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__18183\,
            I => \N__18180\
        );

    \I__3789\ : IoSpan4Mux
    port map (
            O => \N__18180\,
            I => \N__18177\
        );

    \I__3788\ : Span4Mux_s3_h
    port map (
            O => \N__18177\,
            I => \N__18173\
        );

    \I__3787\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18170\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__18173\,
            I => \N__18167\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__18170\,
            I => \N__18164\
        );

    \I__3784\ : Span4Mux_h
    port map (
            O => \N__18167\,
            I => \N__18160\
        );

    \I__3783\ : Span4Mux_h
    port map (
            O => \N__18164\,
            I => \N__18157\
        );

    \I__3782\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18154\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__18160\,
            I => \DEBUG_c_0\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__18157\,
            I => \DEBUG_c_0\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__18154\,
            I => \DEBUG_c_0\
        );

    \I__3778\ : IoInMux
    port map (
            O => \N__18147\,
            I => \N__18144\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__3776\ : Span4Mux_s3_v
    port map (
            O => \N__18141\,
            I => \N__18138\
        );

    \I__3775\ : Span4Mux_h
    port map (
            O => \N__18138\,
            I => \N__18135\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__18135\,
            I => \LED_c\
        );

    \I__3773\ : InMux
    port map (
            O => \N__18132\,
            I => \N__18129\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__18129\,
            I => \N__18126\
        );

    \I__3771\ : Sp12to4
    port map (
            O => \N__18126\,
            I => \N__18123\
        );

    \I__3770\ : Span12Mux_v
    port map (
            O => \N__18123\,
            I => \N__18120\
        );

    \I__3769\ : Span12Mux_h
    port map (
            O => \N__18120\,
            I => \N__18117\
        );

    \I__3768\ : Odrv12
    port map (
            O => \N__18117\,
            I => \TVP_VIDEO_c_2\
        );

    \I__3767\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18111\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__18111\,
            I => \tvp_video_buffer.BUFFER_0_2\
        );

    \I__3765\ : SRMux
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__18105\,
            I => \N__18101\
        );

    \I__3763\ : SRMux
    port map (
            O => \N__18104\,
            I => \N__18098\
        );

    \I__3762\ : Span4Mux_v
    port map (
            O => \N__18101\,
            I => \N__18092\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__18098\,
            I => \N__18092\
        );

    \I__3760\ : SRMux
    port map (
            O => \N__18097\,
            I => \N__18088\
        );

    \I__3759\ : Span4Mux_v
    port map (
            O => \N__18092\,
            I => \N__18085\
        );

    \I__3758\ : SRMux
    port map (
            O => \N__18091\,
            I => \N__18082\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__18088\,
            I => \N__18075\
        );

    \I__3756\ : Sp12to4
    port map (
            O => \N__18085\,
            I => \N__18075\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__18082\,
            I => \N__18075\
        );

    \I__3754\ : Span12Mux_v
    port map (
            O => \N__18075\,
            I => \N__18072\
        );

    \I__3753\ : Odrv12
    port map (
            O => \N__18072\,
            I => \line_buffer.n474\
        );

    \I__3752\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18066\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__18066\,
            I => \N__18063\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__18063\,
            I => \receive_module.n128\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__18060\,
            I => \N__18056\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__18059\,
            I => \N__18053\
        );

    \I__3747\ : CascadeBuf
    port map (
            O => \N__18056\,
            I => \N__18050\
        );

    \I__3746\ : CascadeBuf
    port map (
            O => \N__18053\,
            I => \N__18047\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \N__18044\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__18047\,
            I => \N__18041\
        );

    \I__3743\ : CascadeBuf
    port map (
            O => \N__18044\,
            I => \N__18038\
        );

    \I__3742\ : CascadeBuf
    port map (
            O => \N__18041\,
            I => \N__18035\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__18038\,
            I => \N__18032\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__18035\,
            I => \N__18029\
        );

    \I__3739\ : CascadeBuf
    port map (
            O => \N__18032\,
            I => \N__18026\
        );

    \I__3738\ : CascadeBuf
    port map (
            O => \N__18029\,
            I => \N__18023\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__18026\,
            I => \N__18020\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__18023\,
            I => \N__18017\
        );

    \I__3735\ : CascadeBuf
    port map (
            O => \N__18020\,
            I => \N__18014\
        );

    \I__3734\ : CascadeBuf
    port map (
            O => \N__18017\,
            I => \N__18011\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__18014\,
            I => \N__18008\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__18011\,
            I => \N__18005\
        );

    \I__3731\ : CascadeBuf
    port map (
            O => \N__18008\,
            I => \N__18002\
        );

    \I__3730\ : CascadeBuf
    port map (
            O => \N__18005\,
            I => \N__17999\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__18002\,
            I => \N__17996\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__17999\,
            I => \N__17993\
        );

    \I__3727\ : CascadeBuf
    port map (
            O => \N__17996\,
            I => \N__17990\
        );

    \I__3726\ : CascadeBuf
    port map (
            O => \N__17993\,
            I => \N__17987\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__17990\,
            I => \N__17984\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__17987\,
            I => \N__17981\
        );

    \I__3723\ : CascadeBuf
    port map (
            O => \N__17984\,
            I => \N__17978\
        );

    \I__3722\ : CascadeBuf
    port map (
            O => \N__17981\,
            I => \N__17975\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__17978\,
            I => \N__17972\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__17975\,
            I => \N__17969\
        );

    \I__3719\ : CascadeBuf
    port map (
            O => \N__17972\,
            I => \N__17966\
        );

    \I__3718\ : CascadeBuf
    port map (
            O => \N__17969\,
            I => \N__17963\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__17966\,
            I => \N__17960\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__17963\,
            I => \N__17957\
        );

    \I__3715\ : CascadeBuf
    port map (
            O => \N__17960\,
            I => \N__17954\
        );

    \I__3714\ : CascadeBuf
    port map (
            O => \N__17957\,
            I => \N__17951\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__17954\,
            I => \N__17948\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__17951\,
            I => \N__17945\
        );

    \I__3711\ : CascadeBuf
    port map (
            O => \N__17948\,
            I => \N__17942\
        );

    \I__3710\ : CascadeBuf
    port map (
            O => \N__17945\,
            I => \N__17939\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__17942\,
            I => \N__17936\
        );

    \I__3708\ : CascadeMux
    port map (
            O => \N__17939\,
            I => \N__17933\
        );

    \I__3707\ : CascadeBuf
    port map (
            O => \N__17936\,
            I => \N__17930\
        );

    \I__3706\ : CascadeBuf
    port map (
            O => \N__17933\,
            I => \N__17927\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17930\,
            I => \N__17924\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__17927\,
            I => \N__17921\
        );

    \I__3703\ : CascadeBuf
    port map (
            O => \N__17924\,
            I => \N__17918\
        );

    \I__3702\ : CascadeBuf
    port map (
            O => \N__17921\,
            I => \N__17915\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__17918\,
            I => \N__17912\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__17915\,
            I => \N__17909\
        );

    \I__3699\ : CascadeBuf
    port map (
            O => \N__17912\,
            I => \N__17906\
        );

    \I__3698\ : CascadeBuf
    port map (
            O => \N__17909\,
            I => \N__17903\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__17906\,
            I => \N__17900\
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__17903\,
            I => \N__17897\
        );

    \I__3695\ : CascadeBuf
    port map (
            O => \N__17900\,
            I => \N__17894\
        );

    \I__3694\ : CascadeBuf
    port map (
            O => \N__17897\,
            I => \N__17891\
        );

    \I__3693\ : CascadeMux
    port map (
            O => \N__17894\,
            I => \N__17888\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__17891\,
            I => \N__17885\
        );

    \I__3691\ : CascadeBuf
    port map (
            O => \N__17888\,
            I => \N__17882\
        );

    \I__3690\ : CascadeBuf
    port map (
            O => \N__17885\,
            I => \N__17879\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__17882\,
            I => \N__17876\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__17879\,
            I => \N__17873\
        );

    \I__3687\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17870\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17867\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__17870\,
            I => \N__17864\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__17867\,
            I => \N__17861\
        );

    \I__3683\ : Span4Mux_s1_v
    port map (
            O => \N__17864\,
            I => \N__17858\
        );

    \I__3682\ : Span4Mux_s1_v
    port map (
            O => \N__17861\,
            I => \N__17855\
        );

    \I__3681\ : Span4Mux_v
    port map (
            O => \N__17858\,
            I => \N__17850\
        );

    \I__3680\ : Span4Mux_v
    port map (
            O => \N__17855\,
            I => \N__17847\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__17854\,
            I => \N__17844\
        );

    \I__3678\ : InMux
    port map (
            O => \N__17853\,
            I => \N__17841\
        );

    \I__3677\ : Sp12to4
    port map (
            O => \N__17850\,
            I => \N__17838\
        );

    \I__3676\ : Sp12to4
    port map (
            O => \N__17847\,
            I => \N__17835\
        );

    \I__3675\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17832\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__17841\,
            I => \N__17829\
        );

    \I__3673\ : Span12Mux_h
    port map (
            O => \N__17838\,
            I => \N__17824\
        );

    \I__3672\ : Span12Mux_h
    port map (
            O => \N__17835\,
            I => \N__17824\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__17832\,
            I => \RX_ADDR_9\
        );

    \I__3670\ : Odrv4
    port map (
            O => \N__17829\,
            I => \RX_ADDR_9\
        );

    \I__3669\ : Odrv12
    port map (
            O => \N__17824\,
            I => \RX_ADDR_9\
        );

    \I__3668\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17814\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__17814\,
            I => \N__17811\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__17811\,
            I => \receive_module.n134\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__17808\,
            I => \N__17805\
        );

    \I__3664\ : CascadeBuf
    port map (
            O => \N__17805\,
            I => \N__17801\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__17804\,
            I => \N__17798\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__17801\,
            I => \N__17795\
        );

    \I__3661\ : CascadeBuf
    port map (
            O => \N__17798\,
            I => \N__17792\
        );

    \I__3660\ : CascadeBuf
    port map (
            O => \N__17795\,
            I => \N__17789\
        );

    \I__3659\ : CascadeMux
    port map (
            O => \N__17792\,
            I => \N__17786\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__17789\,
            I => \N__17783\
        );

    \I__3657\ : CascadeBuf
    port map (
            O => \N__17786\,
            I => \N__17780\
        );

    \I__3656\ : CascadeBuf
    port map (
            O => \N__17783\,
            I => \N__17777\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__17780\,
            I => \N__17774\
        );

    \I__3654\ : CascadeMux
    port map (
            O => \N__17777\,
            I => \N__17771\
        );

    \I__3653\ : CascadeBuf
    port map (
            O => \N__17774\,
            I => \N__17768\
        );

    \I__3652\ : CascadeBuf
    port map (
            O => \N__17771\,
            I => \N__17765\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__17768\,
            I => \N__17762\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__17765\,
            I => \N__17759\
        );

    \I__3649\ : CascadeBuf
    port map (
            O => \N__17762\,
            I => \N__17756\
        );

    \I__3648\ : CascadeBuf
    port map (
            O => \N__17759\,
            I => \N__17753\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__17756\,
            I => \N__17750\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__17753\,
            I => \N__17747\
        );

    \I__3645\ : CascadeBuf
    port map (
            O => \N__17750\,
            I => \N__17744\
        );

    \I__3644\ : CascadeBuf
    port map (
            O => \N__17747\,
            I => \N__17741\
        );

    \I__3643\ : CascadeMux
    port map (
            O => \N__17744\,
            I => \N__17738\
        );

    \I__3642\ : CascadeMux
    port map (
            O => \N__17741\,
            I => \N__17735\
        );

    \I__3641\ : CascadeBuf
    port map (
            O => \N__17738\,
            I => \N__17732\
        );

    \I__3640\ : CascadeBuf
    port map (
            O => \N__17735\,
            I => \N__17729\
        );

    \I__3639\ : CascadeMux
    port map (
            O => \N__17732\,
            I => \N__17726\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__17729\,
            I => \N__17723\
        );

    \I__3637\ : CascadeBuf
    port map (
            O => \N__17726\,
            I => \N__17720\
        );

    \I__3636\ : CascadeBuf
    port map (
            O => \N__17723\,
            I => \N__17717\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__17720\,
            I => \N__17714\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__17717\,
            I => \N__17711\
        );

    \I__3633\ : CascadeBuf
    port map (
            O => \N__17714\,
            I => \N__17708\
        );

    \I__3632\ : CascadeBuf
    port map (
            O => \N__17711\,
            I => \N__17705\
        );

    \I__3631\ : CascadeMux
    port map (
            O => \N__17708\,
            I => \N__17702\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__17705\,
            I => \N__17699\
        );

    \I__3629\ : CascadeBuf
    port map (
            O => \N__17702\,
            I => \N__17696\
        );

    \I__3628\ : CascadeBuf
    port map (
            O => \N__17699\,
            I => \N__17693\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__17696\,
            I => \N__17690\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__17693\,
            I => \N__17687\
        );

    \I__3625\ : CascadeBuf
    port map (
            O => \N__17690\,
            I => \N__17684\
        );

    \I__3624\ : CascadeBuf
    port map (
            O => \N__17687\,
            I => \N__17681\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__17684\,
            I => \N__17678\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__17681\,
            I => \N__17675\
        );

    \I__3621\ : CascadeBuf
    port map (
            O => \N__17678\,
            I => \N__17672\
        );

    \I__3620\ : CascadeBuf
    port map (
            O => \N__17675\,
            I => \N__17669\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__17672\,
            I => \N__17666\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__17669\,
            I => \N__17663\
        );

    \I__3617\ : CascadeBuf
    port map (
            O => \N__17666\,
            I => \N__17660\
        );

    \I__3616\ : CascadeBuf
    port map (
            O => \N__17663\,
            I => \N__17657\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__17660\,
            I => \N__17654\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__17657\,
            I => \N__17651\
        );

    \I__3613\ : CascadeBuf
    port map (
            O => \N__17654\,
            I => \N__17648\
        );

    \I__3612\ : CascadeBuf
    port map (
            O => \N__17651\,
            I => \N__17645\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__17648\,
            I => \N__17642\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__17645\,
            I => \N__17639\
        );

    \I__3609\ : CascadeBuf
    port map (
            O => \N__17642\,
            I => \N__17636\
        );

    \I__3608\ : CascadeBuf
    port map (
            O => \N__17639\,
            I => \N__17633\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__17636\,
            I => \N__17630\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__17633\,
            I => \N__17627\
        );

    \I__3605\ : CascadeBuf
    port map (
            O => \N__17630\,
            I => \N__17624\
        );

    \I__3604\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17621\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__17624\,
            I => \N__17618\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__17621\,
            I => \N__17614\
        );

    \I__3601\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17611\
        );

    \I__3600\ : InMux
    port map (
            O => \N__17617\,
            I => \N__17608\
        );

    \I__3599\ : Span4Mux_s2_v
    port map (
            O => \N__17614\,
            I => \N__17605\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__17611\,
            I => \N__17602\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__17608\,
            I => \N__17599\
        );

    \I__3596\ : Sp12to4
    port map (
            O => \N__17605\,
            I => \N__17595\
        );

    \I__3595\ : Sp12to4
    port map (
            O => \N__17602\,
            I => \N__17592\
        );

    \I__3594\ : Span4Mux_h
    port map (
            O => \N__17599\,
            I => \N__17589\
        );

    \I__3593\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17586\
        );

    \I__3592\ : Span12Mux_h
    port map (
            O => \N__17595\,
            I => \N__17583\
        );

    \I__3591\ : Span12Mux_v
    port map (
            O => \N__17592\,
            I => \N__17580\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__17589\,
            I => \RX_ADDR_3\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__17586\,
            I => \RX_ADDR_3\
        );

    \I__3588\ : Odrv12
    port map (
            O => \N__17583\,
            I => \RX_ADDR_3\
        );

    \I__3587\ : Odrv12
    port map (
            O => \N__17580\,
            I => \RX_ADDR_3\
        );

    \I__3586\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17568\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__17568\,
            I => \N__17565\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__17565\,
            I => \receive_module.n133\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__17562\,
            I => \N__17558\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__17561\,
            I => \N__17555\
        );

    \I__3581\ : CascadeBuf
    port map (
            O => \N__17558\,
            I => \N__17552\
        );

    \I__3580\ : CascadeBuf
    port map (
            O => \N__17555\,
            I => \N__17549\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__17552\,
            I => \N__17546\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__17549\,
            I => \N__17543\
        );

    \I__3577\ : CascadeBuf
    port map (
            O => \N__17546\,
            I => \N__17540\
        );

    \I__3576\ : CascadeBuf
    port map (
            O => \N__17543\,
            I => \N__17537\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__17540\,
            I => \N__17534\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__17537\,
            I => \N__17531\
        );

    \I__3573\ : CascadeBuf
    port map (
            O => \N__17534\,
            I => \N__17528\
        );

    \I__3572\ : CascadeBuf
    port map (
            O => \N__17531\,
            I => \N__17525\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__17528\,
            I => \N__17522\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__17525\,
            I => \N__17519\
        );

    \I__3569\ : CascadeBuf
    port map (
            O => \N__17522\,
            I => \N__17516\
        );

    \I__3568\ : CascadeBuf
    port map (
            O => \N__17519\,
            I => \N__17513\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__17516\,
            I => \N__17510\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__17513\,
            I => \N__17507\
        );

    \I__3565\ : CascadeBuf
    port map (
            O => \N__17510\,
            I => \N__17504\
        );

    \I__3564\ : CascadeBuf
    port map (
            O => \N__17507\,
            I => \N__17501\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__17504\,
            I => \N__17498\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__17501\,
            I => \N__17495\
        );

    \I__3561\ : CascadeBuf
    port map (
            O => \N__17498\,
            I => \N__17492\
        );

    \I__3560\ : CascadeBuf
    port map (
            O => \N__17495\,
            I => \N__17489\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__17492\,
            I => \N__17486\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__17489\,
            I => \N__17483\
        );

    \I__3557\ : CascadeBuf
    port map (
            O => \N__17486\,
            I => \N__17480\
        );

    \I__3556\ : CascadeBuf
    port map (
            O => \N__17483\,
            I => \N__17477\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__17480\,
            I => \N__17474\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__17477\,
            I => \N__17471\
        );

    \I__3553\ : CascadeBuf
    port map (
            O => \N__17474\,
            I => \N__17468\
        );

    \I__3552\ : CascadeBuf
    port map (
            O => \N__17471\,
            I => \N__17465\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__17468\,
            I => \N__17462\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__17465\,
            I => \N__17459\
        );

    \I__3549\ : CascadeBuf
    port map (
            O => \N__17462\,
            I => \N__17456\
        );

    \I__3548\ : CascadeBuf
    port map (
            O => \N__17459\,
            I => \N__17453\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__17456\,
            I => \N__17450\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__17453\,
            I => \N__17447\
        );

    \I__3545\ : CascadeBuf
    port map (
            O => \N__17450\,
            I => \N__17444\
        );

    \I__3544\ : CascadeBuf
    port map (
            O => \N__17447\,
            I => \N__17441\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__17444\,
            I => \N__17438\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__17441\,
            I => \N__17435\
        );

    \I__3541\ : CascadeBuf
    port map (
            O => \N__17438\,
            I => \N__17432\
        );

    \I__3540\ : CascadeBuf
    port map (
            O => \N__17435\,
            I => \N__17429\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__17432\,
            I => \N__17426\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__17429\,
            I => \N__17423\
        );

    \I__3537\ : CascadeBuf
    port map (
            O => \N__17426\,
            I => \N__17420\
        );

    \I__3536\ : CascadeBuf
    port map (
            O => \N__17423\,
            I => \N__17417\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__17420\,
            I => \N__17414\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__17417\,
            I => \N__17411\
        );

    \I__3533\ : CascadeBuf
    port map (
            O => \N__17414\,
            I => \N__17408\
        );

    \I__3532\ : CascadeBuf
    port map (
            O => \N__17411\,
            I => \N__17405\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__17408\,
            I => \N__17402\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__17405\,
            I => \N__17399\
        );

    \I__3529\ : CascadeBuf
    port map (
            O => \N__17402\,
            I => \N__17396\
        );

    \I__3528\ : CascadeBuf
    port map (
            O => \N__17399\,
            I => \N__17393\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__17396\,
            I => \N__17390\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__17393\,
            I => \N__17387\
        );

    \I__3525\ : CascadeBuf
    port map (
            O => \N__17390\,
            I => \N__17384\
        );

    \I__3524\ : CascadeBuf
    port map (
            O => \N__17387\,
            I => \N__17381\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__17384\,
            I => \N__17378\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__17381\,
            I => \N__17375\
        );

    \I__3521\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17372\
        );

    \I__3520\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17369\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__17372\,
            I => \N__17366\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__17369\,
            I => \N__17363\
        );

    \I__3517\ : Span4Mux_s1_v
    port map (
            O => \N__17366\,
            I => \N__17358\
        );

    \I__3516\ : Span4Mux_s1_v
    port map (
            O => \N__17363\,
            I => \N__17355\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__17362\,
            I => \N__17352\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__17361\,
            I => \N__17349\
        );

    \I__3513\ : Sp12to4
    port map (
            O => \N__17358\,
            I => \N__17346\
        );

    \I__3512\ : Sp12to4
    port map (
            O => \N__17355\,
            I => \N__17343\
        );

    \I__3511\ : InMux
    port map (
            O => \N__17352\,
            I => \N__17340\
        );

    \I__3510\ : InMux
    port map (
            O => \N__17349\,
            I => \N__17337\
        );

    \I__3509\ : Span12Mux_h
    port map (
            O => \N__17346\,
            I => \N__17332\
        );

    \I__3508\ : Span12Mux_h
    port map (
            O => \N__17343\,
            I => \N__17332\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__17340\,
            I => \N__17329\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__17337\,
            I => \N__17324\
        );

    \I__3505\ : Span12Mux_v
    port map (
            O => \N__17332\,
            I => \N__17324\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__17329\,
            I => \RX_ADDR_4\
        );

    \I__3503\ : Odrv12
    port map (
            O => \N__17324\,
            I => \RX_ADDR_4\
        );

    \I__3502\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17316\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__17316\,
            I => \N__17313\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__17313\,
            I => \receive_module.n129\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__17310\,
            I => \N__17306\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__17309\,
            I => \N__17303\
        );

    \I__3497\ : CascadeBuf
    port map (
            O => \N__17306\,
            I => \N__17300\
        );

    \I__3496\ : CascadeBuf
    port map (
            O => \N__17303\,
            I => \N__17297\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__17300\,
            I => \N__17294\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__17297\,
            I => \N__17291\
        );

    \I__3493\ : CascadeBuf
    port map (
            O => \N__17294\,
            I => \N__17288\
        );

    \I__3492\ : CascadeBuf
    port map (
            O => \N__17291\,
            I => \N__17285\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__17288\,
            I => \N__17282\
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__17285\,
            I => \N__17279\
        );

    \I__3489\ : CascadeBuf
    port map (
            O => \N__17282\,
            I => \N__17276\
        );

    \I__3488\ : CascadeBuf
    port map (
            O => \N__17279\,
            I => \N__17273\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__17276\,
            I => \N__17270\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__17273\,
            I => \N__17267\
        );

    \I__3485\ : CascadeBuf
    port map (
            O => \N__17270\,
            I => \N__17264\
        );

    \I__3484\ : CascadeBuf
    port map (
            O => \N__17267\,
            I => \N__17261\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__17264\,
            I => \N__17258\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__17261\,
            I => \N__17255\
        );

    \I__3481\ : CascadeBuf
    port map (
            O => \N__17258\,
            I => \N__17252\
        );

    \I__3480\ : CascadeBuf
    port map (
            O => \N__17255\,
            I => \N__17249\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__17252\,
            I => \N__17246\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__17249\,
            I => \N__17243\
        );

    \I__3477\ : CascadeBuf
    port map (
            O => \N__17246\,
            I => \N__17240\
        );

    \I__3476\ : CascadeBuf
    port map (
            O => \N__17243\,
            I => \N__17237\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__17240\,
            I => \N__17234\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__17237\,
            I => \N__17231\
        );

    \I__3473\ : CascadeBuf
    port map (
            O => \N__17234\,
            I => \N__17228\
        );

    \I__3472\ : CascadeBuf
    port map (
            O => \N__17231\,
            I => \N__17225\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__17228\,
            I => \N__17222\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__17225\,
            I => \N__17219\
        );

    \I__3469\ : CascadeBuf
    port map (
            O => \N__17222\,
            I => \N__17216\
        );

    \I__3468\ : CascadeBuf
    port map (
            O => \N__17219\,
            I => \N__17213\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__17216\,
            I => \N__17210\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__17213\,
            I => \N__17207\
        );

    \I__3465\ : CascadeBuf
    port map (
            O => \N__17210\,
            I => \N__17204\
        );

    \I__3464\ : CascadeBuf
    port map (
            O => \N__17207\,
            I => \N__17201\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__17204\,
            I => \N__17198\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__17201\,
            I => \N__17195\
        );

    \I__3461\ : CascadeBuf
    port map (
            O => \N__17198\,
            I => \N__17192\
        );

    \I__3460\ : CascadeBuf
    port map (
            O => \N__17195\,
            I => \N__17189\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__17192\,
            I => \N__17186\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__17189\,
            I => \N__17183\
        );

    \I__3457\ : CascadeBuf
    port map (
            O => \N__17186\,
            I => \N__17180\
        );

    \I__3456\ : CascadeBuf
    port map (
            O => \N__17183\,
            I => \N__17177\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__17180\,
            I => \N__17174\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__17177\,
            I => \N__17171\
        );

    \I__3453\ : CascadeBuf
    port map (
            O => \N__17174\,
            I => \N__17168\
        );

    \I__3452\ : CascadeBuf
    port map (
            O => \N__17171\,
            I => \N__17165\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__17168\,
            I => \N__17162\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__17165\,
            I => \N__17159\
        );

    \I__3449\ : CascadeBuf
    port map (
            O => \N__17162\,
            I => \N__17156\
        );

    \I__3448\ : CascadeBuf
    port map (
            O => \N__17159\,
            I => \N__17153\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__17156\,
            I => \N__17150\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__17153\,
            I => \N__17147\
        );

    \I__3445\ : CascadeBuf
    port map (
            O => \N__17150\,
            I => \N__17144\
        );

    \I__3444\ : CascadeBuf
    port map (
            O => \N__17147\,
            I => \N__17141\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__17144\,
            I => \N__17138\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__17141\,
            I => \N__17135\
        );

    \I__3441\ : CascadeBuf
    port map (
            O => \N__17138\,
            I => \N__17132\
        );

    \I__3440\ : CascadeBuf
    port map (
            O => \N__17135\,
            I => \N__17129\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__17132\,
            I => \N__17126\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__17129\,
            I => \N__17123\
        );

    \I__3437\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17120\
        );

    \I__3436\ : InMux
    port map (
            O => \N__17123\,
            I => \N__17117\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__17120\,
            I => \N__17113\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__17117\,
            I => \N__17110\
        );

    \I__3433\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17107\
        );

    \I__3432\ : Span4Mux_h
    port map (
            O => \N__17113\,
            I => \N__17104\
        );

    \I__3431\ : Span4Mux_h
    port map (
            O => \N__17110\,
            I => \N__17101\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__17107\,
            I => \N__17097\
        );

    \I__3429\ : Sp12to4
    port map (
            O => \N__17104\,
            I => \N__17094\
        );

    \I__3428\ : Sp12to4
    port map (
            O => \N__17101\,
            I => \N__17091\
        );

    \I__3427\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17088\
        );

    \I__3426\ : Span12Mux_v
    port map (
            O => \N__17097\,
            I => \N__17083\
        );

    \I__3425\ : Span12Mux_v
    port map (
            O => \N__17094\,
            I => \N__17083\
        );

    \I__3424\ : Span12Mux_v
    port map (
            O => \N__17091\,
            I => \N__17080\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__17088\,
            I => \RX_ADDR_8\
        );

    \I__3422\ : Odrv12
    port map (
            O => \N__17083\,
            I => \RX_ADDR_8\
        );

    \I__3421\ : Odrv12
    port map (
            O => \N__17080\,
            I => \RX_ADDR_8\
        );

    \I__3420\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17070\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__17070\,
            I => \N__17067\
        );

    \I__3418\ : Span4Mux_h
    port map (
            O => \N__17067\,
            I => \N__17064\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__17064\,
            I => \receive_module.n131\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__17061\,
            I => \N__17057\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__17060\,
            I => \N__17054\
        );

    \I__3414\ : CascadeBuf
    port map (
            O => \N__17057\,
            I => \N__17051\
        );

    \I__3413\ : CascadeBuf
    port map (
            O => \N__17054\,
            I => \N__17048\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__17051\,
            I => \N__17045\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__17048\,
            I => \N__17042\
        );

    \I__3410\ : CascadeBuf
    port map (
            O => \N__17045\,
            I => \N__17039\
        );

    \I__3409\ : CascadeBuf
    port map (
            O => \N__17042\,
            I => \N__17036\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__17039\,
            I => \N__17033\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__17036\,
            I => \N__17030\
        );

    \I__3406\ : CascadeBuf
    port map (
            O => \N__17033\,
            I => \N__17027\
        );

    \I__3405\ : CascadeBuf
    port map (
            O => \N__17030\,
            I => \N__17024\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__17027\,
            I => \N__17021\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__17024\,
            I => \N__17018\
        );

    \I__3402\ : CascadeBuf
    port map (
            O => \N__17021\,
            I => \N__17015\
        );

    \I__3401\ : CascadeBuf
    port map (
            O => \N__17018\,
            I => \N__17012\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__17015\,
            I => \N__17009\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__17012\,
            I => \N__17006\
        );

    \I__3398\ : CascadeBuf
    port map (
            O => \N__17009\,
            I => \N__17003\
        );

    \I__3397\ : CascadeBuf
    port map (
            O => \N__17006\,
            I => \N__17000\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__17003\,
            I => \N__16997\
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__17000\,
            I => \N__16994\
        );

    \I__3394\ : CascadeBuf
    port map (
            O => \N__16997\,
            I => \N__16991\
        );

    \I__3393\ : CascadeBuf
    port map (
            O => \N__16994\,
            I => \N__16988\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__16991\,
            I => \N__16985\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__16988\,
            I => \N__16982\
        );

    \I__3390\ : CascadeBuf
    port map (
            O => \N__16985\,
            I => \N__16979\
        );

    \I__3389\ : CascadeBuf
    port map (
            O => \N__16982\,
            I => \N__16976\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__16979\,
            I => \N__16973\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__16976\,
            I => \N__16970\
        );

    \I__3386\ : CascadeBuf
    port map (
            O => \N__16973\,
            I => \N__16967\
        );

    \I__3385\ : CascadeBuf
    port map (
            O => \N__16970\,
            I => \N__16964\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__16967\,
            I => \N__16961\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__16964\,
            I => \N__16958\
        );

    \I__3382\ : CascadeBuf
    port map (
            O => \N__16961\,
            I => \N__16955\
        );

    \I__3381\ : CascadeBuf
    port map (
            O => \N__16958\,
            I => \N__16952\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__16955\,
            I => \N__16949\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__16952\,
            I => \N__16946\
        );

    \I__3378\ : CascadeBuf
    port map (
            O => \N__16949\,
            I => \N__16943\
        );

    \I__3377\ : CascadeBuf
    port map (
            O => \N__16946\,
            I => \N__16940\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__16943\,
            I => \N__16937\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__16940\,
            I => \N__16934\
        );

    \I__3374\ : CascadeBuf
    port map (
            O => \N__16937\,
            I => \N__16931\
        );

    \I__3373\ : CascadeBuf
    port map (
            O => \N__16934\,
            I => \N__16928\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__16931\,
            I => \N__16925\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__16928\,
            I => \N__16922\
        );

    \I__3370\ : CascadeBuf
    port map (
            O => \N__16925\,
            I => \N__16919\
        );

    \I__3369\ : CascadeBuf
    port map (
            O => \N__16922\,
            I => \N__16916\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__16919\,
            I => \N__16913\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__16916\,
            I => \N__16910\
        );

    \I__3366\ : CascadeBuf
    port map (
            O => \N__16913\,
            I => \N__16907\
        );

    \I__3365\ : CascadeBuf
    port map (
            O => \N__16910\,
            I => \N__16904\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__16907\,
            I => \N__16901\
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__16904\,
            I => \N__16898\
        );

    \I__3362\ : CascadeBuf
    port map (
            O => \N__16901\,
            I => \N__16895\
        );

    \I__3361\ : CascadeBuf
    port map (
            O => \N__16898\,
            I => \N__16892\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__16895\,
            I => \N__16889\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__16892\,
            I => \N__16886\
        );

    \I__3358\ : CascadeBuf
    port map (
            O => \N__16889\,
            I => \N__16883\
        );

    \I__3357\ : CascadeBuf
    port map (
            O => \N__16886\,
            I => \N__16880\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__16883\,
            I => \N__16877\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__16880\,
            I => \N__16874\
        );

    \I__3354\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16871\
        );

    \I__3353\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16868\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__16871\,
            I => \N__16865\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__16868\,
            I => \N__16861\
        );

    \I__3350\ : Span4Mux_s1_v
    port map (
            O => \N__16865\,
            I => \N__16858\
        );

    \I__3349\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16854\
        );

    \I__3348\ : Span4Mux_s1_v
    port map (
            O => \N__16861\,
            I => \N__16851\
        );

    \I__3347\ : Sp12to4
    port map (
            O => \N__16858\,
            I => \N__16848\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__16857\,
            I => \N__16845\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16854\,
            I => \N__16842\
        );

    \I__3344\ : Sp12to4
    port map (
            O => \N__16851\,
            I => \N__16839\
        );

    \I__3343\ : Span12Mux_h
    port map (
            O => \N__16848\,
            I => \N__16836\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16833\
        );

    \I__3341\ : Span4Mux_h
    port map (
            O => \N__16842\,
            I => \N__16830\
        );

    \I__3340\ : Span12Mux_v
    port map (
            O => \N__16839\,
            I => \N__16825\
        );

    \I__3339\ : Span12Mux_v
    port map (
            O => \N__16836\,
            I => \N__16825\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__16833\,
            I => \RX_ADDR_6\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__16830\,
            I => \RX_ADDR_6\
        );

    \I__3336\ : Odrv12
    port map (
            O => \N__16825\,
            I => \RX_ADDR_6\
        );

    \I__3335\ : InMux
    port map (
            O => \N__16818\,
            I => \N__16815\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__16815\,
            I => \N__16812\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__16812\,
            I => \receive_module.n130\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__16809\,
            I => \N__16805\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__16808\,
            I => \N__16802\
        );

    \I__3330\ : CascadeBuf
    port map (
            O => \N__16805\,
            I => \N__16799\
        );

    \I__3329\ : CascadeBuf
    port map (
            O => \N__16802\,
            I => \N__16796\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__16799\,
            I => \N__16793\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__16796\,
            I => \N__16790\
        );

    \I__3326\ : CascadeBuf
    port map (
            O => \N__16793\,
            I => \N__16787\
        );

    \I__3325\ : CascadeBuf
    port map (
            O => \N__16790\,
            I => \N__16784\
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__16787\,
            I => \N__16781\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__16784\,
            I => \N__16778\
        );

    \I__3322\ : CascadeBuf
    port map (
            O => \N__16781\,
            I => \N__16775\
        );

    \I__3321\ : CascadeBuf
    port map (
            O => \N__16778\,
            I => \N__16772\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__16775\,
            I => \N__16769\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__16772\,
            I => \N__16766\
        );

    \I__3318\ : CascadeBuf
    port map (
            O => \N__16769\,
            I => \N__16763\
        );

    \I__3317\ : CascadeBuf
    port map (
            O => \N__16766\,
            I => \N__16760\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__16763\,
            I => \N__16757\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__16760\,
            I => \N__16754\
        );

    \I__3314\ : CascadeBuf
    port map (
            O => \N__16757\,
            I => \N__16751\
        );

    \I__3313\ : CascadeBuf
    port map (
            O => \N__16754\,
            I => \N__16748\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__16751\,
            I => \N__16745\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__16748\,
            I => \N__16742\
        );

    \I__3310\ : CascadeBuf
    port map (
            O => \N__16745\,
            I => \N__16739\
        );

    \I__3309\ : CascadeBuf
    port map (
            O => \N__16742\,
            I => \N__16736\
        );

    \I__3308\ : CascadeMux
    port map (
            O => \N__16739\,
            I => \N__16733\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__16736\,
            I => \N__16730\
        );

    \I__3306\ : CascadeBuf
    port map (
            O => \N__16733\,
            I => \N__16727\
        );

    \I__3305\ : CascadeBuf
    port map (
            O => \N__16730\,
            I => \N__16724\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__16727\,
            I => \N__16721\
        );

    \I__3303\ : CascadeMux
    port map (
            O => \N__16724\,
            I => \N__16718\
        );

    \I__3302\ : CascadeBuf
    port map (
            O => \N__16721\,
            I => \N__16715\
        );

    \I__3301\ : CascadeBuf
    port map (
            O => \N__16718\,
            I => \N__16712\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__16715\,
            I => \N__16709\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__16712\,
            I => \N__16706\
        );

    \I__3298\ : CascadeBuf
    port map (
            O => \N__16709\,
            I => \N__16703\
        );

    \I__3297\ : CascadeBuf
    port map (
            O => \N__16706\,
            I => \N__16700\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__16703\,
            I => \N__16697\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__16700\,
            I => \N__16694\
        );

    \I__3294\ : CascadeBuf
    port map (
            O => \N__16697\,
            I => \N__16691\
        );

    \I__3293\ : CascadeBuf
    port map (
            O => \N__16694\,
            I => \N__16688\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__16691\,
            I => \N__16685\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__16688\,
            I => \N__16682\
        );

    \I__3290\ : CascadeBuf
    port map (
            O => \N__16685\,
            I => \N__16679\
        );

    \I__3289\ : CascadeBuf
    port map (
            O => \N__16682\,
            I => \N__16676\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__16679\,
            I => \N__16673\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__16676\,
            I => \N__16670\
        );

    \I__3286\ : CascadeBuf
    port map (
            O => \N__16673\,
            I => \N__16667\
        );

    \I__3285\ : CascadeBuf
    port map (
            O => \N__16670\,
            I => \N__16664\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__16667\,
            I => \N__16661\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__16664\,
            I => \N__16658\
        );

    \I__3282\ : CascadeBuf
    port map (
            O => \N__16661\,
            I => \N__16655\
        );

    \I__3281\ : CascadeBuf
    port map (
            O => \N__16658\,
            I => \N__16652\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__16655\,
            I => \N__16649\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__16652\,
            I => \N__16646\
        );

    \I__3278\ : CascadeBuf
    port map (
            O => \N__16649\,
            I => \N__16643\
        );

    \I__3277\ : CascadeBuf
    port map (
            O => \N__16646\,
            I => \N__16640\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__16643\,
            I => \N__16637\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__16640\,
            I => \N__16634\
        );

    \I__3274\ : CascadeBuf
    port map (
            O => \N__16637\,
            I => \N__16631\
        );

    \I__3273\ : CascadeBuf
    port map (
            O => \N__16634\,
            I => \N__16628\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__16631\,
            I => \N__16625\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__16628\,
            I => \N__16622\
        );

    \I__3270\ : InMux
    port map (
            O => \N__16625\,
            I => \N__16619\
        );

    \I__3269\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16615\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__16619\,
            I => \N__16612\
        );

    \I__3267\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16609\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__16615\,
            I => \N__16606\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__16612\,
            I => \N__16603\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__16609\,
            I => \N__16600\
        );

    \I__3263\ : Span12Mux_s1_v
    port map (
            O => \N__16606\,
            I => \N__16596\
        );

    \I__3262\ : Sp12to4
    port map (
            O => \N__16603\,
            I => \N__16593\
        );

    \I__3261\ : Span4Mux_h
    port map (
            O => \N__16600\,
            I => \N__16590\
        );

    \I__3260\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16587\
        );

    \I__3259\ : Span12Mux_v
    port map (
            O => \N__16596\,
            I => \N__16584\
        );

    \I__3258\ : Span12Mux_v
    port map (
            O => \N__16593\,
            I => \N__16581\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__16590\,
            I => \RX_ADDR_7\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__16587\,
            I => \RX_ADDR_7\
        );

    \I__3255\ : Odrv12
    port map (
            O => \N__16584\,
            I => \RX_ADDR_7\
        );

    \I__3254\ : Odrv12
    port map (
            O => \N__16581\,
            I => \RX_ADDR_7\
        );

    \I__3253\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16569\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16566\
        );

    \I__3251\ : Span4Mux_v
    port map (
            O => \N__16566\,
            I => \N__16563\
        );

    \I__3250\ : Span4Mux_h
    port map (
            O => \N__16563\,
            I => \N__16560\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__16560\,
            I => \N__16557\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__16557\,
            I => \N__16554\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__16554\,
            I => \line_buffer.n564\
        );

    \I__3246\ : InMux
    port map (
            O => \N__16551\,
            I => \N__16548\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16545\
        );

    \I__3244\ : Span4Mux_v
    port map (
            O => \N__16545\,
            I => \N__16542\
        );

    \I__3243\ : Span4Mux_h
    port map (
            O => \N__16542\,
            I => \N__16539\
        );

    \I__3242\ : Span4Mux_h
    port map (
            O => \N__16539\,
            I => \N__16536\
        );

    \I__3241\ : Odrv4
    port map (
            O => \N__16536\,
            I => \line_buffer.n556\
        );

    \I__3240\ : SRMux
    port map (
            O => \N__16533\,
            I => \N__16529\
        );

    \I__3239\ : SRMux
    port map (
            O => \N__16532\,
            I => \N__16524\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__16529\,
            I => \N__16521\
        );

    \I__3237\ : SRMux
    port map (
            O => \N__16528\,
            I => \N__16518\
        );

    \I__3236\ : SRMux
    port map (
            O => \N__16527\,
            I => \N__16515\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__16524\,
            I => \N__16512\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__16521\,
            I => \N__16509\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__16518\,
            I => \N__16506\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__16515\,
            I => \N__16503\
        );

    \I__3231\ : Span4Mux_h
    port map (
            O => \N__16512\,
            I => \N__16500\
        );

    \I__3230\ : Span4Mux_h
    port map (
            O => \N__16509\,
            I => \N__16497\
        );

    \I__3229\ : Span4Mux_h
    port map (
            O => \N__16506\,
            I => \N__16492\
        );

    \I__3228\ : Span4Mux_v
    port map (
            O => \N__16503\,
            I => \N__16492\
        );

    \I__3227\ : Sp12to4
    port map (
            O => \N__16500\,
            I => \N__16489\
        );

    \I__3226\ : Sp12to4
    port map (
            O => \N__16497\,
            I => \N__16486\
        );

    \I__3225\ : Sp12to4
    port map (
            O => \N__16492\,
            I => \N__16481\
        );

    \I__3224\ : Span12Mux_s5_v
    port map (
            O => \N__16489\,
            I => \N__16481\
        );

    \I__3223\ : Span12Mux_v
    port map (
            O => \N__16486\,
            I => \N__16476\
        );

    \I__3222\ : Span12Mux_v
    port map (
            O => \N__16481\,
            I => \N__16476\
        );

    \I__3221\ : Odrv12
    port map (
            O => \N__16476\,
            I => \line_buffer.n473\
        );

    \I__3220\ : SRMux
    port map (
            O => \N__16473\,
            I => \N__16470\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__16470\,
            I => \N__16467\
        );

    \I__3218\ : Span4Mux_v
    port map (
            O => \N__16467\,
            I => \N__16461\
        );

    \I__3217\ : SRMux
    port map (
            O => \N__16466\,
            I => \N__16458\
        );

    \I__3216\ : SRMux
    port map (
            O => \N__16465\,
            I => \N__16455\
        );

    \I__3215\ : SRMux
    port map (
            O => \N__16464\,
            I => \N__16452\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__16461\,
            I => \N__16447\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__16458\,
            I => \N__16447\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__16455\,
            I => \N__16442\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__16452\,
            I => \N__16442\
        );

    \I__3210\ : Span4Mux_v
    port map (
            O => \N__16447\,
            I => \N__16437\
        );

    \I__3209\ : Span4Mux_v
    port map (
            O => \N__16442\,
            I => \N__16437\
        );

    \I__3208\ : Span4Mux_h
    port map (
            O => \N__16437\,
            I => \N__16434\
        );

    \I__3207\ : Span4Mux_h
    port map (
            O => \N__16434\,
            I => \N__16431\
        );

    \I__3206\ : Odrv4
    port map (
            O => \N__16431\,
            I => \line_buffer.n570\
        );

    \I__3205\ : SRMux
    port map (
            O => \N__16428\,
            I => \N__16424\
        );

    \I__3204\ : SRMux
    port map (
            O => \N__16427\,
            I => \N__16420\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__16424\,
            I => \N__16417\
        );

    \I__3202\ : SRMux
    port map (
            O => \N__16423\,
            I => \N__16414\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__16420\,
            I => \N__16410\
        );

    \I__3200\ : Span4Mux_h
    port map (
            O => \N__16417\,
            I => \N__16405\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__16414\,
            I => \N__16405\
        );

    \I__3198\ : SRMux
    port map (
            O => \N__16413\,
            I => \N__16402\
        );

    \I__3197\ : Span4Mux_v
    port map (
            O => \N__16410\,
            I => \N__16399\
        );

    \I__3196\ : Span4Mux_v
    port map (
            O => \N__16405\,
            I => \N__16394\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__16402\,
            I => \N__16394\
        );

    \I__3194\ : Sp12to4
    port map (
            O => \N__16399\,
            I => \N__16391\
        );

    \I__3193\ : Span4Mux_h
    port map (
            O => \N__16394\,
            I => \N__16388\
        );

    \I__3192\ : Span12Mux_h
    port map (
            O => \N__16391\,
            I => \N__16385\
        );

    \I__3191\ : Span4Mux_h
    port map (
            O => \N__16388\,
            I => \N__16382\
        );

    \I__3190\ : Odrv12
    port map (
            O => \N__16385\,
            I => \line_buffer.n571\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__16382\,
            I => \line_buffer.n571\
        );

    \I__3188\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16374\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__16374\,
            I => \N__16371\
        );

    \I__3186\ : Span4Mux_h
    port map (
            O => \N__16371\,
            I => \N__16368\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__16368\,
            I => \transmit_module.ADDR_Y_COMPONENT_11\
        );

    \I__3184\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16362\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__16362\,
            I => \N__16359\
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__16359\,
            I => \transmit_module.n121\
        );

    \I__3181\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16353\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__16353\,
            I => \N__16350\
        );

    \I__3179\ : Span4Mux_h
    port map (
            O => \N__16350\,
            I => \N__16347\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__16347\,
            I => \transmit_module.ADDR_Y_COMPONENT_13\
        );

    \I__3177\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16341\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__16341\,
            I => \N__16338\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__16338\,
            I => \transmit_module.n119\
        );

    \I__3174\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16332\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__16332\,
            I => \N__16329\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__16329\,
            I => \N__16326\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__16326\,
            I => \transmit_module.ADDR_Y_COMPONENT_12\
        );

    \I__3170\ : InMux
    port map (
            O => \N__16323\,
            I => \N__16309\
        );

    \I__3169\ : InMux
    port map (
            O => \N__16322\,
            I => \N__16309\
        );

    \I__3168\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16301\
        );

    \I__3167\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16291\
        );

    \I__3166\ : InMux
    port map (
            O => \N__16319\,
            I => \N__16291\
        );

    \I__3165\ : InMux
    port map (
            O => \N__16318\,
            I => \N__16291\
        );

    \I__3164\ : InMux
    port map (
            O => \N__16317\,
            I => \N__16282\
        );

    \I__3163\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16282\
        );

    \I__3162\ : InMux
    port map (
            O => \N__16315\,
            I => \N__16282\
        );

    \I__3161\ : InMux
    port map (
            O => \N__16314\,
            I => \N__16282\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__16309\,
            I => \N__16279\
        );

    \I__3159\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16276\
        );

    \I__3158\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16267\
        );

    \I__3157\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16267\
        );

    \I__3156\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16267\
        );

    \I__3155\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16267\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__16301\,
            I => \N__16261\
        );

    \I__3153\ : InMux
    port map (
            O => \N__16300\,
            I => \N__16254\
        );

    \I__3152\ : InMux
    port map (
            O => \N__16299\,
            I => \N__16254\
        );

    \I__3151\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16254\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__16291\,
            I => \N__16251\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__16282\,
            I => \N__16242\
        );

    \I__3148\ : Span4Mux_v
    port map (
            O => \N__16279\,
            I => \N__16242\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__16276\,
            I => \N__16242\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__16267\,
            I => \N__16242\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__16266\,
            I => \N__16234\
        );

    \I__3144\ : InMux
    port map (
            O => \N__16265\,
            I => \N__16230\
        );

    \I__3143\ : InMux
    port map (
            O => \N__16264\,
            I => \N__16227\
        );

    \I__3142\ : Sp12to4
    port map (
            O => \N__16261\,
            I => \N__16222\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__16254\,
            I => \N__16222\
        );

    \I__3140\ : Span4Mux_v
    port map (
            O => \N__16251\,
            I => \N__16217\
        );

    \I__3139\ : Span4Mux_v
    port map (
            O => \N__16242\,
            I => \N__16217\
        );

    \I__3138\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16210\
        );

    \I__3137\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16210\
        );

    \I__3136\ : InMux
    port map (
            O => \N__16239\,
            I => \N__16210\
        );

    \I__3135\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16201\
        );

    \I__3134\ : InMux
    port map (
            O => \N__16237\,
            I => \N__16201\
        );

    \I__3133\ : InMux
    port map (
            O => \N__16234\,
            I => \N__16201\
        );

    \I__3132\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16201\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__16230\,
            I => \transmit_module.n3675\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__16227\,
            I => \transmit_module.n3675\
        );

    \I__3129\ : Odrv12
    port map (
            O => \N__16222\,
            I => \transmit_module.n3675\
        );

    \I__3128\ : Odrv4
    port map (
            O => \N__16217\,
            I => \transmit_module.n3675\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__16210\,
            I => \transmit_module.n3675\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__16201\,
            I => \transmit_module.n3675\
        );

    \I__3125\ : InMux
    port map (
            O => \N__16188\,
            I => \N__16185\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__16185\,
            I => \N__16182\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__16182\,
            I => \transmit_module.n120\
        );

    \I__3122\ : CEMux
    port map (
            O => \N__16179\,
            I => \N__16176\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__16176\,
            I => \N__16173\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__16173\,
            I => \N__16170\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__16170\,
            I => \N__16167\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__16167\,
            I => \transmit_module.n2070\
        );

    \I__3117\ : CEMux
    port map (
            O => \N__16164\,
            I => \N__16161\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__16161\,
            I => \N__16158\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__16158\,
            I => \N__16155\
        );

    \I__3114\ : Odrv4
    port map (
            O => \N__16155\,
            I => \receive_module.n3671\
        );

    \I__3113\ : SRMux
    port map (
            O => \N__16152\,
            I => \N__16149\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__16149\,
            I => \N__16145\
        );

    \I__3111\ : SRMux
    port map (
            O => \N__16148\,
            I => \N__16142\
        );

    \I__3110\ : Span4Mux_v
    port map (
            O => \N__16145\,
            I => \N__16135\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__16142\,
            I => \N__16135\
        );

    \I__3108\ : SRMux
    port map (
            O => \N__16141\,
            I => \N__16132\
        );

    \I__3107\ : SRMux
    port map (
            O => \N__16140\,
            I => \N__16129\
        );

    \I__3106\ : Span4Mux_v
    port map (
            O => \N__16135\,
            I => \N__16124\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__16132\,
            I => \N__16124\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__16129\,
            I => \N__16121\
        );

    \I__3103\ : Span4Mux_h
    port map (
            O => \N__16124\,
            I => \N__16118\
        );

    \I__3102\ : Span4Mux_h
    port map (
            O => \N__16121\,
            I => \N__16115\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__16118\,
            I => \N__16112\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__16115\,
            I => \N__16107\
        );

    \I__3099\ : Span4Mux_h
    port map (
            O => \N__16112\,
            I => \N__16107\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__16107\,
            I => \line_buffer.n603\
        );

    \I__3097\ : SRMux
    port map (
            O => \N__16104\,
            I => \N__16100\
        );

    \I__3096\ : SRMux
    port map (
            O => \N__16103\,
            I => \N__16097\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__16100\,
            I => \N__16091\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__16097\,
            I => \N__16091\
        );

    \I__3093\ : SRMux
    port map (
            O => \N__16096\,
            I => \N__16088\
        );

    \I__3092\ : Span4Mux_v
    port map (
            O => \N__16091\,
            I => \N__16082\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__16088\,
            I => \N__16082\
        );

    \I__3090\ : SRMux
    port map (
            O => \N__16087\,
            I => \N__16079\
        );

    \I__3089\ : Span4Mux_v
    port map (
            O => \N__16082\,
            I => \N__16076\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__16079\,
            I => \N__16073\
        );

    \I__3087\ : Span4Mux_v
    port map (
            O => \N__16076\,
            I => \N__16070\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__16073\,
            I => \N__16067\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__16070\,
            I => \N__16064\
        );

    \I__3084\ : Span4Mux_h
    port map (
            O => \N__16067\,
            I => \N__16061\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__16064\,
            I => \N__16058\
        );

    \I__3082\ : Span4Mux_h
    port map (
            O => \N__16061\,
            I => \N__16055\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__16058\,
            I => \line_buffer.n539\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__16055\,
            I => \line_buffer.n539\
        );

    \I__3079\ : InMux
    port map (
            O => \N__16050\,
            I => \receive_module.rx_counter.n3205\
        );

    \I__3078\ : InMux
    port map (
            O => \N__16047\,
            I => \receive_module.rx_counter.n3206\
        );

    \I__3077\ : InMux
    port map (
            O => \N__16044\,
            I => \N__16041\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__16041\,
            I => \receive_module.rx_counter.n6\
        );

    \I__3075\ : InMux
    port map (
            O => \N__16038\,
            I => \N__16035\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__16035\,
            I => \receive_module.rx_counter.n7\
        );

    \I__3073\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16028\
        );

    \I__3072\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16025\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__16028\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__16025\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__3069\ : InMux
    port map (
            O => \N__16020\,
            I => \N__16016\
        );

    \I__3068\ : InMux
    port map (
            O => \N__16019\,
            I => \N__16013\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__16016\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__16013\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__3065\ : InMux
    port map (
            O => \N__16008\,
            I => \N__16005\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__16005\,
            I => \N__16000\
        );

    \I__3063\ : InMux
    port map (
            O => \N__16004\,
            I => \N__15997\
        );

    \I__3062\ : InMux
    port map (
            O => \N__16003\,
            I => \N__15994\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__16000\,
            I => \N__15991\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__15997\,
            I => \N__15988\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__15994\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__15991\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__15988\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15978\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__15978\,
            I => \N__15973\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15970\
        );

    \I__3053\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15967\
        );

    \I__3052\ : Span4Mux_v
    port map (
            O => \N__15973\,
            I => \N__15964\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__15970\,
            I => \N__15961\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15967\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__15964\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__15961\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__15954\,
            I => \N__15951\
        );

    \I__3046\ : InMux
    port map (
            O => \N__15951\,
            I => \N__15947\
        );

    \I__3045\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15943\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15940\
        );

    \I__3043\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15937\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15943\,
            I => \N__15934\
        );

    \I__3041\ : Span4Mux_v
    port map (
            O => \N__15940\,
            I => \N__15931\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15937\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__15934\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__15931\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__3037\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15920\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15917\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__15920\,
            I => \N__15912\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__15917\,
            I => \N__15912\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__15912\,
            I => \receive_module.rx_counter.n3222\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__15909\,
            I => \N__15905\
        );

    \I__3031\ : InMux
    port map (
            O => \N__15908\,
            I => \N__15902\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15905\,
            I => \N__15898\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15902\,
            I => \N__15895\
        );

    \I__3028\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15892\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__15898\,
            I => \N__15889\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__15895\,
            I => \N__15886\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__15892\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__15889\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__3023\ : Odrv4
    port map (
            O => \N__15886\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__15879\,
            I => \receive_module.rx_counter.n3455_cascade_\
        );

    \I__3021\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15873\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__15873\,
            I => \N__15868\
        );

    \I__3019\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15865\
        );

    \I__3018\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15862\
        );

    \I__3017\ : Span4Mux_v
    port map (
            O => \N__15868\,
            I => \N__15859\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__15865\,
            I => \N__15856\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__15862\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__15859\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__15856\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__3012\ : InMux
    port map (
            O => \N__15849\,
            I => \N__15843\
        );

    \I__3011\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15843\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__15843\,
            I => \N__15839\
        );

    \I__3009\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15836\
        );

    \I__3008\ : Span4Mux_v
    port map (
            O => \N__15839\,
            I => \N__15833\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__15836\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__3006\ : Odrv4
    port map (
            O => \N__15833\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15825\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__15825\,
            I => \N__15821\
        );

    \I__3003\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15818\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__15821\,
            I => \N__15815\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__15818\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__15815\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__15810\,
            I => \receive_module.rx_counter.n39_cascade_\
        );

    \I__2998\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15804\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__15804\,
            I => \receive_module.rx_counter.n3426\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15801\,
            I => \N__15798\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__15798\,
            I => \N__15795\
        );

    \I__2994\ : Odrv12
    port map (
            O => \N__15795\,
            I => \receive_module.rx_counter.n3478\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__15792\,
            I => \receive_module.rx_counter.n54_cascade_\
        );

    \I__2992\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15786\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__15786\,
            I => \N__15783\
        );

    \I__2990\ : Odrv12
    port map (
            O => \N__15783\,
            I => \receive_module.rx_counter.n4_adj_612\
        );

    \I__2989\ : InMux
    port map (
            O => \N__15780\,
            I => \N__15777\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__15777\,
            I => \N__15774\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__15774\,
            I => \receive_module.rx_counter.n4\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__15771\,
            I => \receive_module.rx_counter.n5_cascade_\
        );

    \I__2985\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15765\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__15765\,
            I => \receive_module.rx_counter.n3450\
        );

    \I__2983\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15758\
        );

    \I__2982\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15755\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__15758\,
            I => \receive_module.rx_counter.n3677\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__15755\,
            I => \receive_module.rx_counter.n3677\
        );

    \I__2979\ : SRMux
    port map (
            O => \N__15750\,
            I => \N__15747\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__15747\,
            I => \N__15743\
        );

    \I__2977\ : SRMux
    port map (
            O => \N__15746\,
            I => \N__15740\
        );

    \I__2976\ : Span4Mux_h
    port map (
            O => \N__15743\,
            I => \N__15737\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__15740\,
            I => \N__15734\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__15737\,
            I => \receive_module.rx_counter.n3\
        );

    \I__2973\ : Odrv12
    port map (
            O => \N__15734\,
            I => \receive_module.rx_counter.n3\
        );

    \I__2972\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15725\
        );

    \I__2971\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15722\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__15725\,
            I => \receive_module.rx_counter.X_1\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__15722\,
            I => \receive_module.rx_counter.X_1\
        );

    \I__2968\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15713\
        );

    \I__2967\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15710\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__15713\,
            I => \receive_module.rx_counter.X_2\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__15710\,
            I => \receive_module.rx_counter.X_2\
        );

    \I__2964\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15701\
        );

    \I__2963\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15698\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__15701\,
            I => \receive_module.rx_counter.X_0\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__15698\,
            I => \receive_module.rx_counter.X_0\
        );

    \I__2960\ : InMux
    port map (
            O => \N__15693\,
            I => \bfn_16_12_0_\
        );

    \I__2959\ : InMux
    port map (
            O => \N__15690\,
            I => \receive_module.rx_counter.n3202\
        );

    \I__2958\ : InMux
    port map (
            O => \N__15687\,
            I => \receive_module.rx_counter.n3203\
        );

    \I__2957\ : InMux
    port map (
            O => \N__15684\,
            I => \receive_module.rx_counter.n3204\
        );

    \I__2956\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15678\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__15678\,
            I => \N__15675\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__15675\,
            I => \tvp_video_buffer.BUFFER_0_5\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__15672\,
            I => \receive_module.rx_counter.n3452_cascade_\
        );

    \I__2952\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15666\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__15666\,
            I => \N__15663\
        );

    \I__2950\ : Span4Mux_v
    port map (
            O => \N__15663\,
            I => \N__15660\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__15660\,
            I => \tvp_video_buffer.BUFFER_1_5\
        );

    \I__2948\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15654\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__15654\,
            I => \N__15650\
        );

    \I__2946\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15647\
        );

    \I__2945\ : Span4Mux_s3_v
    port map (
            O => \N__15650\,
            I => \N__15644\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__15647\,
            I => \N__15641\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__15644\,
            I => \N__15637\
        );

    \I__2942\ : Span4Mux_v
    port map (
            O => \N__15641\,
            I => \N__15632\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15628\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__15637\,
            I => \N__15625\
        );

    \I__2939\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15622\
        );

    \I__2938\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15619\
        );

    \I__2937\ : Span4Mux_v
    port map (
            O => \N__15632\,
            I => \N__15616\
        );

    \I__2936\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15613\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__15628\,
            I => \N__15610\
        );

    \I__2934\ : Span4Mux_v
    port map (
            O => \N__15625\,
            I => \N__15605\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N__15605\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__15619\,
            I => \N__15602\
        );

    \I__2931\ : Sp12to4
    port map (
            O => \N__15616\,
            I => \N__15597\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__15613\,
            I => \N__15597\
        );

    \I__2929\ : Span4Mux_v
    port map (
            O => \N__15610\,
            I => \N__15594\
        );

    \I__2928\ : Span4Mux_v
    port map (
            O => \N__15605\,
            I => \N__15590\
        );

    \I__2927\ : Span4Mux_v
    port map (
            O => \N__15602\,
            I => \N__15587\
        );

    \I__2926\ : Span12Mux_h
    port map (
            O => \N__15597\,
            I => \N__15583\
        );

    \I__2925\ : Span4Mux_v
    port map (
            O => \N__15594\,
            I => \N__15580\
        );

    \I__2924\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15577\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__15590\,
            I => \N__15572\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__15587\,
            I => \N__15572\
        );

    \I__2921\ : InMux
    port map (
            O => \N__15586\,
            I => \N__15569\
        );

    \I__2920\ : Span12Mux_v
    port map (
            O => \N__15583\,
            I => \N__15562\
        );

    \I__2919\ : Sp12to4
    port map (
            O => \N__15580\,
            I => \N__15562\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__15577\,
            I => \N__15562\
        );

    \I__2917\ : Sp12to4
    port map (
            O => \N__15572\,
            I => \N__15557\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__15569\,
            I => \N__15557\
        );

    \I__2915\ : Odrv12
    port map (
            O => \N__15562\,
            I => \RX_DATA_3\
        );

    \I__2914\ : Odrv12
    port map (
            O => \N__15557\,
            I => \RX_DATA_3\
        );

    \I__2913\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15549\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__15549\,
            I => \N__15546\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__15546\,
            I => \receive_module.rx_counter.n10\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__15543\,
            I => \receive_module.rx_counter.n14_cascade_\
        );

    \I__2909\ : InMux
    port map (
            O => \N__15540\,
            I => \N__15537\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__15537\,
            I => \N__15534\
        );

    \I__2907\ : Span4Mux_h
    port map (
            O => \N__15534\,
            I => \N__15531\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__15531\,
            I => \RX_TX_SYNC\
        );

    \I__2905\ : InMux
    port map (
            O => \N__15528\,
            I => \receive_module.n3158\
        );

    \I__2904\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15521\
        );

    \I__2903\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15518\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__15521\,
            I => \N__15515\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__15518\,
            I => \N__15508\
        );

    \I__2900\ : Span4Mux_v
    port map (
            O => \N__15515\,
            I => \N__15508\
        );

    \I__2899\ : InMux
    port map (
            O => \N__15514\,
            I => \N__15505\
        );

    \I__2898\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15502\
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__15508\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__15505\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__15502\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15492\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__15492\,
            I => \transmit_module.ADDR_Y_COMPONENT_4\
        );

    \I__2892\ : InMux
    port map (
            O => \N__15489\,
            I => \N__15484\
        );

    \I__2891\ : InMux
    port map (
            O => \N__15488\,
            I => \N__15481\
        );

    \I__2890\ : InMux
    port map (
            O => \N__15487\,
            I => \N__15478\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__15484\,
            I => \N__15474\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__15481\,
            I => \N__15469\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__15478\,
            I => \N__15469\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__15477\,
            I => \N__15466\
        );

    \I__2885\ : Span4Mux_h
    port map (
            O => \N__15474\,
            I => \N__15463\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__15469\,
            I => \N__15460\
        );

    \I__2883\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15457\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__15463\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__15460\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__15457\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2879\ : InMux
    port map (
            O => \N__15450\,
            I => \N__15447\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__15447\,
            I => \transmit_module.ADDR_Y_COMPONENT_7\
        );

    \I__2877\ : InMux
    port map (
            O => \N__15444\,
            I => \N__15440\
        );

    \I__2876\ : InMux
    port map (
            O => \N__15443\,
            I => \N__15436\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__15440\,
            I => \N__15433\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__15439\,
            I => \N__15429\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__15436\,
            I => \N__15426\
        );

    \I__2872\ : Span4Mux_v
    port map (
            O => \N__15433\,
            I => \N__15423\
        );

    \I__2871\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15420\
        );

    \I__2870\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15417\
        );

    \I__2869\ : Odrv12
    port map (
            O => \N__15426\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__15423\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__15420\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__15417\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2865\ : InMux
    port map (
            O => \N__15408\,
            I => \N__15405\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__15405\,
            I => \transmit_module.ADDR_Y_COMPONENT_6\
        );

    \I__2863\ : CEMux
    port map (
            O => \N__15402\,
            I => \N__15398\
        );

    \I__2862\ : CEMux
    port map (
            O => \N__15401\,
            I => \N__15394\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__15398\,
            I => \N__15391\
        );

    \I__2860\ : CEMux
    port map (
            O => \N__15397\,
            I => \N__15385\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__15394\,
            I => \N__15382\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__15391\,
            I => \N__15379\
        );

    \I__2857\ : CEMux
    port map (
            O => \N__15390\,
            I => \N__15376\
        );

    \I__2856\ : CEMux
    port map (
            O => \N__15389\,
            I => \N__15373\
        );

    \I__2855\ : CEMux
    port map (
            O => \N__15388\,
            I => \N__15370\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15367\
        );

    \I__2853\ : Span4Mux_v
    port map (
            O => \N__15382\,
            I => \N__15364\
        );

    \I__2852\ : Span4Mux_h
    port map (
            O => \N__15379\,
            I => \N__15361\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__15376\,
            I => \N__15358\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__15373\,
            I => \N__15355\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__15370\,
            I => \N__15350\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__15367\,
            I => \N__15350\
        );

    \I__2847\ : Span4Mux_h
    port map (
            O => \N__15364\,
            I => \N__15345\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__15361\,
            I => \N__15345\
        );

    \I__2845\ : Span4Mux_v
    port map (
            O => \N__15358\,
            I => \N__15342\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__15355\,
            I => \N__15339\
        );

    \I__2843\ : Span4Mux_h
    port map (
            O => \N__15350\,
            I => \N__15336\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__15345\,
            I => \transmit_module.n2310\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__15342\,
            I => \transmit_module.n2310\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__15339\,
            I => \transmit_module.n2310\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__15336\,
            I => \transmit_module.n2310\
        );

    \I__2838\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15324\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__15324\,
            I => \N__15321\
        );

    \I__2836\ : Odrv12
    port map (
            O => \N__15321\,
            I => \receive_module.n136\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__15318\,
            I => \N__15314\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__15317\,
            I => \N__15311\
        );

    \I__2833\ : CascadeBuf
    port map (
            O => \N__15314\,
            I => \N__15308\
        );

    \I__2832\ : CascadeBuf
    port map (
            O => \N__15311\,
            I => \N__15305\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__15308\,
            I => \N__15302\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__15305\,
            I => \N__15299\
        );

    \I__2829\ : CascadeBuf
    port map (
            O => \N__15302\,
            I => \N__15296\
        );

    \I__2828\ : CascadeBuf
    port map (
            O => \N__15299\,
            I => \N__15293\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__15296\,
            I => \N__15290\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__15293\,
            I => \N__15287\
        );

    \I__2825\ : CascadeBuf
    port map (
            O => \N__15290\,
            I => \N__15284\
        );

    \I__2824\ : CascadeBuf
    port map (
            O => \N__15287\,
            I => \N__15281\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__15284\,
            I => \N__15278\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__15281\,
            I => \N__15275\
        );

    \I__2821\ : CascadeBuf
    port map (
            O => \N__15278\,
            I => \N__15272\
        );

    \I__2820\ : CascadeBuf
    port map (
            O => \N__15275\,
            I => \N__15269\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \N__15266\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__15269\,
            I => \N__15263\
        );

    \I__2817\ : CascadeBuf
    port map (
            O => \N__15266\,
            I => \N__15260\
        );

    \I__2816\ : CascadeBuf
    port map (
            O => \N__15263\,
            I => \N__15257\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__15260\,
            I => \N__15254\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \N__15251\
        );

    \I__2813\ : CascadeBuf
    port map (
            O => \N__15254\,
            I => \N__15248\
        );

    \I__2812\ : CascadeBuf
    port map (
            O => \N__15251\,
            I => \N__15245\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__15248\,
            I => \N__15242\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__15245\,
            I => \N__15239\
        );

    \I__2809\ : CascadeBuf
    port map (
            O => \N__15242\,
            I => \N__15236\
        );

    \I__2808\ : CascadeBuf
    port map (
            O => \N__15239\,
            I => \N__15233\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__15236\,
            I => \N__15230\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__15233\,
            I => \N__15227\
        );

    \I__2805\ : CascadeBuf
    port map (
            O => \N__15230\,
            I => \N__15224\
        );

    \I__2804\ : CascadeBuf
    port map (
            O => \N__15227\,
            I => \N__15221\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \N__15218\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__15221\,
            I => \N__15215\
        );

    \I__2801\ : CascadeBuf
    port map (
            O => \N__15218\,
            I => \N__15212\
        );

    \I__2800\ : CascadeBuf
    port map (
            O => \N__15215\,
            I => \N__15209\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__15212\,
            I => \N__15206\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \N__15203\
        );

    \I__2797\ : CascadeBuf
    port map (
            O => \N__15206\,
            I => \N__15200\
        );

    \I__2796\ : CascadeBuf
    port map (
            O => \N__15203\,
            I => \N__15197\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__15200\,
            I => \N__15194\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__15197\,
            I => \N__15191\
        );

    \I__2793\ : CascadeBuf
    port map (
            O => \N__15194\,
            I => \N__15188\
        );

    \I__2792\ : CascadeBuf
    port map (
            O => \N__15191\,
            I => \N__15185\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__15188\,
            I => \N__15182\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__15185\,
            I => \N__15179\
        );

    \I__2789\ : CascadeBuf
    port map (
            O => \N__15182\,
            I => \N__15176\
        );

    \I__2788\ : CascadeBuf
    port map (
            O => \N__15179\,
            I => \N__15173\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__15176\,
            I => \N__15170\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__15173\,
            I => \N__15167\
        );

    \I__2785\ : CascadeBuf
    port map (
            O => \N__15170\,
            I => \N__15164\
        );

    \I__2784\ : CascadeBuf
    port map (
            O => \N__15167\,
            I => \N__15161\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__15164\,
            I => \N__15158\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__15161\,
            I => \N__15155\
        );

    \I__2781\ : CascadeBuf
    port map (
            O => \N__15158\,
            I => \N__15152\
        );

    \I__2780\ : CascadeBuf
    port map (
            O => \N__15155\,
            I => \N__15149\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__15152\,
            I => \N__15146\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__15149\,
            I => \N__15143\
        );

    \I__2777\ : CascadeBuf
    port map (
            O => \N__15146\,
            I => \N__15140\
        );

    \I__2776\ : CascadeBuf
    port map (
            O => \N__15143\,
            I => \N__15137\
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__15140\,
            I => \N__15134\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__15137\,
            I => \N__15131\
        );

    \I__2773\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15128\
        );

    \I__2772\ : InMux
    port map (
            O => \N__15131\,
            I => \N__15125\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__15128\,
            I => \N__15120\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__15125\,
            I => \N__15117\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__15124\,
            I => \N__15114\
        );

    \I__2768\ : InMux
    port map (
            O => \N__15123\,
            I => \N__15111\
        );

    \I__2767\ : Span12Mux_h
    port map (
            O => \N__15120\,
            I => \N__15106\
        );

    \I__2766\ : Span12Mux_h
    port map (
            O => \N__15117\,
            I => \N__15106\
        );

    \I__2765\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15103\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__15111\,
            I => \N__15100\
        );

    \I__2763\ : Span12Mux_v
    port map (
            O => \N__15106\,
            I => \N__15097\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__15103\,
            I => \RX_ADDR_1\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__15100\,
            I => \RX_ADDR_1\
        );

    \I__2760\ : Odrv12
    port map (
            O => \N__15097\,
            I => \RX_ADDR_1\
        );

    \I__2759\ : InMux
    port map (
            O => \N__15090\,
            I => \N__15087\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__15087\,
            I => \N__15084\
        );

    \I__2757\ : Odrv12
    port map (
            O => \N__15084\,
            I => \receive_module.n127\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__15081\,
            I => \N__15077\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__15080\,
            I => \N__15074\
        );

    \I__2754\ : CascadeBuf
    port map (
            O => \N__15077\,
            I => \N__15071\
        );

    \I__2753\ : CascadeBuf
    port map (
            O => \N__15074\,
            I => \N__15068\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__15071\,
            I => \N__15065\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__15068\,
            I => \N__15062\
        );

    \I__2750\ : CascadeBuf
    port map (
            O => \N__15065\,
            I => \N__15059\
        );

    \I__2749\ : CascadeBuf
    port map (
            O => \N__15062\,
            I => \N__15056\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__15059\,
            I => \N__15053\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__15056\,
            I => \N__15050\
        );

    \I__2746\ : CascadeBuf
    port map (
            O => \N__15053\,
            I => \N__15047\
        );

    \I__2745\ : CascadeBuf
    port map (
            O => \N__15050\,
            I => \N__15044\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__15047\,
            I => \N__15041\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__15044\,
            I => \N__15038\
        );

    \I__2742\ : CascadeBuf
    port map (
            O => \N__15041\,
            I => \N__15035\
        );

    \I__2741\ : CascadeBuf
    port map (
            O => \N__15038\,
            I => \N__15032\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__15035\,
            I => \N__15029\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__15032\,
            I => \N__15026\
        );

    \I__2738\ : CascadeBuf
    port map (
            O => \N__15029\,
            I => \N__15023\
        );

    \I__2737\ : CascadeBuf
    port map (
            O => \N__15026\,
            I => \N__15020\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__15023\,
            I => \N__15017\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__15020\,
            I => \N__15014\
        );

    \I__2734\ : CascadeBuf
    port map (
            O => \N__15017\,
            I => \N__15011\
        );

    \I__2733\ : CascadeBuf
    port map (
            O => \N__15014\,
            I => \N__15008\
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__15011\,
            I => \N__15005\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__15008\,
            I => \N__15002\
        );

    \I__2730\ : CascadeBuf
    port map (
            O => \N__15005\,
            I => \N__14999\
        );

    \I__2729\ : CascadeBuf
    port map (
            O => \N__15002\,
            I => \N__14996\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__14999\,
            I => \N__14993\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__14996\,
            I => \N__14990\
        );

    \I__2726\ : CascadeBuf
    port map (
            O => \N__14993\,
            I => \N__14987\
        );

    \I__2725\ : CascadeBuf
    port map (
            O => \N__14990\,
            I => \N__14984\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__14987\,
            I => \N__14981\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__14984\,
            I => \N__14978\
        );

    \I__2722\ : CascadeBuf
    port map (
            O => \N__14981\,
            I => \N__14975\
        );

    \I__2721\ : CascadeBuf
    port map (
            O => \N__14978\,
            I => \N__14972\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__14975\,
            I => \N__14969\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__14972\,
            I => \N__14966\
        );

    \I__2718\ : CascadeBuf
    port map (
            O => \N__14969\,
            I => \N__14963\
        );

    \I__2717\ : CascadeBuf
    port map (
            O => \N__14966\,
            I => \N__14960\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__14963\,
            I => \N__14957\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__14960\,
            I => \N__14954\
        );

    \I__2714\ : CascadeBuf
    port map (
            O => \N__14957\,
            I => \N__14951\
        );

    \I__2713\ : CascadeBuf
    port map (
            O => \N__14954\,
            I => \N__14948\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__14951\,
            I => \N__14945\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__14948\,
            I => \N__14942\
        );

    \I__2710\ : CascadeBuf
    port map (
            O => \N__14945\,
            I => \N__14939\
        );

    \I__2709\ : CascadeBuf
    port map (
            O => \N__14942\,
            I => \N__14936\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__14939\,
            I => \N__14933\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__14936\,
            I => \N__14930\
        );

    \I__2706\ : CascadeBuf
    port map (
            O => \N__14933\,
            I => \N__14927\
        );

    \I__2705\ : CascadeBuf
    port map (
            O => \N__14930\,
            I => \N__14924\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__14927\,
            I => \N__14921\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__14924\,
            I => \N__14918\
        );

    \I__2702\ : CascadeBuf
    port map (
            O => \N__14921\,
            I => \N__14915\
        );

    \I__2701\ : CascadeBuf
    port map (
            O => \N__14918\,
            I => \N__14912\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__14915\,
            I => \N__14909\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__14912\,
            I => \N__14906\
        );

    \I__2698\ : CascadeBuf
    port map (
            O => \N__14909\,
            I => \N__14903\
        );

    \I__2697\ : CascadeBuf
    port map (
            O => \N__14906\,
            I => \N__14900\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__14903\,
            I => \N__14897\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \N__14894\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14891\
        );

    \I__2693\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14888\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14891\,
            I => \N__14885\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__14888\,
            I => \N__14882\
        );

    \I__2690\ : Span4Mux_s3_v
    port map (
            O => \N__14885\,
            I => \N__14877\
        );

    \I__2689\ : Span4Mux_s3_v
    port map (
            O => \N__14882\,
            I => \N__14874\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__14881\,
            I => \N__14871\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14880\,
            I => \N__14868\
        );

    \I__2686\ : Sp12to4
    port map (
            O => \N__14877\,
            I => \N__14865\
        );

    \I__2685\ : Sp12to4
    port map (
            O => \N__14874\,
            I => \N__14862\
        );

    \I__2684\ : InMux
    port map (
            O => \N__14871\,
            I => \N__14859\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14868\,
            I => \N__14856\
        );

    \I__2682\ : Span12Mux_h
    port map (
            O => \N__14865\,
            I => \N__14851\
        );

    \I__2681\ : Span12Mux_h
    port map (
            O => \N__14862\,
            I => \N__14851\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__14859\,
            I => \RX_ADDR_10\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__14856\,
            I => \RX_ADDR_10\
        );

    \I__2678\ : Odrv12
    port map (
            O => \N__14851\,
            I => \RX_ADDR_10\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14841\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__14841\,
            I => \N__14838\
        );

    \I__2675\ : Odrv12
    port map (
            O => \N__14838\,
            I => \receive_module.n137\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__14835\,
            I => \N__14831\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__14834\,
            I => \N__14828\
        );

    \I__2672\ : CascadeBuf
    port map (
            O => \N__14831\,
            I => \N__14825\
        );

    \I__2671\ : CascadeBuf
    port map (
            O => \N__14828\,
            I => \N__14822\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__14825\,
            I => \N__14819\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__14822\,
            I => \N__14816\
        );

    \I__2668\ : CascadeBuf
    port map (
            O => \N__14819\,
            I => \N__14813\
        );

    \I__2667\ : CascadeBuf
    port map (
            O => \N__14816\,
            I => \N__14810\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__14813\,
            I => \N__14807\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__14810\,
            I => \N__14804\
        );

    \I__2664\ : CascadeBuf
    port map (
            O => \N__14807\,
            I => \N__14801\
        );

    \I__2663\ : CascadeBuf
    port map (
            O => \N__14804\,
            I => \N__14798\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__14801\,
            I => \N__14795\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__14798\,
            I => \N__14792\
        );

    \I__2660\ : CascadeBuf
    port map (
            O => \N__14795\,
            I => \N__14789\
        );

    \I__2659\ : CascadeBuf
    port map (
            O => \N__14792\,
            I => \N__14786\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__14789\,
            I => \N__14783\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__14786\,
            I => \N__14780\
        );

    \I__2656\ : CascadeBuf
    port map (
            O => \N__14783\,
            I => \N__14777\
        );

    \I__2655\ : CascadeBuf
    port map (
            O => \N__14780\,
            I => \N__14774\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__14777\,
            I => \N__14771\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__14774\,
            I => \N__14768\
        );

    \I__2652\ : CascadeBuf
    port map (
            O => \N__14771\,
            I => \N__14765\
        );

    \I__2651\ : CascadeBuf
    port map (
            O => \N__14768\,
            I => \N__14762\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__14765\,
            I => \N__14759\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__14762\,
            I => \N__14756\
        );

    \I__2648\ : CascadeBuf
    port map (
            O => \N__14759\,
            I => \N__14753\
        );

    \I__2647\ : CascadeBuf
    port map (
            O => \N__14756\,
            I => \N__14750\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__14753\,
            I => \N__14747\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__14750\,
            I => \N__14744\
        );

    \I__2644\ : CascadeBuf
    port map (
            O => \N__14747\,
            I => \N__14741\
        );

    \I__2643\ : CascadeBuf
    port map (
            O => \N__14744\,
            I => \N__14738\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__14741\,
            I => \N__14735\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__14738\,
            I => \N__14732\
        );

    \I__2640\ : CascadeBuf
    port map (
            O => \N__14735\,
            I => \N__14729\
        );

    \I__2639\ : CascadeBuf
    port map (
            O => \N__14732\,
            I => \N__14726\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__14729\,
            I => \N__14723\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__14726\,
            I => \N__14720\
        );

    \I__2636\ : CascadeBuf
    port map (
            O => \N__14723\,
            I => \N__14717\
        );

    \I__2635\ : CascadeBuf
    port map (
            O => \N__14720\,
            I => \N__14714\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__14717\,
            I => \N__14711\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__14714\,
            I => \N__14708\
        );

    \I__2632\ : CascadeBuf
    port map (
            O => \N__14711\,
            I => \N__14705\
        );

    \I__2631\ : CascadeBuf
    port map (
            O => \N__14708\,
            I => \N__14702\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__14705\,
            I => \N__14699\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__14702\,
            I => \N__14696\
        );

    \I__2628\ : CascadeBuf
    port map (
            O => \N__14699\,
            I => \N__14693\
        );

    \I__2627\ : CascadeBuf
    port map (
            O => \N__14696\,
            I => \N__14690\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__14693\,
            I => \N__14687\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__14690\,
            I => \N__14684\
        );

    \I__2624\ : CascadeBuf
    port map (
            O => \N__14687\,
            I => \N__14681\
        );

    \I__2623\ : CascadeBuf
    port map (
            O => \N__14684\,
            I => \N__14678\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__14681\,
            I => \N__14675\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__14678\,
            I => \N__14672\
        );

    \I__2620\ : CascadeBuf
    port map (
            O => \N__14675\,
            I => \N__14669\
        );

    \I__2619\ : CascadeBuf
    port map (
            O => \N__14672\,
            I => \N__14666\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__14669\,
            I => \N__14663\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__14666\,
            I => \N__14660\
        );

    \I__2616\ : CascadeBuf
    port map (
            O => \N__14663\,
            I => \N__14657\
        );

    \I__2615\ : CascadeBuf
    port map (
            O => \N__14660\,
            I => \N__14654\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__14657\,
            I => \N__14651\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__14654\,
            I => \N__14648\
        );

    \I__2612\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14645\
        );

    \I__2611\ : InMux
    port map (
            O => \N__14648\,
            I => \N__14642\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__14645\,
            I => \N__14639\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__14642\,
            I => \N__14634\
        );

    \I__2608\ : Span4Mux_s2_v
    port map (
            O => \N__14639\,
            I => \N__14631\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__14638\,
            I => \N__14628\
        );

    \I__2606\ : InMux
    port map (
            O => \N__14637\,
            I => \N__14625\
        );

    \I__2605\ : Span12Mux_s1_v
    port map (
            O => \N__14634\,
            I => \N__14622\
        );

    \I__2604\ : Sp12to4
    port map (
            O => \N__14631\,
            I => \N__14619\
        );

    \I__2603\ : InMux
    port map (
            O => \N__14628\,
            I => \N__14616\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__14625\,
            I => \N__14613\
        );

    \I__2601\ : Span12Mux_v
    port map (
            O => \N__14622\,
            I => \N__14610\
        );

    \I__2600\ : Span12Mux_h
    port map (
            O => \N__14619\,
            I => \N__14607\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__14616\,
            I => \RX_ADDR_0\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__14613\,
            I => \RX_ADDR_0\
        );

    \I__2597\ : Odrv12
    port map (
            O => \N__14610\,
            I => \RX_ADDR_0\
        );

    \I__2596\ : Odrv12
    port map (
            O => \N__14607\,
            I => \RX_ADDR_0\
        );

    \I__2595\ : IoInMux
    port map (
            O => \N__14598\,
            I => \N__14594\
        );

    \I__2594\ : IoInMux
    port map (
            O => \N__14597\,
            I => \N__14590\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__14594\,
            I => \N__14587\
        );

    \I__2592\ : IoInMux
    port map (
            O => \N__14593\,
            I => \N__14584\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__14590\,
            I => \N__14581\
        );

    \I__2590\ : Span4Mux_s1_h
    port map (
            O => \N__14587\,
            I => \N__14578\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__14584\,
            I => \N__14575\
        );

    \I__2588\ : Sp12to4
    port map (
            O => \N__14581\,
            I => \N__14570\
        );

    \I__2587\ : Sp12to4
    port map (
            O => \N__14578\,
            I => \N__14570\
        );

    \I__2586\ : IoSpan4Mux
    port map (
            O => \N__14575\,
            I => \N__14567\
        );

    \I__2585\ : Span12Mux_v
    port map (
            O => \N__14570\,
            I => \N__14564\
        );

    \I__2584\ : Sp12to4
    port map (
            O => \N__14567\,
            I => \N__14561\
        );

    \I__2583\ : Span12Mux_h
    port map (
            O => \N__14564\,
            I => \N__14556\
        );

    \I__2582\ : Span12Mux_v
    port map (
            O => \N__14561\,
            I => \N__14556\
        );

    \I__2581\ : Odrv12
    port map (
            O => \N__14556\,
            I => n1818
        );

    \I__2580\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14550\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__14550\,
            I => \N__14547\
        );

    \I__2578\ : Span12Mux_s6_v
    port map (
            O => \N__14547\,
            I => \N__14544\
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__14544\,
            I => \receive_module.n135\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__14541\,
            I => \N__14538\
        );

    \I__2575\ : CascadeBuf
    port map (
            O => \N__14538\,
            I => \N__14534\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__14537\,
            I => \N__14531\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__14534\,
            I => \N__14528\
        );

    \I__2572\ : CascadeBuf
    port map (
            O => \N__14531\,
            I => \N__14525\
        );

    \I__2571\ : CascadeBuf
    port map (
            O => \N__14528\,
            I => \N__14522\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__14525\,
            I => \N__14519\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__14522\,
            I => \N__14516\
        );

    \I__2568\ : CascadeBuf
    port map (
            O => \N__14519\,
            I => \N__14513\
        );

    \I__2567\ : CascadeBuf
    port map (
            O => \N__14516\,
            I => \N__14510\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__14513\,
            I => \N__14507\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__14510\,
            I => \N__14504\
        );

    \I__2564\ : CascadeBuf
    port map (
            O => \N__14507\,
            I => \N__14501\
        );

    \I__2563\ : CascadeBuf
    port map (
            O => \N__14504\,
            I => \N__14498\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__14501\,
            I => \N__14495\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__14498\,
            I => \N__14492\
        );

    \I__2560\ : CascadeBuf
    port map (
            O => \N__14495\,
            I => \N__14489\
        );

    \I__2559\ : CascadeBuf
    port map (
            O => \N__14492\,
            I => \N__14486\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__14489\,
            I => \N__14483\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__14486\,
            I => \N__14480\
        );

    \I__2556\ : CascadeBuf
    port map (
            O => \N__14483\,
            I => \N__14477\
        );

    \I__2555\ : CascadeBuf
    port map (
            O => \N__14480\,
            I => \N__14474\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__14477\,
            I => \N__14471\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__14474\,
            I => \N__14468\
        );

    \I__2552\ : CascadeBuf
    port map (
            O => \N__14471\,
            I => \N__14465\
        );

    \I__2551\ : CascadeBuf
    port map (
            O => \N__14468\,
            I => \N__14462\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__14465\,
            I => \N__14459\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__14462\,
            I => \N__14456\
        );

    \I__2548\ : CascadeBuf
    port map (
            O => \N__14459\,
            I => \N__14453\
        );

    \I__2547\ : CascadeBuf
    port map (
            O => \N__14456\,
            I => \N__14450\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__14453\,
            I => \N__14447\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__14450\,
            I => \N__14444\
        );

    \I__2544\ : CascadeBuf
    port map (
            O => \N__14447\,
            I => \N__14441\
        );

    \I__2543\ : CascadeBuf
    port map (
            O => \N__14444\,
            I => \N__14438\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__14441\,
            I => \N__14435\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__14438\,
            I => \N__14432\
        );

    \I__2540\ : CascadeBuf
    port map (
            O => \N__14435\,
            I => \N__14429\
        );

    \I__2539\ : CascadeBuf
    port map (
            O => \N__14432\,
            I => \N__14426\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__14429\,
            I => \N__14423\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__14426\,
            I => \N__14420\
        );

    \I__2536\ : CascadeBuf
    port map (
            O => \N__14423\,
            I => \N__14417\
        );

    \I__2535\ : CascadeBuf
    port map (
            O => \N__14420\,
            I => \N__14414\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__14417\,
            I => \N__14411\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__14414\,
            I => \N__14408\
        );

    \I__2532\ : CascadeBuf
    port map (
            O => \N__14411\,
            I => \N__14405\
        );

    \I__2531\ : CascadeBuf
    port map (
            O => \N__14408\,
            I => \N__14402\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__14405\,
            I => \N__14399\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__14402\,
            I => \N__14396\
        );

    \I__2528\ : CascadeBuf
    port map (
            O => \N__14399\,
            I => \N__14393\
        );

    \I__2527\ : CascadeBuf
    port map (
            O => \N__14396\,
            I => \N__14390\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__14393\,
            I => \N__14387\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__14390\,
            I => \N__14384\
        );

    \I__2524\ : CascadeBuf
    port map (
            O => \N__14387\,
            I => \N__14381\
        );

    \I__2523\ : CascadeBuf
    port map (
            O => \N__14384\,
            I => \N__14378\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__14381\,
            I => \N__14375\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__14378\,
            I => \N__14372\
        );

    \I__2520\ : CascadeBuf
    port map (
            O => \N__14375\,
            I => \N__14369\
        );

    \I__2519\ : CascadeBuf
    port map (
            O => \N__14372\,
            I => \N__14366\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__14369\,
            I => \N__14363\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__14366\,
            I => \N__14360\
        );

    \I__2516\ : CascadeBuf
    port map (
            O => \N__14363\,
            I => \N__14357\
        );

    \I__2515\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14353\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__14357\,
            I => \N__14350\
        );

    \I__2513\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14347\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__14353\,
            I => \N__14344\
        );

    \I__2511\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14341\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__14347\,
            I => \N__14338\
        );

    \I__2509\ : Span4Mux_s1_v
    port map (
            O => \N__14344\,
            I => \N__14335\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__14341\,
            I => \N__14332\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__14338\,
            I => \N__14329\
        );

    \I__2506\ : Span4Mux_h
    port map (
            O => \N__14335\,
            I => \N__14325\
        );

    \I__2505\ : Span4Mux_s1_v
    port map (
            O => \N__14332\,
            I => \N__14322\
        );

    \I__2504\ : Sp12to4
    port map (
            O => \N__14329\,
            I => \N__14319\
        );

    \I__2503\ : InMux
    port map (
            O => \N__14328\,
            I => \N__14316\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__14325\,
            I => \N__14313\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__14322\,
            I => \N__14310\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__14319\,
            I => \RX_ADDR_2\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__14316\,
            I => \RX_ADDR_2\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__14313\,
            I => \RX_ADDR_2\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__14310\,
            I => \RX_ADDR_2\
        );

    \I__2496\ : InMux
    port map (
            O => \N__14301\,
            I => \receive_module.n3149\
        );

    \I__2495\ : InMux
    port map (
            O => \N__14298\,
            I => \receive_module.n3150\
        );

    \I__2494\ : InMux
    port map (
            O => \N__14295\,
            I => \receive_module.n3151\
        );

    \I__2493\ : InMux
    port map (
            O => \N__14292\,
            I => \receive_module.n3152\
        );

    \I__2492\ : InMux
    port map (
            O => \N__14289\,
            I => \bfn_15_17_0_\
        );

    \I__2491\ : InMux
    port map (
            O => \N__14286\,
            I => \receive_module.n3154\
        );

    \I__2490\ : InMux
    port map (
            O => \N__14283\,
            I => \receive_module.n3155\
        );

    \I__2489\ : InMux
    port map (
            O => \N__14280\,
            I => \receive_module.n3156\
        );

    \I__2488\ : InMux
    port map (
            O => \N__14277\,
            I => \receive_module.n3157\
        );

    \I__2487\ : InMux
    port map (
            O => \N__14274\,
            I => \N__14271\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__14271\,
            I => \transmit_module.n132\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__14268\,
            I => \transmit_module.n147_cascade_\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__14265\,
            I => \N__14262\
        );

    \I__2483\ : CascadeBuf
    port map (
            O => \N__14262\,
            I => \N__14259\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__14259\,
            I => \N__14255\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__14258\,
            I => \N__14252\
        );

    \I__2480\ : CascadeBuf
    port map (
            O => \N__14255\,
            I => \N__14249\
        );

    \I__2479\ : CascadeBuf
    port map (
            O => \N__14252\,
            I => \N__14246\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__14249\,
            I => \N__14243\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__14246\,
            I => \N__14240\
        );

    \I__2476\ : CascadeBuf
    port map (
            O => \N__14243\,
            I => \N__14237\
        );

    \I__2475\ : CascadeBuf
    port map (
            O => \N__14240\,
            I => \N__14234\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__14237\,
            I => \N__14231\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__14234\,
            I => \N__14228\
        );

    \I__2472\ : CascadeBuf
    port map (
            O => \N__14231\,
            I => \N__14225\
        );

    \I__2471\ : CascadeBuf
    port map (
            O => \N__14228\,
            I => \N__14222\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__14225\,
            I => \N__14219\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__14222\,
            I => \N__14216\
        );

    \I__2468\ : CascadeBuf
    port map (
            O => \N__14219\,
            I => \N__14213\
        );

    \I__2467\ : CascadeBuf
    port map (
            O => \N__14216\,
            I => \N__14210\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__14213\,
            I => \N__14207\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__14210\,
            I => \N__14204\
        );

    \I__2464\ : CascadeBuf
    port map (
            O => \N__14207\,
            I => \N__14201\
        );

    \I__2463\ : CascadeBuf
    port map (
            O => \N__14204\,
            I => \N__14198\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__14201\,
            I => \N__14195\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__14198\,
            I => \N__14192\
        );

    \I__2460\ : CascadeBuf
    port map (
            O => \N__14195\,
            I => \N__14189\
        );

    \I__2459\ : CascadeBuf
    port map (
            O => \N__14192\,
            I => \N__14186\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__14189\,
            I => \N__14183\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__14186\,
            I => \N__14180\
        );

    \I__2456\ : CascadeBuf
    port map (
            O => \N__14183\,
            I => \N__14177\
        );

    \I__2455\ : CascadeBuf
    port map (
            O => \N__14180\,
            I => \N__14174\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__14177\,
            I => \N__14171\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__14174\,
            I => \N__14168\
        );

    \I__2452\ : CascadeBuf
    port map (
            O => \N__14171\,
            I => \N__14165\
        );

    \I__2451\ : CascadeBuf
    port map (
            O => \N__14168\,
            I => \N__14162\
        );

    \I__2450\ : CascadeMux
    port map (
            O => \N__14165\,
            I => \N__14159\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__14162\,
            I => \N__14156\
        );

    \I__2448\ : CascadeBuf
    port map (
            O => \N__14159\,
            I => \N__14153\
        );

    \I__2447\ : CascadeBuf
    port map (
            O => \N__14156\,
            I => \N__14150\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__14153\,
            I => \N__14147\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__14150\,
            I => \N__14144\
        );

    \I__2444\ : CascadeBuf
    port map (
            O => \N__14147\,
            I => \N__14141\
        );

    \I__2443\ : CascadeBuf
    port map (
            O => \N__14144\,
            I => \N__14138\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__14141\,
            I => \N__14135\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__14138\,
            I => \N__14132\
        );

    \I__2440\ : CascadeBuf
    port map (
            O => \N__14135\,
            I => \N__14129\
        );

    \I__2439\ : CascadeBuf
    port map (
            O => \N__14132\,
            I => \N__14126\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__14129\,
            I => \N__14123\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__14126\,
            I => \N__14120\
        );

    \I__2436\ : CascadeBuf
    port map (
            O => \N__14123\,
            I => \N__14117\
        );

    \I__2435\ : CascadeBuf
    port map (
            O => \N__14120\,
            I => \N__14114\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__14117\,
            I => \N__14111\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__14114\,
            I => \N__14108\
        );

    \I__2432\ : CascadeBuf
    port map (
            O => \N__14111\,
            I => \N__14105\
        );

    \I__2431\ : CascadeBuf
    port map (
            O => \N__14108\,
            I => \N__14102\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__14105\,
            I => \N__14099\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__14102\,
            I => \N__14096\
        );

    \I__2428\ : CascadeBuf
    port map (
            O => \N__14099\,
            I => \N__14093\
        );

    \I__2427\ : CascadeBuf
    port map (
            O => \N__14096\,
            I => \N__14090\
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__14093\,
            I => \N__14087\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__14090\,
            I => \N__14084\
        );

    \I__2424\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14081\
        );

    \I__2423\ : CascadeBuf
    port map (
            O => \N__14084\,
            I => \N__14078\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__14081\,
            I => \N__14075\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__14078\,
            I => \N__14072\
        );

    \I__2420\ : Span4Mux_s2_v
    port map (
            O => \N__14075\,
            I => \N__14069\
        );

    \I__2419\ : InMux
    port map (
            O => \N__14072\,
            I => \N__14066\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__14069\,
            I => \N__14063\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__14066\,
            I => \N__14060\
        );

    \I__2416\ : Sp12to4
    port map (
            O => \N__14063\,
            I => \N__14057\
        );

    \I__2415\ : Span12Mux_s5_v
    port map (
            O => \N__14060\,
            I => \N__14054\
        );

    \I__2414\ : Span12Mux_h
    port map (
            O => \N__14057\,
            I => \N__14051\
        );

    \I__2413\ : Span12Mux_v
    port map (
            O => \N__14054\,
            I => \N__14048\
        );

    \I__2412\ : Odrv12
    port map (
            O => \N__14051\,
            I => n28
        );

    \I__2411\ : Odrv12
    port map (
            O => \N__14048\,
            I => n28
        );

    \I__2410\ : InMux
    port map (
            O => \N__14043\,
            I => \N__14036\
        );

    \I__2409\ : InMux
    port map (
            O => \N__14042\,
            I => \N__14033\
        );

    \I__2408\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14030\
        );

    \I__2407\ : InMux
    port map (
            O => \N__14040\,
            I => \N__14021\
        );

    \I__2406\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14018\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__14036\,
            I => \N__14011\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__14033\,
            I => \N__14011\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__14030\,
            I => \N__14011\
        );

    \I__2402\ : InMux
    port map (
            O => \N__14029\,
            I => \N__14006\
        );

    \I__2401\ : InMux
    port map (
            O => \N__14028\,
            I => \N__14006\
        );

    \I__2400\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14003\
        );

    \I__2399\ : InMux
    port map (
            O => \N__14026\,
            I => \N__13995\
        );

    \I__2398\ : InMux
    port map (
            O => \N__14025\,
            I => \N__13995\
        );

    \I__2397\ : InMux
    port map (
            O => \N__14024\,
            I => \N__13992\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__14021\,
            I => \N__13987\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__14018\,
            I => \N__13987\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__14011\,
            I => \N__13980\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__14006\,
            I => \N__13980\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__14003\,
            I => \N__13980\
        );

    \I__2391\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13973\
        );

    \I__2390\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13973\
        );

    \I__2389\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13973\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__13995\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__13992\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2386\ : Odrv12
    port map (
            O => \N__13987\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__13980\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__13973\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13959\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13959\,
            I => \transmit_module.n128\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13956\,
            I => \N__13953\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13953\,
            I => \N__13950\
        );

    \I__2379\ : Span4Mux_v
    port map (
            O => \N__13950\,
            I => \N__13947\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__13947\,
            I => \transmit_module.n143\
        );

    \I__2377\ : InMux
    port map (
            O => \N__13944\,
            I => \N__13941\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__13941\,
            I => \N__13938\
        );

    \I__2375\ : Span4Mux_h
    port map (
            O => \N__13938\,
            I => \N__13935\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__13935\,
            I => \transmit_module.n112\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__13932\,
            I => \transmit_module.n143_cascade_\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13923\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13923\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__13923\,
            I => \transmit_module.n116\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13920\,
            I => \N__13917\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__13917\,
            I => \transmit_module.n147\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13914\,
            I => \N__13910\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__13913\,
            I => \N__13905\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13910\,
            I => \N__13902\
        );

    \I__2364\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13899\
        );

    \I__2363\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13896\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13905\,
            I => \N__13893\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__13902\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__13899\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__13896\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13893\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13884\,
            I => \bfn_15_16_0_\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13881\,
            I => \receive_module.n3146\
        );

    \I__2355\ : InMux
    port map (
            O => \N__13878\,
            I => \receive_module.n3147\
        );

    \I__2354\ : InMux
    port map (
            O => \N__13875\,
            I => \receive_module.n3148\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13872\,
            I => \N__13869\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__13869\,
            I => \transmit_module.X_DELTA_PATTERN_8\
        );

    \I__2351\ : InMux
    port map (
            O => \N__13866\,
            I => \N__13863\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__13863\,
            I => \N__13860\
        );

    \I__2349\ : Span4Mux_v
    port map (
            O => \N__13860\,
            I => \N__13857\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__13857\,
            I => \transmit_module.X_DELTA_PATTERN_7\
        );

    \I__2347\ : InMux
    port map (
            O => \N__13854\,
            I => \N__13851\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13851\,
            I => \N__13848\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__13848\,
            I => \transmit_module.X_DELTA_PATTERN_3\
        );

    \I__2344\ : InMux
    port map (
            O => \N__13845\,
            I => \N__13842\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__13842\,
            I => \transmit_module.X_DELTA_PATTERN_9\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13836\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13836\,
            I => \transmit_module.X_DELTA_PATTERN_10\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13830\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__13830\,
            I => \N__13827\
        );

    \I__2338\ : Span4Mux_v
    port map (
            O => \N__13827\,
            I => \N__13824\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__13824\,
            I => \transmit_module.X_DELTA_PATTERN_12\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13821\,
            I => \N__13818\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__13818\,
            I => \transmit_module.X_DELTA_PATTERN_11\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13812\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__13812\,
            I => \transmit_module.X_DELTA_PATTERN_2\
        );

    \I__2332\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13806\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__13806\,
            I => \transmit_module.X_DELTA_PATTERN_1\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13800\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13800\,
            I => \transmit_module.n126\
        );

    \I__2328\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13794\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__13794\,
            I => \N__13791\
        );

    \I__2326\ : Span4Mux_v
    port map (
            O => \N__13791\,
            I => \N__13788\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__13788\,
            I => \transmit_module.n141\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__13785\,
            I => \transmit_module.n141_cascade_\
        );

    \I__2323\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13779\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13779\,
            I => \N__13775\
        );

    \I__2321\ : InMux
    port map (
            O => \N__13778\,
            I => \N__13772\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__13775\,
            I => \transmit_module.n110\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__13772\,
            I => \transmit_module.n110\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13767\,
            I => \N__13764\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13764\,
            I => \N__13761\
        );

    \I__2316\ : Odrv12
    port map (
            O => \N__13761\,
            I => \tvp_vs_buffer.BUFFER_2_0\
        );

    \I__2315\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13754\
        );

    \I__2314\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13750\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__13754\,
            I => \N__13747\
        );

    \I__2312\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13744\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__13750\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__2310\ : Odrv4
    port map (
            O => \N__13747\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__13744\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__2308\ : InMux
    port map (
            O => \N__13737\,
            I => \N__13733\
        );

    \I__2307\ : InMux
    port map (
            O => \N__13736\,
            I => \N__13730\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__13733\,
            I => \N__13724\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__13730\,
            I => \N__13724\
        );

    \I__2304\ : InMux
    port map (
            O => \N__13729\,
            I => \N__13721\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__13724\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__13721\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13713\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__13713\,
            I => \transmit_module.video_signal_controller.n3461\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13706\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13703\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__13706\,
            I => \transmit_module.video_signal_controller.n3375\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__13703\,
            I => \transmit_module.video_signal_controller.n3375\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__13698\,
            I => \transmit_module.video_signal_controller.n3673_cascade_\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13695\,
            I => \N__13691\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13687\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__13691\,
            I => \N__13684\
        );

    \I__2291\ : InMux
    port map (
            O => \N__13690\,
            I => \N__13681\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__13687\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__13684\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__13681\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13670\
        );

    \I__2286\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13667\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__13670\,
            I => \transmit_module.video_signal_controller.n3379\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__13667\,
            I => \transmit_module.video_signal_controller.n3379\
        );

    \I__2283\ : InMux
    port map (
            O => \N__13662\,
            I => \receive_module.rx_counter.n3207\
        );

    \I__2282\ : InMux
    port map (
            O => \N__13659\,
            I => \receive_module.rx_counter.n3208\
        );

    \I__2281\ : InMux
    port map (
            O => \N__13656\,
            I => \receive_module.rx_counter.n3209\
        );

    \I__2280\ : InMux
    port map (
            O => \N__13653\,
            I => \receive_module.rx_counter.n3210\
        );

    \I__2279\ : InMux
    port map (
            O => \N__13650\,
            I => \receive_module.rx_counter.n3211\
        );

    \I__2278\ : InMux
    port map (
            O => \N__13647\,
            I => \receive_module.rx_counter.n3212\
        );

    \I__2277\ : InMux
    port map (
            O => \N__13644\,
            I => \receive_module.rx_counter.n3213\
        );

    \I__2276\ : InMux
    port map (
            O => \N__13641\,
            I => \bfn_15_11_0_\
        );

    \I__2275\ : InMux
    port map (
            O => \N__13638\,
            I => \receive_module.rx_counter.n3215\
        );

    \I__2274\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13632\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__13632\,
            I => \N__13629\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__13629\,
            I => \N__13626\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__13626\,
            I => \TVP_VIDEO_c_5\
        );

    \I__2270\ : IoInMux
    port map (
            O => \N__13623\,
            I => \N__13620\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__13620\,
            I => \N__13617\
        );

    \I__2268\ : IoSpan4Mux
    port map (
            O => \N__13617\,
            I => \N__13614\
        );

    \I__2267\ : Span4Mux_s1_h
    port map (
            O => \N__13614\,
            I => \N__13611\
        );

    \I__2266\ : Sp12to4
    port map (
            O => \N__13611\,
            I => \N__13607\
        );

    \I__2265\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13604\
        );

    \I__2264\ : Span12Mux_h
    port map (
            O => \N__13607\,
            I => \N__13601\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__13604\,
            I => \N__13598\
        );

    \I__2262\ : Odrv12
    port map (
            O => \N__13601\,
            I => \DEBUG_c_1_c\
        );

    \I__2261\ : Odrv12
    port map (
            O => \N__13598\,
            I => \DEBUG_c_1_c\
        );

    \I__2260\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13590\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__13590\,
            I => \tvp_vs_buffer.BUFFER_0_0\
        );

    \I__2258\ : InMux
    port map (
            O => \N__13587\,
            I => \N__13584\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__13584\,
            I => \tvp_vs_buffer.BUFFER_1_0\
        );

    \I__2256\ : InMux
    port map (
            O => \N__13581\,
            I => \N__13577\
        );

    \I__2255\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13574\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__13577\,
            I => \N__13567\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__13574\,
            I => \N__13564\
        );

    \I__2252\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13561\
        );

    \I__2251\ : InMux
    port map (
            O => \N__13572\,
            I => \N__13558\
        );

    \I__2250\ : InMux
    port map (
            O => \N__13571\,
            I => \N__13555\
        );

    \I__2249\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13550\
        );

    \I__2248\ : Span12Mux_s8_h
    port map (
            O => \N__13567\,
            I => \N__13546\
        );

    \I__2247\ : Span12Mux_s7_v
    port map (
            O => \N__13564\,
            I => \N__13541\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__13561\,
            I => \N__13541\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__13558\,
            I => \N__13536\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__13555\,
            I => \N__13536\
        );

    \I__2243\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13533\
        );

    \I__2242\ : InMux
    port map (
            O => \N__13553\,
            I => \N__13530\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__13550\,
            I => \N__13527\
        );

    \I__2240\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13524\
        );

    \I__2239\ : Span12Mux_v
    port map (
            O => \N__13546\,
            I => \N__13521\
        );

    \I__2238\ : Span12Mux_v
    port map (
            O => \N__13541\,
            I => \N__13518\
        );

    \I__2237\ : Span12Mux_v
    port map (
            O => \N__13536\,
            I => \N__13515\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__13533\,
            I => \N__13512\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__13530\,
            I => \N__13509\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__13527\,
            I => \N__13506\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__13524\,
            I => \N__13503\
        );

    \I__2232\ : Span12Mux_v
    port map (
            O => \N__13521\,
            I => \N__13500\
        );

    \I__2231\ : Span12Mux_h
    port map (
            O => \N__13518\,
            I => \N__13491\
        );

    \I__2230\ : Span12Mux_h
    port map (
            O => \N__13515\,
            I => \N__13491\
        );

    \I__2229\ : Span12Mux_h
    port map (
            O => \N__13512\,
            I => \N__13491\
        );

    \I__2228\ : Span12Mux_h
    port map (
            O => \N__13509\,
            I => \N__13491\
        );

    \I__2227\ : Span4Mux_h
    port map (
            O => \N__13506\,
            I => \N__13488\
        );

    \I__2226\ : Span4Mux_v
    port map (
            O => \N__13503\,
            I => \N__13485\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__13500\,
            I => \RX_DATA_5\
        );

    \I__2224\ : Odrv12
    port map (
            O => \N__13491\,
            I => \RX_DATA_5\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__13488\,
            I => \RX_DATA_5\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__13485\,
            I => \RX_DATA_5\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__13476\,
            I => \receive_module.sync_wd.n6_cascade_\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__13473\,
            I => \receive_module.sync_wd.n4_cascade_\
        );

    \I__2219\ : InMux
    port map (
            O => \N__13470\,
            I => \N__13467\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__13467\,
            I => \receive_module.sync_wd.old_visible\
        );

    \I__2217\ : InMux
    port map (
            O => \N__13464\,
            I => \bfn_15_10_0_\
        );

    \I__2216\ : CascadeMux
    port map (
            O => \N__13461\,
            I => \N__13457\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__13460\,
            I => \N__13454\
        );

    \I__2214\ : CascadeBuf
    port map (
            O => \N__13457\,
            I => \N__13451\
        );

    \I__2213\ : CascadeBuf
    port map (
            O => \N__13454\,
            I => \N__13448\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__13451\,
            I => \N__13445\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__13448\,
            I => \N__13442\
        );

    \I__2210\ : CascadeBuf
    port map (
            O => \N__13445\,
            I => \N__13439\
        );

    \I__2209\ : CascadeBuf
    port map (
            O => \N__13442\,
            I => \N__13436\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__13439\,
            I => \N__13433\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__13436\,
            I => \N__13430\
        );

    \I__2206\ : CascadeBuf
    port map (
            O => \N__13433\,
            I => \N__13427\
        );

    \I__2205\ : CascadeBuf
    port map (
            O => \N__13430\,
            I => \N__13424\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__13427\,
            I => \N__13421\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__13424\,
            I => \N__13418\
        );

    \I__2202\ : CascadeBuf
    port map (
            O => \N__13421\,
            I => \N__13415\
        );

    \I__2201\ : CascadeBuf
    port map (
            O => \N__13418\,
            I => \N__13412\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__13415\,
            I => \N__13409\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__13412\,
            I => \N__13406\
        );

    \I__2198\ : CascadeBuf
    port map (
            O => \N__13409\,
            I => \N__13403\
        );

    \I__2197\ : CascadeBuf
    port map (
            O => \N__13406\,
            I => \N__13400\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__13403\,
            I => \N__13397\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__13400\,
            I => \N__13394\
        );

    \I__2194\ : CascadeBuf
    port map (
            O => \N__13397\,
            I => \N__13391\
        );

    \I__2193\ : CascadeBuf
    port map (
            O => \N__13394\,
            I => \N__13388\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__13391\,
            I => \N__13385\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__13388\,
            I => \N__13382\
        );

    \I__2190\ : CascadeBuf
    port map (
            O => \N__13385\,
            I => \N__13379\
        );

    \I__2189\ : CascadeBuf
    port map (
            O => \N__13382\,
            I => \N__13376\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__13379\,
            I => \N__13373\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__13376\,
            I => \N__13370\
        );

    \I__2186\ : CascadeBuf
    port map (
            O => \N__13373\,
            I => \N__13367\
        );

    \I__2185\ : CascadeBuf
    port map (
            O => \N__13370\,
            I => \N__13364\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__13367\,
            I => \N__13361\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__13364\,
            I => \N__13358\
        );

    \I__2182\ : CascadeBuf
    port map (
            O => \N__13361\,
            I => \N__13355\
        );

    \I__2181\ : CascadeBuf
    port map (
            O => \N__13358\,
            I => \N__13352\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__13355\,
            I => \N__13349\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__13352\,
            I => \N__13346\
        );

    \I__2178\ : CascadeBuf
    port map (
            O => \N__13349\,
            I => \N__13343\
        );

    \I__2177\ : CascadeBuf
    port map (
            O => \N__13346\,
            I => \N__13340\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__13343\,
            I => \N__13337\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__13340\,
            I => \N__13334\
        );

    \I__2174\ : CascadeBuf
    port map (
            O => \N__13337\,
            I => \N__13331\
        );

    \I__2173\ : CascadeBuf
    port map (
            O => \N__13334\,
            I => \N__13328\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__13331\,
            I => \N__13325\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__13328\,
            I => \N__13322\
        );

    \I__2170\ : CascadeBuf
    port map (
            O => \N__13325\,
            I => \N__13319\
        );

    \I__2169\ : CascadeBuf
    port map (
            O => \N__13322\,
            I => \N__13316\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__13319\,
            I => \N__13313\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__13316\,
            I => \N__13310\
        );

    \I__2166\ : CascadeBuf
    port map (
            O => \N__13313\,
            I => \N__13307\
        );

    \I__2165\ : CascadeBuf
    port map (
            O => \N__13310\,
            I => \N__13304\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__13307\,
            I => \N__13301\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__13304\,
            I => \N__13298\
        );

    \I__2162\ : CascadeBuf
    port map (
            O => \N__13301\,
            I => \N__13295\
        );

    \I__2161\ : CascadeBuf
    port map (
            O => \N__13298\,
            I => \N__13292\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__13295\,
            I => \N__13289\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__13292\,
            I => \N__13286\
        );

    \I__2158\ : CascadeBuf
    port map (
            O => \N__13289\,
            I => \N__13283\
        );

    \I__2157\ : CascadeBuf
    port map (
            O => \N__13286\,
            I => \N__13280\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__13283\,
            I => \N__13277\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__13280\,
            I => \N__13274\
        );

    \I__2154\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13271\
        );

    \I__2153\ : InMux
    port map (
            O => \N__13274\,
            I => \N__13268\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__13271\,
            I => \N__13265\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__13268\,
            I => \N__13262\
        );

    \I__2150\ : Sp12to4
    port map (
            O => \N__13265\,
            I => \N__13259\
        );

    \I__2149\ : Span12Mux_s9_h
    port map (
            O => \N__13262\,
            I => \N__13256\
        );

    \I__2148\ : Span12Mux_s5_v
    port map (
            O => \N__13259\,
            I => \N__13253\
        );

    \I__2147\ : Span12Mux_v
    port map (
            O => \N__13256\,
            I => \N__13250\
        );

    \I__2146\ : Span12Mux_h
    port map (
            O => \N__13253\,
            I => \N__13247\
        );

    \I__2145\ : Odrv12
    port map (
            O => \N__13250\,
            I => n22
        );

    \I__2144\ : Odrv12
    port map (
            O => \N__13247\,
            I => n22
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__13242\,
            I => \transmit_module.n112_cascade_\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__13239\,
            I => \N__13236\
        );

    \I__2141\ : CascadeBuf
    port map (
            O => \N__13236\,
            I => \N__13232\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__13235\,
            I => \N__13229\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__13232\,
            I => \N__13226\
        );

    \I__2138\ : CascadeBuf
    port map (
            O => \N__13229\,
            I => \N__13223\
        );

    \I__2137\ : CascadeBuf
    port map (
            O => \N__13226\,
            I => \N__13220\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__13223\,
            I => \N__13217\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__13220\,
            I => \N__13214\
        );

    \I__2134\ : CascadeBuf
    port map (
            O => \N__13217\,
            I => \N__13211\
        );

    \I__2133\ : CascadeBuf
    port map (
            O => \N__13214\,
            I => \N__13208\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__13211\,
            I => \N__13205\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__13208\,
            I => \N__13202\
        );

    \I__2130\ : CascadeBuf
    port map (
            O => \N__13205\,
            I => \N__13199\
        );

    \I__2129\ : CascadeBuf
    port map (
            O => \N__13202\,
            I => \N__13196\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__13199\,
            I => \N__13193\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__13196\,
            I => \N__13190\
        );

    \I__2126\ : CascadeBuf
    port map (
            O => \N__13193\,
            I => \N__13187\
        );

    \I__2125\ : CascadeBuf
    port map (
            O => \N__13190\,
            I => \N__13184\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__13187\,
            I => \N__13181\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__13184\,
            I => \N__13178\
        );

    \I__2122\ : CascadeBuf
    port map (
            O => \N__13181\,
            I => \N__13175\
        );

    \I__2121\ : CascadeBuf
    port map (
            O => \N__13178\,
            I => \N__13172\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__13175\,
            I => \N__13169\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__13172\,
            I => \N__13166\
        );

    \I__2118\ : CascadeBuf
    port map (
            O => \N__13169\,
            I => \N__13163\
        );

    \I__2117\ : CascadeBuf
    port map (
            O => \N__13166\,
            I => \N__13160\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__13163\,
            I => \N__13157\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__13160\,
            I => \N__13154\
        );

    \I__2114\ : CascadeBuf
    port map (
            O => \N__13157\,
            I => \N__13151\
        );

    \I__2113\ : CascadeBuf
    port map (
            O => \N__13154\,
            I => \N__13148\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__13151\,
            I => \N__13145\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__13148\,
            I => \N__13142\
        );

    \I__2110\ : CascadeBuf
    port map (
            O => \N__13145\,
            I => \N__13139\
        );

    \I__2109\ : CascadeBuf
    port map (
            O => \N__13142\,
            I => \N__13136\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__13139\,
            I => \N__13133\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__13136\,
            I => \N__13130\
        );

    \I__2106\ : CascadeBuf
    port map (
            O => \N__13133\,
            I => \N__13127\
        );

    \I__2105\ : CascadeBuf
    port map (
            O => \N__13130\,
            I => \N__13124\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__13127\,
            I => \N__13121\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__13124\,
            I => \N__13118\
        );

    \I__2102\ : CascadeBuf
    port map (
            O => \N__13121\,
            I => \N__13115\
        );

    \I__2101\ : CascadeBuf
    port map (
            O => \N__13118\,
            I => \N__13112\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__13115\,
            I => \N__13109\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__13112\,
            I => \N__13106\
        );

    \I__2098\ : CascadeBuf
    port map (
            O => \N__13109\,
            I => \N__13103\
        );

    \I__2097\ : CascadeBuf
    port map (
            O => \N__13106\,
            I => \N__13100\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__13103\,
            I => \N__13097\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__13100\,
            I => \N__13094\
        );

    \I__2094\ : CascadeBuf
    port map (
            O => \N__13097\,
            I => \N__13091\
        );

    \I__2093\ : CascadeBuf
    port map (
            O => \N__13094\,
            I => \N__13088\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__13091\,
            I => \N__13085\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__13088\,
            I => \N__13082\
        );

    \I__2090\ : CascadeBuf
    port map (
            O => \N__13085\,
            I => \N__13079\
        );

    \I__2089\ : CascadeBuf
    port map (
            O => \N__13082\,
            I => \N__13076\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__13079\,
            I => \N__13073\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__13076\,
            I => \N__13070\
        );

    \I__2086\ : CascadeBuf
    port map (
            O => \N__13073\,
            I => \N__13067\
        );

    \I__2085\ : CascadeBuf
    port map (
            O => \N__13070\,
            I => \N__13064\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__13067\,
            I => \N__13061\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__13064\,
            I => \N__13058\
        );

    \I__2082\ : CascadeBuf
    port map (
            O => \N__13061\,
            I => \N__13055\
        );

    \I__2081\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13052\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__13055\,
            I => \N__13049\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__13052\,
            I => \N__13046\
        );

    \I__2078\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13043\
        );

    \I__2077\ : Span12Mux_h
    port map (
            O => \N__13046\,
            I => \N__13040\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__13043\,
            I => \N__13037\
        );

    \I__2075\ : Span12Mux_v
    port map (
            O => \N__13040\,
            I => \N__13032\
        );

    \I__2074\ : Span12Mux_v
    port map (
            O => \N__13037\,
            I => \N__13032\
        );

    \I__2073\ : Odrv12
    port map (
            O => \N__13032\,
            I => n24
        );

    \I__2072\ : InMux
    port map (
            O => \N__13029\,
            I => \N__13026\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__13026\,
            I => \N__13023\
        );

    \I__2070\ : Odrv12
    port map (
            O => \N__13023\,
            I => \transmit_module.n125\
        );

    \I__2069\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13017\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__13017\,
            I => \N__13014\
        );

    \I__2067\ : Span4Mux_h
    port map (
            O => \N__13014\,
            I => \N__13011\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__13011\,
            I => \transmit_module.n140\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__13008\,
            I => \transmit_module.n140_cascade_\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__13005\,
            I => \N__13002\
        );

    \I__2063\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12999\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12999\,
            I => \N__12996\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__12996\,
            I => \N__12992\
        );

    \I__2060\ : InMux
    port map (
            O => \N__12995\,
            I => \N__12989\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__12992\,
            I => \transmit_module.n109\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__12989\,
            I => \transmit_module.n109\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__12984\,
            I => \N__12981\
        );

    \I__2056\ : CascadeBuf
    port map (
            O => \N__12981\,
            I => \N__12977\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__12980\,
            I => \N__12974\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__12977\,
            I => \N__12971\
        );

    \I__2053\ : CascadeBuf
    port map (
            O => \N__12974\,
            I => \N__12968\
        );

    \I__2052\ : CascadeBuf
    port map (
            O => \N__12971\,
            I => \N__12965\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__12968\,
            I => \N__12962\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__12965\,
            I => \N__12959\
        );

    \I__2049\ : CascadeBuf
    port map (
            O => \N__12962\,
            I => \N__12956\
        );

    \I__2048\ : CascadeBuf
    port map (
            O => \N__12959\,
            I => \N__12953\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__12956\,
            I => \N__12950\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__12953\,
            I => \N__12947\
        );

    \I__2045\ : CascadeBuf
    port map (
            O => \N__12950\,
            I => \N__12944\
        );

    \I__2044\ : CascadeBuf
    port map (
            O => \N__12947\,
            I => \N__12941\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__12944\,
            I => \N__12938\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__12941\,
            I => \N__12935\
        );

    \I__2041\ : CascadeBuf
    port map (
            O => \N__12938\,
            I => \N__12932\
        );

    \I__2040\ : CascadeBuf
    port map (
            O => \N__12935\,
            I => \N__12929\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__12932\,
            I => \N__12926\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__12929\,
            I => \N__12923\
        );

    \I__2037\ : CascadeBuf
    port map (
            O => \N__12926\,
            I => \N__12920\
        );

    \I__2036\ : CascadeBuf
    port map (
            O => \N__12923\,
            I => \N__12917\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__12920\,
            I => \N__12914\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__12917\,
            I => \N__12911\
        );

    \I__2033\ : CascadeBuf
    port map (
            O => \N__12914\,
            I => \N__12908\
        );

    \I__2032\ : CascadeBuf
    port map (
            O => \N__12911\,
            I => \N__12905\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__12908\,
            I => \N__12902\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__12905\,
            I => \N__12899\
        );

    \I__2029\ : CascadeBuf
    port map (
            O => \N__12902\,
            I => \N__12896\
        );

    \I__2028\ : CascadeBuf
    port map (
            O => \N__12899\,
            I => \N__12893\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__12896\,
            I => \N__12890\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__12893\,
            I => \N__12887\
        );

    \I__2025\ : CascadeBuf
    port map (
            O => \N__12890\,
            I => \N__12884\
        );

    \I__2024\ : CascadeBuf
    port map (
            O => \N__12887\,
            I => \N__12881\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__12884\,
            I => \N__12878\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__12881\,
            I => \N__12875\
        );

    \I__2021\ : CascadeBuf
    port map (
            O => \N__12878\,
            I => \N__12872\
        );

    \I__2020\ : CascadeBuf
    port map (
            O => \N__12875\,
            I => \N__12869\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__12872\,
            I => \N__12866\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__12869\,
            I => \N__12863\
        );

    \I__2017\ : CascadeBuf
    port map (
            O => \N__12866\,
            I => \N__12860\
        );

    \I__2016\ : CascadeBuf
    port map (
            O => \N__12863\,
            I => \N__12857\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__12860\,
            I => \N__12854\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__12857\,
            I => \N__12851\
        );

    \I__2013\ : CascadeBuf
    port map (
            O => \N__12854\,
            I => \N__12848\
        );

    \I__2012\ : CascadeBuf
    port map (
            O => \N__12851\,
            I => \N__12845\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__12848\,
            I => \N__12842\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__12845\,
            I => \N__12839\
        );

    \I__2009\ : CascadeBuf
    port map (
            O => \N__12842\,
            I => \N__12836\
        );

    \I__2008\ : CascadeBuf
    port map (
            O => \N__12839\,
            I => \N__12833\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__12836\,
            I => \N__12830\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__12833\,
            I => \N__12827\
        );

    \I__2005\ : CascadeBuf
    port map (
            O => \N__12830\,
            I => \N__12824\
        );

    \I__2004\ : CascadeBuf
    port map (
            O => \N__12827\,
            I => \N__12821\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__12824\,
            I => \N__12818\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__12821\,
            I => \N__12815\
        );

    \I__2001\ : CascadeBuf
    port map (
            O => \N__12818\,
            I => \N__12812\
        );

    \I__2000\ : CascadeBuf
    port map (
            O => \N__12815\,
            I => \N__12809\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__12812\,
            I => \N__12806\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__12809\,
            I => \N__12803\
        );

    \I__1997\ : CascadeBuf
    port map (
            O => \N__12806\,
            I => \N__12800\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12797\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__12800\,
            I => \N__12794\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__12797\,
            I => \N__12791\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12788\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__12791\,
            I => \N__12785\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__12788\,
            I => \N__12782\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__12785\,
            I => \N__12779\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__12782\,
            I => \N__12776\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__12779\,
            I => \N__12773\
        );

    \I__1987\ : Span4Mux_v
    port map (
            O => \N__12776\,
            I => \N__12770\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__12773\,
            I => \N__12767\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__12770\,
            I => \N__12764\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__12767\,
            I => \N__12759\
        );

    \I__1983\ : Span4Mux_h
    port map (
            O => \N__12764\,
            I => \N__12759\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__12759\,
            I => n21
        );

    \I__1981\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12752\
        );

    \I__1980\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12749\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__12752\,
            I => \transmit_module.n106\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__12749\,
            I => \transmit_module.n106\
        );

    \I__1977\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12740\
        );

    \I__1976\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12737\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__12740\,
            I => \transmit_module.n137\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__12737\,
            I => \transmit_module.n137\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__1972\ : CascadeBuf
    port map (
            O => \N__12729\,
            I => \N__12725\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__12728\,
            I => \N__12722\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__12725\,
            I => \N__12719\
        );

    \I__1969\ : CascadeBuf
    port map (
            O => \N__12722\,
            I => \N__12716\
        );

    \I__1968\ : CascadeBuf
    port map (
            O => \N__12719\,
            I => \N__12713\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__12716\,
            I => \N__12710\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__12713\,
            I => \N__12707\
        );

    \I__1965\ : CascadeBuf
    port map (
            O => \N__12710\,
            I => \N__12704\
        );

    \I__1964\ : CascadeBuf
    port map (
            O => \N__12707\,
            I => \N__12701\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__12704\,
            I => \N__12698\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__12701\,
            I => \N__12695\
        );

    \I__1961\ : CascadeBuf
    port map (
            O => \N__12698\,
            I => \N__12692\
        );

    \I__1960\ : CascadeBuf
    port map (
            O => \N__12695\,
            I => \N__12689\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__12692\,
            I => \N__12686\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__12689\,
            I => \N__12683\
        );

    \I__1957\ : CascadeBuf
    port map (
            O => \N__12686\,
            I => \N__12680\
        );

    \I__1956\ : CascadeBuf
    port map (
            O => \N__12683\,
            I => \N__12677\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__12680\,
            I => \N__12674\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__12677\,
            I => \N__12671\
        );

    \I__1953\ : CascadeBuf
    port map (
            O => \N__12674\,
            I => \N__12668\
        );

    \I__1952\ : CascadeBuf
    port map (
            O => \N__12671\,
            I => \N__12665\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__12668\,
            I => \N__12662\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__12665\,
            I => \N__12659\
        );

    \I__1949\ : CascadeBuf
    port map (
            O => \N__12662\,
            I => \N__12656\
        );

    \I__1948\ : CascadeBuf
    port map (
            O => \N__12659\,
            I => \N__12653\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__12656\,
            I => \N__12650\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__12653\,
            I => \N__12647\
        );

    \I__1945\ : CascadeBuf
    port map (
            O => \N__12650\,
            I => \N__12644\
        );

    \I__1944\ : CascadeBuf
    port map (
            O => \N__12647\,
            I => \N__12641\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__12644\,
            I => \N__12638\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__12641\,
            I => \N__12635\
        );

    \I__1941\ : CascadeBuf
    port map (
            O => \N__12638\,
            I => \N__12632\
        );

    \I__1940\ : CascadeBuf
    port map (
            O => \N__12635\,
            I => \N__12629\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__12632\,
            I => \N__12626\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__12629\,
            I => \N__12623\
        );

    \I__1937\ : CascadeBuf
    port map (
            O => \N__12626\,
            I => \N__12620\
        );

    \I__1936\ : CascadeBuf
    port map (
            O => \N__12623\,
            I => \N__12617\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__12620\,
            I => \N__12614\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__12617\,
            I => \N__12611\
        );

    \I__1933\ : CascadeBuf
    port map (
            O => \N__12614\,
            I => \N__12608\
        );

    \I__1932\ : CascadeBuf
    port map (
            O => \N__12611\,
            I => \N__12605\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__12608\,
            I => \N__12602\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__12605\,
            I => \N__12599\
        );

    \I__1929\ : CascadeBuf
    port map (
            O => \N__12602\,
            I => \N__12596\
        );

    \I__1928\ : CascadeBuf
    port map (
            O => \N__12599\,
            I => \N__12593\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__12596\,
            I => \N__12590\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__12593\,
            I => \N__12587\
        );

    \I__1925\ : CascadeBuf
    port map (
            O => \N__12590\,
            I => \N__12584\
        );

    \I__1924\ : CascadeBuf
    port map (
            O => \N__12587\,
            I => \N__12581\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__12584\,
            I => \N__12578\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__12581\,
            I => \N__12575\
        );

    \I__1921\ : CascadeBuf
    port map (
            O => \N__12578\,
            I => \N__12572\
        );

    \I__1920\ : CascadeBuf
    port map (
            O => \N__12575\,
            I => \N__12569\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__12572\,
            I => \N__12566\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__12569\,
            I => \N__12563\
        );

    \I__1917\ : CascadeBuf
    port map (
            O => \N__12566\,
            I => \N__12560\
        );

    \I__1916\ : CascadeBuf
    port map (
            O => \N__12563\,
            I => \N__12557\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__12560\,
            I => \N__12554\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__12557\,
            I => \N__12551\
        );

    \I__1913\ : CascadeBuf
    port map (
            O => \N__12554\,
            I => \N__12548\
        );

    \I__1912\ : InMux
    port map (
            O => \N__12551\,
            I => \N__12545\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__12548\,
            I => \N__12542\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__12545\,
            I => \N__12539\
        );

    \I__1909\ : InMux
    port map (
            O => \N__12542\,
            I => \N__12536\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__12539\,
            I => \N__12533\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__12536\,
            I => \N__12530\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__12533\,
            I => \N__12527\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__12530\,
            I => \N__12524\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__12527\,
            I => \N__12521\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__12524\,
            I => \N__12518\
        );

    \I__1902\ : Span4Mux_h
    port map (
            O => \N__12521\,
            I => \N__12515\
        );

    \I__1901\ : Span4Mux_v
    port map (
            O => \N__12518\,
            I => \N__12512\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__12515\,
            I => \N__12507\
        );

    \I__1899\ : Span4Mux_h
    port map (
            O => \N__12512\,
            I => \N__12507\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__12507\,
            I => n18
        );

    \I__1897\ : InMux
    port map (
            O => \N__12504\,
            I => \transmit_module.n3171\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__12501\,
            I => \N__12495\
        );

    \I__1895\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12492\
        );

    \I__1894\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12489\
        );

    \I__1893\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12484\
        );

    \I__1892\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12484\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__12492\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__12489\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__12484\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__1888\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12474\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__12474\,
            I => \transmit_module.ADDR_Y_COMPONENT_9\
        );

    \I__1886\ : InMux
    port map (
            O => \N__12471\,
            I => \N__12468\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__12468\,
            I => \N__12465\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__12465\,
            I => \transmit_module.ADDR_Y_COMPONENT_0\
        );

    \I__1883\ : InMux
    port map (
            O => \N__12462\,
            I => \N__12457\
        );

    \I__1882\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12454\
        );

    \I__1881\ : InMux
    port map (
            O => \N__12460\,
            I => \N__12450\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__12457\,
            I => \N__12445\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__12454\,
            I => \N__12445\
        );

    \I__1878\ : InMux
    port map (
            O => \N__12453\,
            I => \N__12442\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__12450\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__12445\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__12442\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__1874\ : InMux
    port map (
            O => \N__12435\,
            I => \N__12432\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__12432\,
            I => \transmit_module.ADDR_Y_COMPONENT_1\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__12429\,
            I => \N__12423\
        );

    \I__1871\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12420\
        );

    \I__1870\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12415\
        );

    \I__1869\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12415\
        );

    \I__1868\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12412\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__12420\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__12415\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__12412\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__1864\ : InMux
    port map (
            O => \N__12405\,
            I => \N__12402\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__12402\,
            I => \transmit_module.ADDR_Y_COMPONENT_8\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__12399\,
            I => \N__12393\
        );

    \I__1861\ : InMux
    port map (
            O => \N__12398\,
            I => \N__12390\
        );

    \I__1860\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12385\
        );

    \I__1859\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12385\
        );

    \I__1858\ : InMux
    port map (
            O => \N__12393\,
            I => \N__12382\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__12390\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__12385\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__12382\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__1854\ : InMux
    port map (
            O => \N__12375\,
            I => \N__12372\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__12372\,
            I => \transmit_module.ADDR_Y_COMPONENT_5\
        );

    \I__1852\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12366\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__12366\,
            I => \N__12363\
        );

    \I__1850\ : Span4Mux_h
    port map (
            O => \N__12363\,
            I => \N__12357\
        );

    \I__1849\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12354\
        );

    \I__1848\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12351\
        );

    \I__1847\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12348\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__12357\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__12354\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__12351\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__12348\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__1842\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12336\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__12336\,
            I => \N__12333\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__12333\,
            I => \transmit_module.n122\
        );

    \I__1839\ : InMux
    port map (
            O => \N__12330\,
            I => \transmit_module.n3162\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__12327\,
            I => \N__12324\
        );

    \I__1837\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12321\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__12321\,
            I => \N__12318\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__12318\,
            I => \transmit_module.n127\
        );

    \I__1834\ : InMux
    port map (
            O => \N__12315\,
            I => \transmit_module.n3163\
        );

    \I__1833\ : InMux
    port map (
            O => \N__12312\,
            I => \transmit_module.n3164\
        );

    \I__1832\ : InMux
    port map (
            O => \N__12309\,
            I => \transmit_module.n3165\
        );

    \I__1831\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12303\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12300\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__12300\,
            I => \transmit_module.n124\
        );

    \I__1828\ : InMux
    port map (
            O => \N__12297\,
            I => \bfn_14_16_0_\
        );

    \I__1827\ : InMux
    port map (
            O => \N__12294\,
            I => \N__12291\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__12291\,
            I => \transmit_module.n123\
        );

    \I__1825\ : InMux
    port map (
            O => \N__12288\,
            I => \transmit_module.n3167\
        );

    \I__1824\ : InMux
    port map (
            O => \N__12285\,
            I => \transmit_module.n3168\
        );

    \I__1823\ : InMux
    port map (
            O => \N__12282\,
            I => \transmit_module.n3169\
        );

    \I__1822\ : InMux
    port map (
            O => \N__12279\,
            I => \transmit_module.n3170\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__12276\,
            I => \transmit_module.video_signal_controller.n6_adj_623_cascade_\
        );

    \I__1820\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12269\
        );

    \I__1819\ : InMux
    port map (
            O => \N__12272\,
            I => \N__12266\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__12269\,
            I => \N__12263\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__12266\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_588\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__12263\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_588\
        );

    \I__1815\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12252\
        );

    \I__1814\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12249\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__12256\,
            I => \N__12246\
        );

    \I__1812\ : InMux
    port map (
            O => \N__12255\,
            I => \N__12243\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__12252\,
            I => \N__12237\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__12249\,
            I => \N__12237\
        );

    \I__1809\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12234\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__12243\,
            I => \N__12231\
        );

    \I__1807\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12228\
        );

    \I__1806\ : Span4Mux_h
    port map (
            O => \N__12237\,
            I => \N__12225\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__12234\,
            I => \N__12220\
        );

    \I__1804\ : Span4Mux_h
    port map (
            O => \N__12231\,
            I => \N__12220\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__12228\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__12225\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__12220\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__12213\,
            I => \transmit_module.video_signal_controller.n7_adj_624_cascade_\
        );

    \I__1799\ : InMux
    port map (
            O => \N__12210\,
            I => \N__12204\
        );

    \I__1798\ : InMux
    port map (
            O => \N__12209\,
            I => \N__12204\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__12204\,
            I => \transmit_module.video_signal_controller.n3004\
        );

    \I__1796\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12194\
        );

    \I__1795\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12194\
        );

    \I__1794\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12190\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__12194\,
            I => \N__12186\
        );

    \I__1792\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12183\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__12190\,
            I => \N__12180\
        );

    \I__1790\ : InMux
    port map (
            O => \N__12189\,
            I => \N__12177\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__12186\,
            I => \N__12174\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__12183\,
            I => \N__12169\
        );

    \I__1787\ : Span4Mux_h
    port map (
            O => \N__12180\,
            I => \N__12169\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__12177\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__12174\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__12169\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1783\ : InMux
    port map (
            O => \N__12162\,
            I => \N__12156\
        );

    \I__1782\ : InMux
    port map (
            O => \N__12161\,
            I => \N__12151\
        );

    \I__1781\ : InMux
    port map (
            O => \N__12160\,
            I => \N__12151\
        );

    \I__1780\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12147\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__12156\,
            I => \N__12144\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__12151\,
            I => \N__12141\
        );

    \I__1777\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12138\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__12147\,
            I => \N__12133\
        );

    \I__1775\ : Span4Mux_h
    port map (
            O => \N__12144\,
            I => \N__12133\
        );

    \I__1774\ : Span4Mux_h
    port map (
            O => \N__12141\,
            I => \N__12130\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__12138\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__12133\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__12130\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1770\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12120\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__12120\,
            I => \transmit_module.video_signal_controller.n3014\
        );

    \I__1768\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12114\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__12114\,
            I => \transmit_module.n131\
        );

    \I__1766\ : InMux
    port map (
            O => \N__12111\,
            I => \transmit_module.n3159\
        );

    \I__1765\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12101\
        );

    \I__1764\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12101\
        );

    \I__1763\ : InMux
    port map (
            O => \N__12106\,
            I => \N__12097\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__12101\,
            I => \N__12094\
        );

    \I__1761\ : InMux
    port map (
            O => \N__12100\,
            I => \N__12091\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__12097\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__12094\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__12091\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__1757\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12081\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__12081\,
            I => \transmit_module.n130\
        );

    \I__1755\ : InMux
    port map (
            O => \N__12078\,
            I => \transmit_module.n3160\
        );

    \I__1754\ : InMux
    port map (
            O => \N__12075\,
            I => \N__12070\
        );

    \I__1753\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12065\
        );

    \I__1752\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12065\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__12070\,
            I => \N__12061\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__12065\,
            I => \N__12058\
        );

    \I__1749\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12055\
        );

    \I__1748\ : Odrv12
    port map (
            O => \N__12061\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__12058\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__12055\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__1745\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12045\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__12045\,
            I => \N__12042\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__12042\,
            I => \N__12039\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__12039\,
            I => \transmit_module.n129\
        );

    \I__1741\ : InMux
    port map (
            O => \N__12036\,
            I => \transmit_module.n3161\
        );

    \I__1740\ : InMux
    port map (
            O => \N__12033\,
            I => \N__12030\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__12030\,
            I => \N__12027\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__12027\,
            I => \N__12021\
        );

    \I__1737\ : InMux
    port map (
            O => \N__12026\,
            I => \N__12018\
        );

    \I__1736\ : InMux
    port map (
            O => \N__12025\,
            I => \N__12013\
        );

    \I__1735\ : InMux
    port map (
            O => \N__12024\,
            I => \N__12013\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__12021\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__12018\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__12013\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1731\ : InMux
    port map (
            O => \N__12006\,
            I => \N__12003\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__12003\,
            I => \transmit_module.video_signal_controller.n3517\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__12000\,
            I => \N__11997\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11997\,
            I => \N__11994\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__11994\,
            I => \N__11988\
        );

    \I__1726\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11985\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11980\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11991\,
            I => \N__11980\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__11988\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11985\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__11980\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11973\,
            I => \N__11969\
        );

    \I__1719\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11966\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__11969\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__11966\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1716\ : InMux
    port map (
            O => \N__11961\,
            I => \N__11958\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__11958\,
            I => \transmit_module.video_signal_controller.n2955\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11950\
        );

    \I__1713\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11944\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11944\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__11950\,
            I => \N__11941\
        );

    \I__1710\ : InMux
    port map (
            O => \N__11949\,
            I => \N__11938\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__11944\,
            I => \N__11933\
        );

    \I__1708\ : Span4Mux_h
    port map (
            O => \N__11941\,
            I => \N__11933\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__11938\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__11933\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__11928\,
            I => \N__11924\
        );

    \I__1704\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11921\
        );

    \I__1703\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11918\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11921\,
            I => \transmit_module.video_signal_controller.n3363\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__11918\,
            I => \transmit_module.video_signal_controller.n3363\
        );

    \I__1700\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11910\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__11910\,
            I => \transmit_module.video_signal_controller.n2014\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__11907\,
            I => \transmit_module.video_signal_controller.n2972_cascade_\
        );

    \I__1697\ : SRMux
    port map (
            O => \N__11904\,
            I => \N__11901\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__11901\,
            I => \N__11895\
        );

    \I__1695\ : SRMux
    port map (
            O => \N__11900\,
            I => \N__11892\
        );

    \I__1694\ : CEMux
    port map (
            O => \N__11899\,
            I => \N__11888\
        );

    \I__1693\ : CEMux
    port map (
            O => \N__11898\,
            I => \N__11885\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__11895\,
            I => \N__11882\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__11892\,
            I => \N__11879\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11876\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__11888\,
            I => \N__11873\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__11885\,
            I => \N__11864\
        );

    \I__1687\ : Span4Mux_v
    port map (
            O => \N__11882\,
            I => \N__11864\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__11879\,
            I => \N__11864\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__11876\,
            I => \N__11864\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__11873\,
            I => \transmit_module.video_signal_controller.n2047\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__11864\,
            I => \transmit_module.video_signal_controller.n2047\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__11859\,
            I => \N__11854\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__11858\,
            I => \N__11851\
        );

    \I__1680\ : InMux
    port map (
            O => \N__11857\,
            I => \N__11847\
        );

    \I__1679\ : InMux
    port map (
            O => \N__11854\,
            I => \N__11842\
        );

    \I__1678\ : InMux
    port map (
            O => \N__11851\,
            I => \N__11842\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11850\,
            I => \N__11839\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__11847\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__11842\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__11839\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__1673\ : IoInMux
    port map (
            O => \N__11832\,
            I => \N__11829\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__11829\,
            I => \N__11826\
        );

    \I__1671\ : IoSpan4Mux
    port map (
            O => \N__11826\,
            I => \N__11823\
        );

    \I__1670\ : IoSpan4Mux
    port map (
            O => \N__11823\,
            I => \N__11820\
        );

    \I__1669\ : Sp12to4
    port map (
            O => \N__11820\,
            I => \N__11817\
        );

    \I__1668\ : Span12Mux_h
    port map (
            O => \N__11817\,
            I => \N__11809\
        );

    \I__1667\ : InMux
    port map (
            O => \N__11816\,
            I => \N__11804\
        );

    \I__1666\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11804\
        );

    \I__1665\ : InMux
    port map (
            O => \N__11814\,
            I => \N__11799\
        );

    \I__1664\ : InMux
    port map (
            O => \N__11813\,
            I => \N__11799\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11796\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__11809\,
            I => \ADV_HSYNC_c\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__11804\,
            I => \ADV_HSYNC_c\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__11799\,
            I => \ADV_HSYNC_c\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__11796\,
            I => \ADV_HSYNC_c\
        );

    \I__1658\ : InMux
    port map (
            O => \N__11787\,
            I => \N__11781\
        );

    \I__1657\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11776\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11785\,
            I => \N__11776\
        );

    \I__1655\ : InMux
    port map (
            O => \N__11784\,
            I => \N__11773\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__11781\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__11776\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__11773\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__11766\,
            I => \transmit_module.n3675_cascade_\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__11763\,
            I => \transmit_module.video_signal_controller.n6_adj_622_cascade_\
        );

    \I__1649\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11754\
        );

    \I__1648\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11747\
        );

    \I__1647\ : InMux
    port map (
            O => \N__11758\,
            I => \N__11747\
        );

    \I__1646\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11747\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__11754\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__11747\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11736\
        );

    \I__1642\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11733\
        );

    \I__1641\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11728\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11728\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__11736\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11733\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__11728\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__11721\,
            I => \transmit_module.video_signal_controller.n3482_cascade_\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11718\,
            I => \N__11713\
        );

    \I__1634\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11708\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11708\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__11713\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__11708\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11698\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11693\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11693\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__11698\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__11693\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__11688\,
            I => \transmit_module.video_signal_controller.n6_cascade_\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11679\
        );

    \I__1623\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11679\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__11679\,
            I => \transmit_module.video_signal_controller.n2016\
        );

    \I__1621\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11672\
        );

    \I__1620\ : InMux
    port map (
            O => \N__11675\,
            I => \N__11669\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__11672\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__11669\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__1617\ : InMux
    port map (
            O => \N__11664\,
            I => \N__11660\
        );

    \I__1616\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11657\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__11660\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__11657\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__1613\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11649\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__11649\,
            I => \transmit_module.Y_DELTA_PATTERN_20\
        );

    \I__1611\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11643\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__11643\,
            I => \transmit_module.Y_DELTA_PATTERN_21\
        );

    \I__1609\ : InMux
    port map (
            O => \N__11640\,
            I => \N__11637\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__11637\,
            I => \transmit_module.Y_DELTA_PATTERN_22\
        );

    \I__1607\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11631\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__11631\,
            I => \transmit_module.Y_DELTA_PATTERN_24\
        );

    \I__1605\ : InMux
    port map (
            O => \N__11628\,
            I => \N__11625\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__11625\,
            I => \transmit_module.Y_DELTA_PATTERN_23\
        );

    \I__1603\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11619\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__11619\,
            I => \N__11616\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__11616\,
            I => \transmit_module.X_DELTA_PATTERN_13\
        );

    \I__1600\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11610\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__11610\,
            I => \transmit_module.X_DELTA_PATTERN_14\
        );

    \I__1598\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11604\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__11604\,
            I => \N__11601\
        );

    \I__1596\ : Odrv12
    port map (
            O => \N__11601\,
            I => \transmit_module.X_DELTA_PATTERN_6\
        );

    \I__1595\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11595\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__11595\,
            I => \transmit_module.X_DELTA_PATTERN_5\
        );

    \I__1593\ : InMux
    port map (
            O => \N__11592\,
            I => \N__11589\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11589\,
            I => \transmit_module.X_DELTA_PATTERN_4\
        );

    \I__1591\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11583\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__11583\,
            I => \transmit_module.ADDR_Y_COMPONENT_3\
        );

    \I__1589\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11577\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11574\
        );

    \I__1587\ : Span4Mux_h
    port map (
            O => \N__11574\,
            I => \N__11571\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__11571\,
            I => \N__11568\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__11568\,
            I => \line_buffer.n568\
        );

    \I__1584\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11562\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__11562\,
            I => \N__11559\
        );

    \I__1582\ : Span12Mux_v
    port map (
            O => \N__11559\,
            I => \N__11556\
        );

    \I__1581\ : Span12Mux_v
    port map (
            O => \N__11556\,
            I => \N__11553\
        );

    \I__1580\ : Span12Mux_h
    port map (
            O => \N__11553\,
            I => \N__11550\
        );

    \I__1579\ : Odrv12
    port map (
            O => \N__11550\,
            I => \line_buffer.n560\
        );

    \I__1578\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11544\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__11544\,
            I => \N__11541\
        );

    \I__1576\ : Span4Mux_h
    port map (
            O => \N__11541\,
            I => \N__11538\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__11538\,
            I => \line_buffer.n3530\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__11535\,
            I => \line_buffer.n3531_cascade_\
        );

    \I__1573\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11529\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__11529\,
            I => \line_buffer.n3617\
        );

    \I__1571\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11523\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__11523\,
            I => \TX_DATA_7\
        );

    \I__1569\ : IoInMux
    port map (
            O => \N__11520\,
            I => \N__11515\
        );

    \I__1568\ : IoInMux
    port map (
            O => \N__11519\,
            I => \N__11512\
        );

    \I__1567\ : IoInMux
    port map (
            O => \N__11518\,
            I => \N__11509\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__11515\,
            I => \N__11506\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__11512\,
            I => \N__11503\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__11509\,
            I => \N__11500\
        );

    \I__1563\ : IoSpan4Mux
    port map (
            O => \N__11506\,
            I => \N__11497\
        );

    \I__1562\ : IoSpan4Mux
    port map (
            O => \N__11503\,
            I => \N__11494\
        );

    \I__1561\ : Span12Mux_s10_v
    port map (
            O => \N__11500\,
            I => \N__11491\
        );

    \I__1560\ : Sp12to4
    port map (
            O => \N__11497\,
            I => \N__11488\
        );

    \I__1559\ : Span4Mux_s3_v
    port map (
            O => \N__11494\,
            I => \N__11485\
        );

    \I__1558\ : Span12Mux_h
    port map (
            O => \N__11491\,
            I => \N__11482\
        );

    \I__1557\ : Span12Mux_h
    port map (
            O => \N__11488\,
            I => \N__11479\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__11485\,
            I => \N__11476\
        );

    \I__1555\ : Odrv12
    port map (
            O => \N__11482\,
            I => \ADV_B_c\
        );

    \I__1554\ : Odrv12
    port map (
            O => \N__11479\,
            I => \ADV_B_c\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__11476\,
            I => \ADV_B_c\
        );

    \I__1552\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11466\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__11466\,
            I => \N__11463\
        );

    \I__1550\ : Span12Mux_h
    port map (
            O => \N__11463\,
            I => \N__11460\
        );

    \I__1549\ : Odrv12
    port map (
            O => \N__11460\,
            I => \transmit_module.Y_DELTA_PATTERN_26\
        );

    \I__1548\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11454\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__11454\,
            I => \transmit_module.Y_DELTA_PATTERN_25\
        );

    \I__1546\ : InMux
    port map (
            O => \N__11451\,
            I => \N__11448\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__11448\,
            I => \transmit_module.Y_DELTA_PATTERN_19\
        );

    \I__1544\ : InMux
    port map (
            O => \N__11445\,
            I => \N__11442\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__11442\,
            I => \transmit_module.n139\
        );

    \I__1542\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11435\
        );

    \I__1541\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11432\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__11435\,
            I => \transmit_module.n108\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__11432\,
            I => \transmit_module.n108\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__11427\,
            I => \transmit_module.n139_cascade_\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__11424\,
            I => \N__11421\
        );

    \I__1536\ : CascadeBuf
    port map (
            O => \N__11421\,
            I => \N__11417\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__11420\,
            I => \N__11414\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__11417\,
            I => \N__11411\
        );

    \I__1533\ : CascadeBuf
    port map (
            O => \N__11414\,
            I => \N__11408\
        );

    \I__1532\ : CascadeBuf
    port map (
            O => \N__11411\,
            I => \N__11405\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__11408\,
            I => \N__11402\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__11405\,
            I => \N__11399\
        );

    \I__1529\ : CascadeBuf
    port map (
            O => \N__11402\,
            I => \N__11396\
        );

    \I__1528\ : CascadeBuf
    port map (
            O => \N__11399\,
            I => \N__11393\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__11396\,
            I => \N__11390\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__11393\,
            I => \N__11387\
        );

    \I__1525\ : CascadeBuf
    port map (
            O => \N__11390\,
            I => \N__11384\
        );

    \I__1524\ : CascadeBuf
    port map (
            O => \N__11387\,
            I => \N__11381\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__11384\,
            I => \N__11378\
        );

    \I__1522\ : CascadeMux
    port map (
            O => \N__11381\,
            I => \N__11375\
        );

    \I__1521\ : CascadeBuf
    port map (
            O => \N__11378\,
            I => \N__11372\
        );

    \I__1520\ : CascadeBuf
    port map (
            O => \N__11375\,
            I => \N__11369\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__11372\,
            I => \N__11366\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__11369\,
            I => \N__11363\
        );

    \I__1517\ : CascadeBuf
    port map (
            O => \N__11366\,
            I => \N__11360\
        );

    \I__1516\ : CascadeBuf
    port map (
            O => \N__11363\,
            I => \N__11357\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__11360\,
            I => \N__11354\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__11357\,
            I => \N__11351\
        );

    \I__1513\ : CascadeBuf
    port map (
            O => \N__11354\,
            I => \N__11348\
        );

    \I__1512\ : CascadeBuf
    port map (
            O => \N__11351\,
            I => \N__11345\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__11348\,
            I => \N__11342\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__11345\,
            I => \N__11339\
        );

    \I__1509\ : CascadeBuf
    port map (
            O => \N__11342\,
            I => \N__11336\
        );

    \I__1508\ : CascadeBuf
    port map (
            O => \N__11339\,
            I => \N__11333\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__11336\,
            I => \N__11330\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__11333\,
            I => \N__11327\
        );

    \I__1505\ : CascadeBuf
    port map (
            O => \N__11330\,
            I => \N__11324\
        );

    \I__1504\ : CascadeBuf
    port map (
            O => \N__11327\,
            I => \N__11321\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__11324\,
            I => \N__11318\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__11321\,
            I => \N__11315\
        );

    \I__1501\ : CascadeBuf
    port map (
            O => \N__11318\,
            I => \N__11312\
        );

    \I__1500\ : CascadeBuf
    port map (
            O => \N__11315\,
            I => \N__11309\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__11312\,
            I => \N__11306\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__11309\,
            I => \N__11303\
        );

    \I__1497\ : CascadeBuf
    port map (
            O => \N__11306\,
            I => \N__11300\
        );

    \I__1496\ : CascadeBuf
    port map (
            O => \N__11303\,
            I => \N__11297\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__11300\,
            I => \N__11294\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__11297\,
            I => \N__11291\
        );

    \I__1493\ : CascadeBuf
    port map (
            O => \N__11294\,
            I => \N__11288\
        );

    \I__1492\ : CascadeBuf
    port map (
            O => \N__11291\,
            I => \N__11285\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__11288\,
            I => \N__11282\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__11285\,
            I => \N__11279\
        );

    \I__1489\ : CascadeBuf
    port map (
            O => \N__11282\,
            I => \N__11276\
        );

    \I__1488\ : CascadeBuf
    port map (
            O => \N__11279\,
            I => \N__11273\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__11276\,
            I => \N__11270\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__11273\,
            I => \N__11267\
        );

    \I__1485\ : CascadeBuf
    port map (
            O => \N__11270\,
            I => \N__11264\
        );

    \I__1484\ : CascadeBuf
    port map (
            O => \N__11267\,
            I => \N__11261\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__11264\,
            I => \N__11258\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__11261\,
            I => \N__11255\
        );

    \I__1481\ : CascadeBuf
    port map (
            O => \N__11258\,
            I => \N__11252\
        );

    \I__1480\ : CascadeBuf
    port map (
            O => \N__11255\,
            I => \N__11249\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__11252\,
            I => \N__11246\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__11249\,
            I => \N__11243\
        );

    \I__1477\ : CascadeBuf
    port map (
            O => \N__11246\,
            I => \N__11240\
        );

    \I__1476\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11237\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__11240\,
            I => \N__11234\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__11237\,
            I => \N__11231\
        );

    \I__1473\ : InMux
    port map (
            O => \N__11234\,
            I => \N__11228\
        );

    \I__1472\ : Span4Mux_s3_v
    port map (
            O => \N__11231\,
            I => \N__11225\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__11228\,
            I => \N__11222\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__11225\,
            I => \N__11219\
        );

    \I__1469\ : Span12Mux_s10_v
    port map (
            O => \N__11222\,
            I => \N__11216\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__11219\,
            I => \N__11213\
        );

    \I__1467\ : Span12Mux_h
    port map (
            O => \N__11216\,
            I => \N__11210\
        );

    \I__1466\ : Span4Mux_h
    port map (
            O => \N__11213\,
            I => \N__11207\
        );

    \I__1465\ : Odrv12
    port map (
            O => \N__11210\,
            I => n20
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__11207\,
            I => n20
        );

    \I__1463\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11199\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__11199\,
            I => \N__11196\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__11196\,
            I => \N__11193\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__11193\,
            I => \transmit_module.ADDR_Y_COMPONENT_10\
        );

    \I__1459\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11187\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__11187\,
            I => \N__11184\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__11184\,
            I => \transmit_module.n145\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__11181\,
            I => \N__11178\
        );

    \I__1455\ : CascadeBuf
    port map (
            O => \N__11178\,
            I => \N__11175\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__11175\,
            I => \N__11172\
        );

    \I__1453\ : CascadeBuf
    port map (
            O => \N__11172\,
            I => \N__11168\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__11171\,
            I => \N__11165\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__11168\,
            I => \N__11162\
        );

    \I__1450\ : CascadeBuf
    port map (
            O => \N__11165\,
            I => \N__11159\
        );

    \I__1449\ : CascadeBuf
    port map (
            O => \N__11162\,
            I => \N__11156\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__11159\,
            I => \N__11153\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__11156\,
            I => \N__11150\
        );

    \I__1446\ : CascadeBuf
    port map (
            O => \N__11153\,
            I => \N__11147\
        );

    \I__1445\ : CascadeBuf
    port map (
            O => \N__11150\,
            I => \N__11144\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__11147\,
            I => \N__11141\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__11144\,
            I => \N__11138\
        );

    \I__1442\ : CascadeBuf
    port map (
            O => \N__11141\,
            I => \N__11135\
        );

    \I__1441\ : CascadeBuf
    port map (
            O => \N__11138\,
            I => \N__11132\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__11135\,
            I => \N__11129\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__11132\,
            I => \N__11126\
        );

    \I__1438\ : CascadeBuf
    port map (
            O => \N__11129\,
            I => \N__11123\
        );

    \I__1437\ : CascadeBuf
    port map (
            O => \N__11126\,
            I => \N__11120\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__11123\,
            I => \N__11117\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__11120\,
            I => \N__11114\
        );

    \I__1434\ : CascadeBuf
    port map (
            O => \N__11117\,
            I => \N__11111\
        );

    \I__1433\ : CascadeBuf
    port map (
            O => \N__11114\,
            I => \N__11108\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__11111\,
            I => \N__11105\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__11108\,
            I => \N__11102\
        );

    \I__1430\ : CascadeBuf
    port map (
            O => \N__11105\,
            I => \N__11099\
        );

    \I__1429\ : CascadeBuf
    port map (
            O => \N__11102\,
            I => \N__11096\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__11099\,
            I => \N__11093\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__11096\,
            I => \N__11090\
        );

    \I__1426\ : CascadeBuf
    port map (
            O => \N__11093\,
            I => \N__11087\
        );

    \I__1425\ : CascadeBuf
    port map (
            O => \N__11090\,
            I => \N__11084\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__11087\,
            I => \N__11081\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__11084\,
            I => \N__11078\
        );

    \I__1422\ : CascadeBuf
    port map (
            O => \N__11081\,
            I => \N__11075\
        );

    \I__1421\ : CascadeBuf
    port map (
            O => \N__11078\,
            I => \N__11072\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__11075\,
            I => \N__11069\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__11072\,
            I => \N__11066\
        );

    \I__1418\ : CascadeBuf
    port map (
            O => \N__11069\,
            I => \N__11063\
        );

    \I__1417\ : CascadeBuf
    port map (
            O => \N__11066\,
            I => \N__11060\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__11063\,
            I => \N__11057\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__11060\,
            I => \N__11054\
        );

    \I__1414\ : CascadeBuf
    port map (
            O => \N__11057\,
            I => \N__11051\
        );

    \I__1413\ : CascadeBuf
    port map (
            O => \N__11054\,
            I => \N__11048\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__11051\,
            I => \N__11045\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__11048\,
            I => \N__11042\
        );

    \I__1410\ : CascadeBuf
    port map (
            O => \N__11045\,
            I => \N__11039\
        );

    \I__1409\ : CascadeBuf
    port map (
            O => \N__11042\,
            I => \N__11036\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__11039\,
            I => \N__11033\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__11036\,
            I => \N__11030\
        );

    \I__1406\ : CascadeBuf
    port map (
            O => \N__11033\,
            I => \N__11027\
        );

    \I__1405\ : CascadeBuf
    port map (
            O => \N__11030\,
            I => \N__11024\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__11027\,
            I => \N__11021\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__11024\,
            I => \N__11018\
        );

    \I__1402\ : CascadeBuf
    port map (
            O => \N__11021\,
            I => \N__11015\
        );

    \I__1401\ : CascadeBuf
    port map (
            O => \N__11018\,
            I => \N__11012\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__11015\,
            I => \N__11009\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__11012\,
            I => \N__11006\
        );

    \I__1398\ : CascadeBuf
    port map (
            O => \N__11009\,
            I => \N__11003\
        );

    \I__1397\ : InMux
    port map (
            O => \N__11006\,
            I => \N__11000\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__11003\,
            I => \N__10997\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__11000\,
            I => \N__10994\
        );

    \I__1394\ : CascadeBuf
    port map (
            O => \N__10997\,
            I => \N__10991\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__10994\,
            I => \N__10988\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__10991\,
            I => \N__10985\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__10988\,
            I => \N__10982\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10979\
        );

    \I__1389\ : Span4Mux_v
    port map (
            O => \N__10982\,
            I => \N__10976\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__10979\,
            I => \N__10973\
        );

    \I__1387\ : Span4Mux_h
    port map (
            O => \N__10976\,
            I => \N__10970\
        );

    \I__1386\ : Sp12to4
    port map (
            O => \N__10973\,
            I => \N__10967\
        );

    \I__1385\ : Span4Mux_h
    port map (
            O => \N__10970\,
            I => \N__10964\
        );

    \I__1384\ : Span12Mux_v
    port map (
            O => \N__10967\,
            I => \N__10961\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__10964\,
            I => n26
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__10961\,
            I => n26
        );

    \I__1381\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10953\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__10953\,
            I => \N__10949\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10946\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__10949\,
            I => \transmit_module.n114\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10946\,
            I => \transmit_module.n114\
        );

    \I__1376\ : InMux
    port map (
            O => \N__10941\,
            I => \N__10938\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__10938\,
            I => \N__10935\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__10935\,
            I => \transmit_module.n144\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__10932\,
            I => \transmit_module.n144_cascade_\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__10929\,
            I => \N__10926\
        );

    \I__1371\ : CascadeBuf
    port map (
            O => \N__10926\,
            I => \N__10923\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__10923\,
            I => \N__10920\
        );

    \I__1369\ : CascadeBuf
    port map (
            O => \N__10920\,
            I => \N__10916\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__10919\,
            I => \N__10913\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__10916\,
            I => \N__10910\
        );

    \I__1366\ : CascadeBuf
    port map (
            O => \N__10913\,
            I => \N__10907\
        );

    \I__1365\ : CascadeBuf
    port map (
            O => \N__10910\,
            I => \N__10904\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__10907\,
            I => \N__10901\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__10904\,
            I => \N__10898\
        );

    \I__1362\ : CascadeBuf
    port map (
            O => \N__10901\,
            I => \N__10895\
        );

    \I__1361\ : CascadeBuf
    port map (
            O => \N__10898\,
            I => \N__10892\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__10895\,
            I => \N__10889\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__10892\,
            I => \N__10886\
        );

    \I__1358\ : CascadeBuf
    port map (
            O => \N__10889\,
            I => \N__10883\
        );

    \I__1357\ : CascadeBuf
    port map (
            O => \N__10886\,
            I => \N__10880\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__10883\,
            I => \N__10877\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__10880\,
            I => \N__10874\
        );

    \I__1354\ : CascadeBuf
    port map (
            O => \N__10877\,
            I => \N__10871\
        );

    \I__1353\ : CascadeBuf
    port map (
            O => \N__10874\,
            I => \N__10868\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__10871\,
            I => \N__10865\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__10868\,
            I => \N__10862\
        );

    \I__1350\ : CascadeBuf
    port map (
            O => \N__10865\,
            I => \N__10859\
        );

    \I__1349\ : CascadeBuf
    port map (
            O => \N__10862\,
            I => \N__10856\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__10859\,
            I => \N__10853\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__10856\,
            I => \N__10850\
        );

    \I__1346\ : CascadeBuf
    port map (
            O => \N__10853\,
            I => \N__10847\
        );

    \I__1345\ : CascadeBuf
    port map (
            O => \N__10850\,
            I => \N__10844\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__10847\,
            I => \N__10841\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__10844\,
            I => \N__10838\
        );

    \I__1342\ : CascadeBuf
    port map (
            O => \N__10841\,
            I => \N__10835\
        );

    \I__1341\ : CascadeBuf
    port map (
            O => \N__10838\,
            I => \N__10832\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__10835\,
            I => \N__10829\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__10832\,
            I => \N__10826\
        );

    \I__1338\ : CascadeBuf
    port map (
            O => \N__10829\,
            I => \N__10823\
        );

    \I__1337\ : CascadeBuf
    port map (
            O => \N__10826\,
            I => \N__10820\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__10823\,
            I => \N__10817\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__10820\,
            I => \N__10814\
        );

    \I__1334\ : CascadeBuf
    port map (
            O => \N__10817\,
            I => \N__10811\
        );

    \I__1333\ : CascadeBuf
    port map (
            O => \N__10814\,
            I => \N__10808\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__10811\,
            I => \N__10805\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__10808\,
            I => \N__10802\
        );

    \I__1330\ : CascadeBuf
    port map (
            O => \N__10805\,
            I => \N__10799\
        );

    \I__1329\ : CascadeBuf
    port map (
            O => \N__10802\,
            I => \N__10796\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__10799\,
            I => \N__10793\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__10796\,
            I => \N__10790\
        );

    \I__1326\ : CascadeBuf
    port map (
            O => \N__10793\,
            I => \N__10787\
        );

    \I__1325\ : CascadeBuf
    port map (
            O => \N__10790\,
            I => \N__10784\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__10787\,
            I => \N__10781\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__10784\,
            I => \N__10778\
        );

    \I__1322\ : CascadeBuf
    port map (
            O => \N__10781\,
            I => \N__10775\
        );

    \I__1321\ : CascadeBuf
    port map (
            O => \N__10778\,
            I => \N__10772\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__10775\,
            I => \N__10769\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__10772\,
            I => \N__10766\
        );

    \I__1318\ : CascadeBuf
    port map (
            O => \N__10769\,
            I => \N__10763\
        );

    \I__1317\ : CascadeBuf
    port map (
            O => \N__10766\,
            I => \N__10760\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__10763\,
            I => \N__10757\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__10760\,
            I => \N__10754\
        );

    \I__1314\ : CascadeBuf
    port map (
            O => \N__10757\,
            I => \N__10751\
        );

    \I__1313\ : InMux
    port map (
            O => \N__10754\,
            I => \N__10748\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__10751\,
            I => \N__10745\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10748\,
            I => \N__10742\
        );

    \I__1310\ : CascadeBuf
    port map (
            O => \N__10745\,
            I => \N__10739\
        );

    \I__1309\ : Span4Mux_v
    port map (
            O => \N__10742\,
            I => \N__10736\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__10739\,
            I => \N__10733\
        );

    \I__1307\ : Span4Mux_v
    port map (
            O => \N__10736\,
            I => \N__10730\
        );

    \I__1306\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10727\
        );

    \I__1305\ : Span4Mux_h
    port map (
            O => \N__10730\,
            I => \N__10724\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__10727\,
            I => \N__10721\
        );

    \I__1303\ : Span4Mux_h
    port map (
            O => \N__10724\,
            I => \N__10718\
        );

    \I__1302\ : Span4Mux_v
    port map (
            O => \N__10721\,
            I => \N__10715\
        );

    \I__1301\ : Span4Mux_h
    port map (
            O => \N__10718\,
            I => \N__10710\
        );

    \I__1300\ : Span4Mux_h
    port map (
            O => \N__10715\,
            I => \N__10710\
        );

    \I__1299\ : Sp12to4
    port map (
            O => \N__10710\,
            I => \N__10707\
        );

    \I__1298\ : Odrv12
    port map (
            O => \N__10707\,
            I => n25
        );

    \I__1297\ : InMux
    port map (
            O => \N__10704\,
            I => \N__10701\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__10701\,
            I => \N__10697\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10694\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__10697\,
            I => \transmit_module.n113\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__10694\,
            I => \transmit_module.n113\
        );

    \I__1292\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10686\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__10686\,
            I => \transmit_module.ADDR_Y_COMPONENT_2\
        );

    \I__1290\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10677\
        );

    \I__1289\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10677\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__10677\,
            I => \transmit_module.n115\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10671\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__10671\,
            I => \transmit_module.n142\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__10668\,
            I => \transmit_module.n142_cascade_\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__10665\,
            I => \N__10662\
        );

    \I__1283\ : CascadeBuf
    port map (
            O => \N__10662\,
            I => \N__10659\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__10659\,
            I => \N__10656\
        );

    \I__1281\ : CascadeBuf
    port map (
            O => \N__10656\,
            I => \N__10652\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__10655\,
            I => \N__10649\
        );

    \I__1279\ : CascadeMux
    port map (
            O => \N__10652\,
            I => \N__10646\
        );

    \I__1278\ : CascadeBuf
    port map (
            O => \N__10649\,
            I => \N__10643\
        );

    \I__1277\ : CascadeBuf
    port map (
            O => \N__10646\,
            I => \N__10640\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__10643\,
            I => \N__10637\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__10640\,
            I => \N__10634\
        );

    \I__1274\ : CascadeBuf
    port map (
            O => \N__10637\,
            I => \N__10631\
        );

    \I__1273\ : CascadeBuf
    port map (
            O => \N__10634\,
            I => \N__10628\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__10631\,
            I => \N__10625\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__10628\,
            I => \N__10622\
        );

    \I__1270\ : CascadeBuf
    port map (
            O => \N__10625\,
            I => \N__10619\
        );

    \I__1269\ : CascadeBuf
    port map (
            O => \N__10622\,
            I => \N__10616\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__10619\,
            I => \N__10613\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__10616\,
            I => \N__10610\
        );

    \I__1266\ : CascadeBuf
    port map (
            O => \N__10613\,
            I => \N__10607\
        );

    \I__1265\ : CascadeBuf
    port map (
            O => \N__10610\,
            I => \N__10604\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__10607\,
            I => \N__10601\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__10604\,
            I => \N__10598\
        );

    \I__1262\ : CascadeBuf
    port map (
            O => \N__10601\,
            I => \N__10595\
        );

    \I__1261\ : CascadeBuf
    port map (
            O => \N__10598\,
            I => \N__10592\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__10595\,
            I => \N__10589\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__10592\,
            I => \N__10586\
        );

    \I__1258\ : CascadeBuf
    port map (
            O => \N__10589\,
            I => \N__10583\
        );

    \I__1257\ : CascadeBuf
    port map (
            O => \N__10586\,
            I => \N__10580\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__10583\,
            I => \N__10577\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__10580\,
            I => \N__10574\
        );

    \I__1254\ : CascadeBuf
    port map (
            O => \N__10577\,
            I => \N__10571\
        );

    \I__1253\ : CascadeBuf
    port map (
            O => \N__10574\,
            I => \N__10568\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__10571\,
            I => \N__10565\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__10568\,
            I => \N__10562\
        );

    \I__1250\ : CascadeBuf
    port map (
            O => \N__10565\,
            I => \N__10559\
        );

    \I__1249\ : CascadeBuf
    port map (
            O => \N__10562\,
            I => \N__10556\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__10559\,
            I => \N__10553\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__10556\,
            I => \N__10550\
        );

    \I__1246\ : CascadeBuf
    port map (
            O => \N__10553\,
            I => \N__10547\
        );

    \I__1245\ : CascadeBuf
    port map (
            O => \N__10550\,
            I => \N__10544\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__10547\,
            I => \N__10541\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__10544\,
            I => \N__10538\
        );

    \I__1242\ : CascadeBuf
    port map (
            O => \N__10541\,
            I => \N__10535\
        );

    \I__1241\ : CascadeBuf
    port map (
            O => \N__10538\,
            I => \N__10532\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__10535\,
            I => \N__10529\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__10532\,
            I => \N__10526\
        );

    \I__1238\ : CascadeBuf
    port map (
            O => \N__10529\,
            I => \N__10523\
        );

    \I__1237\ : CascadeBuf
    port map (
            O => \N__10526\,
            I => \N__10520\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__10523\,
            I => \N__10517\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__10520\,
            I => \N__10514\
        );

    \I__1234\ : CascadeBuf
    port map (
            O => \N__10517\,
            I => \N__10511\
        );

    \I__1233\ : CascadeBuf
    port map (
            O => \N__10514\,
            I => \N__10508\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__10511\,
            I => \N__10505\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__10508\,
            I => \N__10502\
        );

    \I__1230\ : CascadeBuf
    port map (
            O => \N__10505\,
            I => \N__10499\
        );

    \I__1229\ : CascadeBuf
    port map (
            O => \N__10502\,
            I => \N__10496\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__10499\,
            I => \N__10493\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__10496\,
            I => \N__10490\
        );

    \I__1226\ : CascadeBuf
    port map (
            O => \N__10493\,
            I => \N__10487\
        );

    \I__1225\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10484\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__10487\,
            I => \N__10481\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__10484\,
            I => \N__10478\
        );

    \I__1222\ : CascadeBuf
    port map (
            O => \N__10481\,
            I => \N__10475\
        );

    \I__1221\ : Span4Mux_v
    port map (
            O => \N__10478\,
            I => \N__10472\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__10475\,
            I => \N__10469\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__10472\,
            I => \N__10466\
        );

    \I__1218\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10463\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__10466\,
            I => \N__10460\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__10463\,
            I => \N__10457\
        );

    \I__1215\ : Span4Mux_h
    port map (
            O => \N__10460\,
            I => \N__10454\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__10457\,
            I => \N__10451\
        );

    \I__1213\ : Span4Mux_h
    port map (
            O => \N__10454\,
            I => \N__10446\
        );

    \I__1212\ : Span4Mux_h
    port map (
            O => \N__10451\,
            I => \N__10446\
        );

    \I__1211\ : Sp12to4
    port map (
            O => \N__10446\,
            I => \N__10443\
        );

    \I__1210\ : Odrv12
    port map (
            O => \N__10443\,
            I => n23
        );

    \I__1209\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10436\
        );

    \I__1208\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10433\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__10436\,
            I => \transmit_module.n111\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__10433\,
            I => \transmit_module.n111\
        );

    \I__1205\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10425\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__10425\,
            I => \transmit_module.n138\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__10422\,
            I => \transmit_module.n138_cascade_\
        );

    \I__1202\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10416\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__10416\,
            I => \transmit_module.n107\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__10413\,
            I => \N__10410\
        );

    \I__1199\ : CascadeBuf
    port map (
            O => \N__10410\,
            I => \N__10407\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__10407\,
            I => \N__10403\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__10406\,
            I => \N__10400\
        );

    \I__1196\ : CascadeBuf
    port map (
            O => \N__10403\,
            I => \N__10397\
        );

    \I__1195\ : CascadeBuf
    port map (
            O => \N__10400\,
            I => \N__10394\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__10397\,
            I => \N__10391\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__10394\,
            I => \N__10388\
        );

    \I__1192\ : CascadeBuf
    port map (
            O => \N__10391\,
            I => \N__10385\
        );

    \I__1191\ : CascadeBuf
    port map (
            O => \N__10388\,
            I => \N__10382\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__10385\,
            I => \N__10379\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__10382\,
            I => \N__10376\
        );

    \I__1188\ : CascadeBuf
    port map (
            O => \N__10379\,
            I => \N__10373\
        );

    \I__1187\ : CascadeBuf
    port map (
            O => \N__10376\,
            I => \N__10370\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__10373\,
            I => \N__10367\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__10370\,
            I => \N__10364\
        );

    \I__1184\ : CascadeBuf
    port map (
            O => \N__10367\,
            I => \N__10361\
        );

    \I__1183\ : CascadeBuf
    port map (
            O => \N__10364\,
            I => \N__10358\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__10361\,
            I => \N__10355\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__10358\,
            I => \N__10352\
        );

    \I__1180\ : CascadeBuf
    port map (
            O => \N__10355\,
            I => \N__10349\
        );

    \I__1179\ : CascadeBuf
    port map (
            O => \N__10352\,
            I => \N__10346\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__10349\,
            I => \N__10343\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__10346\,
            I => \N__10340\
        );

    \I__1176\ : CascadeBuf
    port map (
            O => \N__10343\,
            I => \N__10337\
        );

    \I__1175\ : CascadeBuf
    port map (
            O => \N__10340\,
            I => \N__10334\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__10337\,
            I => \N__10331\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \N__10328\
        );

    \I__1172\ : CascadeBuf
    port map (
            O => \N__10331\,
            I => \N__10325\
        );

    \I__1171\ : CascadeBuf
    port map (
            O => \N__10328\,
            I => \N__10322\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__10325\,
            I => \N__10319\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__10322\,
            I => \N__10316\
        );

    \I__1168\ : CascadeBuf
    port map (
            O => \N__10319\,
            I => \N__10313\
        );

    \I__1167\ : CascadeBuf
    port map (
            O => \N__10316\,
            I => \N__10310\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__10313\,
            I => \N__10307\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__10310\,
            I => \N__10304\
        );

    \I__1164\ : CascadeBuf
    port map (
            O => \N__10307\,
            I => \N__10301\
        );

    \I__1163\ : CascadeBuf
    port map (
            O => \N__10304\,
            I => \N__10298\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__10301\,
            I => \N__10295\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__10298\,
            I => \N__10292\
        );

    \I__1160\ : CascadeBuf
    port map (
            O => \N__10295\,
            I => \N__10289\
        );

    \I__1159\ : CascadeBuf
    port map (
            O => \N__10292\,
            I => \N__10286\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__10289\,
            I => \N__10283\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \N__10280\
        );

    \I__1156\ : CascadeBuf
    port map (
            O => \N__10283\,
            I => \N__10277\
        );

    \I__1155\ : CascadeBuf
    port map (
            O => \N__10280\,
            I => \N__10274\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__10277\,
            I => \N__10271\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__10274\,
            I => \N__10268\
        );

    \I__1152\ : CascadeBuf
    port map (
            O => \N__10271\,
            I => \N__10265\
        );

    \I__1151\ : CascadeBuf
    port map (
            O => \N__10268\,
            I => \N__10262\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__10265\,
            I => \N__10259\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__10262\,
            I => \N__10256\
        );

    \I__1148\ : CascadeBuf
    port map (
            O => \N__10259\,
            I => \N__10253\
        );

    \I__1147\ : CascadeBuf
    port map (
            O => \N__10256\,
            I => \N__10250\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__10253\,
            I => \N__10247\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__10250\,
            I => \N__10244\
        );

    \I__1144\ : CascadeBuf
    port map (
            O => \N__10247\,
            I => \N__10241\
        );

    \I__1143\ : CascadeBuf
    port map (
            O => \N__10244\,
            I => \N__10238\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__10241\,
            I => \N__10235\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__10238\,
            I => \N__10232\
        );

    \I__1140\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10229\
        );

    \I__1139\ : CascadeBuf
    port map (
            O => \N__10232\,
            I => \N__10226\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__10229\,
            I => \N__10223\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__10226\,
            I => \N__10220\
        );

    \I__1136\ : Span4Mux_v
    port map (
            O => \N__10223\,
            I => \N__10217\
        );

    \I__1135\ : InMux
    port map (
            O => \N__10220\,
            I => \N__10214\
        );

    \I__1134\ : Span4Mux_v
    port map (
            O => \N__10217\,
            I => \N__10211\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__10214\,
            I => \N__10208\
        );

    \I__1132\ : Span4Mux_v
    port map (
            O => \N__10211\,
            I => \N__10205\
        );

    \I__1131\ : Span4Mux_v
    port map (
            O => \N__10208\,
            I => \N__10202\
        );

    \I__1130\ : Span4Mux_h
    port map (
            O => \N__10205\,
            I => \N__10199\
        );

    \I__1129\ : Span4Mux_v
    port map (
            O => \N__10202\,
            I => \N__10196\
        );

    \I__1128\ : Span4Mux_h
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__10196\,
            I => \N__10190\
        );

    \I__1126\ : Span4Mux_h
    port map (
            O => \N__10193\,
            I => \N__10185\
        );

    \I__1125\ : Span4Mux_h
    port map (
            O => \N__10190\,
            I => \N__10185\
        );

    \I__1124\ : Odrv4
    port map (
            O => \N__10185\,
            I => n19
        );

    \I__1123\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10179\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__10179\,
            I => \transmit_module.n146\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__10176\,
            I => \transmit_module.n146_cascade_\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__10173\,
            I => \N__10169\
        );

    \I__1119\ : CascadeMux
    port map (
            O => \N__10172\,
            I => \N__10166\
        );

    \I__1118\ : CascadeBuf
    port map (
            O => \N__10169\,
            I => \N__10163\
        );

    \I__1117\ : CascadeBuf
    port map (
            O => \N__10166\,
            I => \N__10160\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__10163\,
            I => \N__10157\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__10160\,
            I => \N__10154\
        );

    \I__1114\ : CascadeBuf
    port map (
            O => \N__10157\,
            I => \N__10151\
        );

    \I__1113\ : CascadeBuf
    port map (
            O => \N__10154\,
            I => \N__10148\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__10151\,
            I => \N__10145\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__10148\,
            I => \N__10142\
        );

    \I__1110\ : CascadeBuf
    port map (
            O => \N__10145\,
            I => \N__10139\
        );

    \I__1109\ : CascadeBuf
    port map (
            O => \N__10142\,
            I => \N__10136\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__10139\,
            I => \N__10133\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__10136\,
            I => \N__10130\
        );

    \I__1106\ : CascadeBuf
    port map (
            O => \N__10133\,
            I => \N__10127\
        );

    \I__1105\ : CascadeBuf
    port map (
            O => \N__10130\,
            I => \N__10124\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__10127\,
            I => \N__10121\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__10124\,
            I => \N__10118\
        );

    \I__1102\ : CascadeBuf
    port map (
            O => \N__10121\,
            I => \N__10115\
        );

    \I__1101\ : CascadeBuf
    port map (
            O => \N__10118\,
            I => \N__10112\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__10115\,
            I => \N__10109\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__10112\,
            I => \N__10106\
        );

    \I__1098\ : CascadeBuf
    port map (
            O => \N__10109\,
            I => \N__10103\
        );

    \I__1097\ : CascadeBuf
    port map (
            O => \N__10106\,
            I => \N__10100\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__10103\,
            I => \N__10097\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__10100\,
            I => \N__10094\
        );

    \I__1094\ : CascadeBuf
    port map (
            O => \N__10097\,
            I => \N__10091\
        );

    \I__1093\ : CascadeBuf
    port map (
            O => \N__10094\,
            I => \N__10088\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__10091\,
            I => \N__10085\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__10088\,
            I => \N__10082\
        );

    \I__1090\ : CascadeBuf
    port map (
            O => \N__10085\,
            I => \N__10079\
        );

    \I__1089\ : CascadeBuf
    port map (
            O => \N__10082\,
            I => \N__10076\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__10079\,
            I => \N__10073\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__10076\,
            I => \N__10070\
        );

    \I__1086\ : CascadeBuf
    port map (
            O => \N__10073\,
            I => \N__10067\
        );

    \I__1085\ : CascadeBuf
    port map (
            O => \N__10070\,
            I => \N__10064\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__10067\,
            I => \N__10061\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__10064\,
            I => \N__10058\
        );

    \I__1082\ : CascadeBuf
    port map (
            O => \N__10061\,
            I => \N__10055\
        );

    \I__1081\ : CascadeBuf
    port map (
            O => \N__10058\,
            I => \N__10052\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__10055\,
            I => \N__10049\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__10052\,
            I => \N__10046\
        );

    \I__1078\ : CascadeBuf
    port map (
            O => \N__10049\,
            I => \N__10043\
        );

    \I__1077\ : CascadeBuf
    port map (
            O => \N__10046\,
            I => \N__10040\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__10043\,
            I => \N__10037\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__10040\,
            I => \N__10034\
        );

    \I__1074\ : CascadeBuf
    port map (
            O => \N__10037\,
            I => \N__10031\
        );

    \I__1073\ : CascadeBuf
    port map (
            O => \N__10034\,
            I => \N__10028\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__10031\,
            I => \N__10025\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__10028\,
            I => \N__10022\
        );

    \I__1070\ : CascadeBuf
    port map (
            O => \N__10025\,
            I => \N__10019\
        );

    \I__1069\ : CascadeBuf
    port map (
            O => \N__10022\,
            I => \N__10016\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__10019\,
            I => \N__10013\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__10016\,
            I => \N__10010\
        );

    \I__1066\ : CascadeBuf
    port map (
            O => \N__10013\,
            I => \N__10007\
        );

    \I__1065\ : CascadeBuf
    port map (
            O => \N__10010\,
            I => \N__10004\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__10007\,
            I => \N__10001\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__10004\,
            I => \N__9998\
        );

    \I__1062\ : CascadeBuf
    port map (
            O => \N__10001\,
            I => \N__9995\
        );

    \I__1061\ : CascadeBuf
    port map (
            O => \N__9998\,
            I => \N__9992\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__9995\,
            I => \N__9989\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__9992\,
            I => \N__9986\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9983\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9986\,
            I => \N__9980\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__9983\,
            I => \N__9977\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__9980\,
            I => \N__9974\
        );

    \I__1054\ : Span4Mux_v
    port map (
            O => \N__9977\,
            I => \N__9971\
        );

    \I__1053\ : Sp12to4
    port map (
            O => \N__9974\,
            I => \N__9968\
        );

    \I__1052\ : Span4Mux_v
    port map (
            O => \N__9971\,
            I => \N__9965\
        );

    \I__1051\ : Span12Mux_s10_v
    port map (
            O => \N__9968\,
            I => \N__9962\
        );

    \I__1050\ : Span4Mux_h
    port map (
            O => \N__9965\,
            I => \N__9959\
        );

    \I__1049\ : Span12Mux_h
    port map (
            O => \N__9962\,
            I => \N__9954\
        );

    \I__1048\ : Sp12to4
    port map (
            O => \N__9959\,
            I => \N__9954\
        );

    \I__1047\ : Odrv12
    port map (
            O => \N__9954\,
            I => n27
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__9951\,
            I => \transmit_module.n107_cascade_\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__9948\,
            I => \transmit_module.n145_cascade_\
        );

    \I__1044\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9942\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9942\,
            I => \transmit_module.video_signal_controller.n7\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9934\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9931\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9928\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__9934\,
            I => \N__9925\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9931\,
            I => \N__9922\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9928\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__9925\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__9922\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1034\ : CEMux
    port map (
            O => \N__9915\,
            I => \N__9909\
        );

    \I__1033\ : CEMux
    port map (
            O => \N__9914\,
            I => \N__9905\
        );

    \I__1032\ : CEMux
    port map (
            O => \N__9913\,
            I => \N__9901\
        );

    \I__1031\ : CEMux
    port map (
            O => \N__9912\,
            I => \N__9896\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__9909\,
            I => \N__9891\
        );

    \I__1029\ : CEMux
    port map (
            O => \N__9908\,
            I => \N__9888\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__9905\,
            I => \N__9885\
        );

    \I__1027\ : CEMux
    port map (
            O => \N__9904\,
            I => \N__9882\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__9901\,
            I => \N__9879\
        );

    \I__1025\ : CEMux
    port map (
            O => \N__9900\,
            I => \N__9876\
        );

    \I__1024\ : CEMux
    port map (
            O => \N__9899\,
            I => \N__9873\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9869\
        );

    \I__1022\ : CEMux
    port map (
            O => \N__9895\,
            I => \N__9866\
        );

    \I__1021\ : CEMux
    port map (
            O => \N__9894\,
            I => \N__9863\
        );

    \I__1020\ : Span4Mux_v
    port map (
            O => \N__9891\,
            I => \N__9854\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__9888\,
            I => \N__9854\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__9885\,
            I => \N__9854\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__9882\,
            I => \N__9854\
        );

    \I__1016\ : Span4Mux_v
    port map (
            O => \N__9879\,
            I => \N__9847\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__9876\,
            I => \N__9847\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__9873\,
            I => \N__9847\
        );

    \I__1013\ : CEMux
    port map (
            O => \N__9872\,
            I => \N__9844\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__9869\,
            I => \N__9837\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9866\,
            I => \N__9837\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9863\,
            I => \N__9837\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__9854\,
            I => \N__9834\
        );

    \I__1008\ : Span4Mux_h
    port map (
            O => \N__9847\,
            I => \N__9831\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__9844\,
            I => \N__9828\
        );

    \I__1006\ : Span4Mux_h
    port map (
            O => \N__9837\,
            I => \N__9825\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__9834\,
            I => \transmit_module.n3680\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__9831\,
            I => \transmit_module.n3680\
        );

    \I__1003\ : Odrv12
    port map (
            O => \N__9828\,
            I => \transmit_module.n3680\
        );

    \I__1002\ : Odrv4
    port map (
            O => \N__9825\,
            I => \transmit_module.n3680\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__9816\,
            I => \N__9812\
        );

    \I__1000\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9807\
        );

    \I__999\ : InMux
    port map (
            O => \N__9812\,
            I => \N__9804\
        );

    \I__998\ : InMux
    port map (
            O => \N__9811\,
            I => \N__9801\
        );

    \I__997\ : InMux
    port map (
            O => \N__9810\,
            I => \N__9798\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9807\,
            I => \N__9791\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__9804\,
            I => \N__9791\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__9801\,
            I => \N__9791\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9798\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__9791\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__9786\,
            I => \N__9782\
        );

    \I__990\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9775\
        );

    \I__989\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9775\
        );

    \I__988\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9772\
        );

    \I__987\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9769\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__9775\,
            I => \N__9764\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__9772\,
            I => \N__9764\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9769\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__983\ : Odrv4
    port map (
            O => \N__9764\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__982\ : InMux
    port map (
            O => \N__9759\,
            I => \N__9751\
        );

    \I__981\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9751\
        );

    \I__980\ : InMux
    port map (
            O => \N__9757\,
            I => \N__9748\
        );

    \I__979\ : InMux
    port map (
            O => \N__9756\,
            I => \N__9745\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9740\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__9748\,
            I => \N__9740\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__9745\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__9740\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__974\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9727\
        );

    \I__973\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9727\
        );

    \I__972\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9724\
        );

    \I__971\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9721\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__9727\,
            I => \N__9716\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__9724\,
            I => \N__9716\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__9721\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__9716\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__966\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9706\
        );

    \I__965\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9703\
        );

    \I__964\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9700\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__9706\,
            I => \N__9695\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9703\,
            I => \N__9695\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__9700\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__9695\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__9690\,
            I => \transmit_module.video_signal_controller.n2014_cascade_\
        );

    \I__958\ : InMux
    port map (
            O => \N__9687\,
            I => \N__9681\
        );

    \I__957\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9678\
        );

    \I__956\ : InMux
    port map (
            O => \N__9685\,
            I => \N__9675\
        );

    \I__955\ : InMux
    port map (
            O => \N__9684\,
            I => \N__9672\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9681\,
            I => \N__9667\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9667\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9675\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9672\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__9667\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__949\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9656\
        );

    \I__948\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9651\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9656\,
            I => \N__9648\
        );

    \I__946\ : InMux
    port map (
            O => \N__9655\,
            I => \N__9645\
        );

    \I__945\ : InMux
    port map (
            O => \N__9654\,
            I => \N__9642\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__9651\,
            I => \N__9639\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__9648\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__9645\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__9642\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__9639\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__939\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9627\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__9627\,
            I => \transmit_module.video_signal_controller.n3676\
        );

    \I__937\ : InMux
    port map (
            O => \N__9624\,
            I => \transmit_module.video_signal_controller.n3193\
        );

    \I__936\ : InMux
    port map (
            O => \N__9621\,
            I => \transmit_module.video_signal_controller.n3194\
        );

    \I__935\ : InMux
    port map (
            O => \N__9618\,
            I => \transmit_module.video_signal_controller.n3195\
        );

    \I__934\ : InMux
    port map (
            O => \N__9615\,
            I => \transmit_module.video_signal_controller.n3196\
        );

    \I__933\ : InMux
    port map (
            O => \N__9612\,
            I => \transmit_module.video_signal_controller.n3197\
        );

    \I__932\ : InMux
    port map (
            O => \N__9609\,
            I => \bfn_13_13_0_\
        );

    \I__931\ : InMux
    port map (
            O => \N__9606\,
            I => \transmit_module.video_signal_controller.n3199\
        );

    \I__930\ : InMux
    port map (
            O => \N__9603\,
            I => \transmit_module.video_signal_controller.n3200\
        );

    \I__929\ : InMux
    port map (
            O => \N__9600\,
            I => \transmit_module.video_signal_controller.n3201\
        );

    \I__928\ : SRMux
    port map (
            O => \N__9597\,
            I => \N__9594\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__9594\,
            I => \N__9590\
        );

    \I__926\ : SRMux
    port map (
            O => \N__9593\,
            I => \N__9587\
        );

    \I__925\ : Span4Mux_v
    port map (
            O => \N__9590\,
            I => \N__9582\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__9587\,
            I => \N__9582\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__9582\,
            I => \transmit_module.video_signal_controller.n2395\
        );

    \I__922\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9576\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__9576\,
            I => \transmit_module.Y_DELTA_PATTERN_17\
        );

    \I__920\ : InMux
    port map (
            O => \N__9573\,
            I => \N__9570\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__9570\,
            I => \transmit_module.Y_DELTA_PATTERN_16\
        );

    \I__918\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9564\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__9564\,
            I => \transmit_module.Y_DELTA_PATTERN_13\
        );

    \I__916\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9558\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__9558\,
            I => \transmit_module.Y_DELTA_PATTERN_15\
        );

    \I__914\ : InMux
    port map (
            O => \N__9555\,
            I => \N__9552\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__9552\,
            I => \transmit_module.Y_DELTA_PATTERN_14\
        );

    \I__912\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__9546\,
            I => \transmit_module.Y_DELTA_PATTERN_18\
        );

    \I__910\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9540\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__9540\,
            I => \N__9537\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__9537\,
            I => \tvp_video_buffer.BUFFER_1_4\
        );

    \I__907\ : InMux
    port map (
            O => \N__9534\,
            I => \N__9531\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__9531\,
            I => \N__9528\
        );

    \I__905\ : Span4Mux_s1_v
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__904\ : Span4Mux_v
    port map (
            O => \N__9525\,
            I => \N__9521\
        );

    \I__903\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9516\
        );

    \I__902\ : Span4Mux_v
    port map (
            O => \N__9521\,
            I => \N__9510\
        );

    \I__901\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9507\
        );

    \I__900\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9504\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__9516\,
            I => \N__9500\
        );

    \I__898\ : InMux
    port map (
            O => \N__9515\,
            I => \N__9497\
        );

    \I__897\ : InMux
    port map (
            O => \N__9514\,
            I => \N__9494\
        );

    \I__896\ : InMux
    port map (
            O => \N__9513\,
            I => \N__9491\
        );

    \I__895\ : Span4Mux_v
    port map (
            O => \N__9510\,
            I => \N__9486\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9486\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__9504\,
            I => \N__9483\
        );

    \I__892\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9480\
        );

    \I__891\ : Span12Mux_s9_v
    port map (
            O => \N__9500\,
            I => \N__9473\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__9497\,
            I => \N__9473\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__9494\,
            I => \N__9473\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__9491\,
            I => \N__9470\
        );

    \I__887\ : Span4Mux_v
    port map (
            O => \N__9486\,
            I => \N__9467\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__9483\,
            I => \N__9462\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__9480\,
            I => \N__9462\
        );

    \I__884\ : Span12Mux_v
    port map (
            O => \N__9473\,
            I => \N__9457\
        );

    \I__883\ : Span12Mux_s10_v
    port map (
            O => \N__9470\,
            I => \N__9457\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__9467\,
            I => \N__9452\
        );

    \I__881\ : Span4Mux_v
    port map (
            O => \N__9462\,
            I => \N__9452\
        );

    \I__880\ : Span12Mux_h
    port map (
            O => \N__9457\,
            I => \N__9449\
        );

    \I__879\ : Span4Mux_h
    port map (
            O => \N__9452\,
            I => \N__9446\
        );

    \I__878\ : Odrv12
    port map (
            O => \N__9449\,
            I => \RX_DATA_2\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__9446\,
            I => \RX_DATA_2\
        );

    \I__876\ : InMux
    port map (
            O => \N__9441\,
            I => \bfn_13_12_0_\
        );

    \I__875\ : InMux
    port map (
            O => \N__9438\,
            I => \transmit_module.video_signal_controller.n3191\
        );

    \I__874\ : InMux
    port map (
            O => \N__9435\,
            I => \transmit_module.video_signal_controller.n3192\
        );

    \I__873\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__9429\,
            I => \line_buffer.n3527\
        );

    \I__871\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9423\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__9423\,
            I => \TX_DATA_2\
        );

    \I__869\ : IoInMux
    port map (
            O => \N__9420\,
            I => \N__9416\
        );

    \I__868\ : IoInMux
    port map (
            O => \N__9419\,
            I => \N__9413\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__9416\,
            I => \N__9410\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__9413\,
            I => \N__9407\
        );

    \I__865\ : IoSpan4Mux
    port map (
            O => \N__9410\,
            I => \N__9404\
        );

    \I__864\ : IoSpan4Mux
    port map (
            O => \N__9407\,
            I => \N__9401\
        );

    \I__863\ : Span4Mux_s2_v
    port map (
            O => \N__9404\,
            I => \N__9397\
        );

    \I__862\ : Span4Mux_s2_v
    port map (
            O => \N__9401\,
            I => \N__9394\
        );

    \I__861\ : IoInMux
    port map (
            O => \N__9400\,
            I => \N__9391\
        );

    \I__860\ : Sp12to4
    port map (
            O => \N__9397\,
            I => \N__9388\
        );

    \I__859\ : Sp12to4
    port map (
            O => \N__9394\,
            I => \N__9385\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__9391\,
            I => \N__9382\
        );

    \I__857\ : Span12Mux_s10_v
    port map (
            O => \N__9388\,
            I => \N__9379\
        );

    \I__856\ : Span12Mux_s10_v
    port map (
            O => \N__9385\,
            I => \N__9374\
        );

    \I__855\ : Span12Mux_s9_h
    port map (
            O => \N__9382\,
            I => \N__9374\
        );

    \I__854\ : Odrv12
    port map (
            O => \N__9379\,
            I => n1816
        );

    \I__853\ : Odrv12
    port map (
            O => \N__9374\,
            I => n1816
        );

    \I__852\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9366\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__9366\,
            I => \N__9363\
        );

    \I__850\ : Span12Mux_h
    port map (
            O => \N__9363\,
            I => \N__9360\
        );

    \I__849\ : Odrv12
    port map (
            O => \N__9360\,
            I => \line_buffer.n471\
        );

    \I__848\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9354\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__9354\,
            I => \N__9351\
        );

    \I__846\ : Span4Mux_h
    port map (
            O => \N__9351\,
            I => \N__9348\
        );

    \I__845\ : Odrv4
    port map (
            O => \N__9348\,
            I => \line_buffer.n463\
        );

    \I__844\ : InMux
    port map (
            O => \N__9345\,
            I => \N__9342\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__9342\,
            I => \tvp_video_buffer.BUFFER_1_3\
        );

    \I__842\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9336\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__9336\,
            I => \N__9332\
        );

    \I__840\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9328\
        );

    \I__839\ : Span4Mux_v
    port map (
            O => \N__9332\,
            I => \N__9325\
        );

    \I__838\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9322\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__9328\,
            I => \N__9319\
        );

    \I__836\ : Span4Mux_v
    port map (
            O => \N__9325\,
            I => \N__9313\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__9322\,
            I => \N__9313\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__9319\,
            I => \N__9307\
        );

    \I__833\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9304\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__9313\,
            I => \N__9300\
        );

    \I__831\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9297\
        );

    \I__830\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9294\
        );

    \I__829\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9291\
        );

    \I__828\ : Span4Mux_v
    port map (
            O => \N__9307\,
            I => \N__9286\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__9304\,
            I => \N__9286\
        );

    \I__826\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9283\
        );

    \I__825\ : Sp12to4
    port map (
            O => \N__9300\,
            I => \N__9276\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__9297\,
            I => \N__9276\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__9294\,
            I => \N__9276\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__9291\,
            I => \N__9273\
        );

    \I__821\ : Span4Mux_v
    port map (
            O => \N__9286\,
            I => \N__9270\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__9283\,
            I => \N__9267\
        );

    \I__819\ : Span12Mux_v
    port map (
            O => \N__9276\,
            I => \N__9262\
        );

    \I__818\ : Span12Mux_s9_v
    port map (
            O => \N__9273\,
            I => \N__9262\
        );

    \I__817\ : Span4Mux_v
    port map (
            O => \N__9270\,
            I => \N__9257\
        );

    \I__816\ : Span4Mux_h
    port map (
            O => \N__9267\,
            I => \N__9257\
        );

    \I__815\ : Span12Mux_h
    port map (
            O => \N__9262\,
            I => \N__9254\
        );

    \I__814\ : Span4Mux_h
    port map (
            O => \N__9257\,
            I => \N__9251\
        );

    \I__813\ : Odrv12
    port map (
            O => \N__9254\,
            I => \RX_DATA_1\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__9251\,
            I => \RX_DATA_1\
        );

    \I__811\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__9243\,
            I => \tvp_video_buffer.BUFFER_1_7\
        );

    \I__809\ : IoInMux
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__807\ : IoSpan4Mux
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__806\ : Span4Mux_s2_h
    port map (
            O => \N__9231\,
            I => \N__9227\
        );

    \I__805\ : InMux
    port map (
            O => \N__9230\,
            I => \N__9224\
        );

    \I__804\ : Sp12to4
    port map (
            O => \N__9227\,
            I => \N__9221\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__9224\,
            I => \N__9218\
        );

    \I__802\ : Span12Mux_v
    port map (
            O => \N__9221\,
            I => \N__9215\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__9218\,
            I => \N__9212\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__9215\,
            I => \N__9207\
        );

    \I__799\ : Sp12to4
    port map (
            O => \N__9212\,
            I => \N__9207\
        );

    \I__798\ : Odrv12
    port map (
            O => \N__9207\,
            I => \DEBUG_c_6_c\
        );

    \I__797\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__9201\,
            I => \tvp_video_buffer.BUFFER_0_7\
        );

    \I__795\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9195\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__9195\,
            I => \N__9192\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__9192\,
            I => \tvp_video_buffer.BUFFER_0_4\
        );

    \I__792\ : InMux
    port map (
            O => \N__9189\,
            I => \bfn_12_17_0_\
        );

    \I__791\ : InMux
    port map (
            O => \N__9186\,
            I => \transmit_module.video_signal_controller.n3188\
        );

    \I__790\ : InMux
    port map (
            O => \N__9183\,
            I => \transmit_module.video_signal_controller.n3189\
        );

    \I__789\ : InMux
    port map (
            O => \N__9180\,
            I => \transmit_module.video_signal_controller.n3190\
        );

    \I__788\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9174\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9171\
        );

    \I__786\ : Odrv4
    port map (
            O => \N__9171\,
            I => \transmit_module.Y_DELTA_PATTERN_3\
        );

    \I__785\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9165\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__9165\,
            I => \transmit_module.Y_DELTA_PATTERN_2\
        );

    \I__783\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9159\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__9159\,
            I => \transmit_module.Y_DELTA_PATTERN_1\
        );

    \I__781\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9153\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__779\ : Span4Mux_v
    port map (
            O => \N__9150\,
            I => \N__9147\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__9147\,
            I => \line_buffer.n536\
        );

    \I__777\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9141\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__9141\,
            I => \N__9138\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__9138\,
            I => \N__9135\
        );

    \I__774\ : Sp12to4
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__773\ : Span12Mux_v
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__772\ : Span12Mux_h
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__771\ : Odrv12
    port map (
            O => \N__9126\,
            I => \line_buffer.n528\
        );

    \I__770\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__9117\,
            I => \line_buffer.n3528\
        );

    \I__767\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9111\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__9111\,
            I => \N__9108\
        );

    \I__765\ : Span12Mux_v
    port map (
            O => \N__9108\,
            I => \N__9105\
        );

    \I__764\ : Odrv12
    port map (
            O => \N__9105\,
            I => \line_buffer.n563\
        );

    \I__763\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__9099\,
            I => \N__9096\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__9096\,
            I => \N__9093\
        );

    \I__760\ : Span4Mux_h
    port map (
            O => \N__9093\,
            I => \N__9090\
        );

    \I__759\ : Sp12to4
    port map (
            O => \N__9090\,
            I => \N__9087\
        );

    \I__758\ : Odrv12
    port map (
            O => \N__9087\,
            I => \line_buffer.n555\
        );

    \I__757\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9081\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__9081\,
            I => \N__9078\
        );

    \I__755\ : Span4Mux_v
    port map (
            O => \N__9078\,
            I => \N__9075\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__9075\,
            I => \line_buffer.n3567\
        );

    \I__753\ : InMux
    port map (
            O => \N__9072\,
            I => \bfn_12_16_0_\
        );

    \I__752\ : InMux
    port map (
            O => \N__9069\,
            I => \transmit_module.video_signal_controller.n3180\
        );

    \I__751\ : InMux
    port map (
            O => \N__9066\,
            I => \transmit_module.video_signal_controller.n3181\
        );

    \I__750\ : InMux
    port map (
            O => \N__9063\,
            I => \transmit_module.video_signal_controller.n3182\
        );

    \I__749\ : InMux
    port map (
            O => \N__9060\,
            I => \transmit_module.video_signal_controller.n3183\
        );

    \I__748\ : InMux
    port map (
            O => \N__9057\,
            I => \transmit_module.video_signal_controller.n3184\
        );

    \I__747\ : InMux
    port map (
            O => \N__9054\,
            I => \transmit_module.video_signal_controller.n3185\
        );

    \I__746\ : InMux
    port map (
            O => \N__9051\,
            I => \transmit_module.video_signal_controller.n3186\
        );

    \I__745\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9045\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__9045\,
            I => \transmit_module.Y_DELTA_PATTERN_12\
        );

    \I__743\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9039\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__9039\,
            I => \transmit_module.Y_DELTA_PATTERN_11\
        );

    \I__741\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9033\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__9033\,
            I => \transmit_module.Y_DELTA_PATTERN_10\
        );

    \I__739\ : InMux
    port map (
            O => \N__9030\,
            I => \N__9027\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__9027\,
            I => \sync_buffer.BUFFER_0_0\
        );

    \I__737\ : InMux
    port map (
            O => \N__9024\,
            I => \N__9021\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__9021\,
            I => \sync_buffer.BUFFER_1_0\
        );

    \I__735\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9015\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__9015\,
            I => \RX_TX_SYNC_BUFF\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__9012\,
            I => \transmit_module.video_signal_controller.n3479_cascade_\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__9009\,
            I => \transmit_module.video_signal_controller.n3475_cascade_\
        );

    \I__731\ : InMux
    port map (
            O => \N__9006\,
            I => \N__9003\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__9003\,
            I => \transmit_module.video_signal_controller.n55\
        );

    \I__729\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8997\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__8997\,
            I => \transmit_module.Y_DELTA_PATTERN_63\
        );

    \I__727\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8991\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__8991\,
            I => \transmit_module.Y_DELTA_PATTERN_62\
        );

    \I__725\ : InMux
    port map (
            O => \N__8988\,
            I => \N__8985\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8982\
        );

    \I__723\ : Span12Mux_v
    port map (
            O => \N__8982\,
            I => \N__8979\
        );

    \I__722\ : Odrv12
    port map (
            O => \N__8979\,
            I => \line_buffer.n3569\
        );

    \I__721\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8973\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__8973\,
            I => \line_buffer.n3566\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__8970\,
            I => \line_buffer.n3599_cascade_\
        );

    \I__718\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8964\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__8964\,
            I => \N__8961\
        );

    \I__716\ : Span4Mux_v
    port map (
            O => \N__8961\,
            I => \N__8958\
        );

    \I__715\ : Odrv4
    port map (
            O => \N__8958\,
            I => \line_buffer.n595\
        );

    \I__714\ : InMux
    port map (
            O => \N__8955\,
            I => \N__8952\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__8952\,
            I => \N__8949\
        );

    \I__712\ : Span4Mux_h
    port map (
            O => \N__8949\,
            I => \N__8946\
        );

    \I__711\ : Span4Mux_v
    port map (
            O => \N__8946\,
            I => \N__8943\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__8943\,
            I => \N__8940\
        );

    \I__709\ : Span4Mux_h
    port map (
            O => \N__8940\,
            I => \N__8937\
        );

    \I__708\ : Span4Mux_h
    port map (
            O => \N__8937\,
            I => \N__8934\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__8934\,
            I => \line_buffer.n587\
        );

    \I__706\ : InMux
    port map (
            O => \N__8931\,
            I => \N__8928\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__8928\,
            I => \line_buffer.n3570\
        );

    \I__704\ : InMux
    port map (
            O => \N__8925\,
            I => \N__8922\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__8922\,
            I => \N__8919\
        );

    \I__702\ : Span4Mux_h
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__701\ : IoSpan4Mux
    port map (
            O => \N__8916\,
            I => \N__8913\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__8913\,
            I => \TVP_VIDEO_c_3\
        );

    \I__699\ : InMux
    port map (
            O => \N__8910\,
            I => \N__8907\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__8907\,
            I => \tvp_video_buffer.BUFFER_0_3\
        );

    \I__697\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8901\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__8901\,
            I => \transmit_module.Y_DELTA_PATTERN_71\
        );

    \I__695\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8895\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__8895\,
            I => \transmit_module.Y_DELTA_PATTERN_79\
        );

    \I__693\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8889\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__8889\,
            I => \transmit_module.Y_DELTA_PATTERN_78\
        );

    \I__691\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8883\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__8883\,
            I => \transmit_module.Y_DELTA_PATTERN_72\
        );

    \I__689\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__8877\,
            I => \transmit_module.Y_DELTA_PATTERN_75\
        );

    \I__687\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8871\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__8871\,
            I => \transmit_module.Y_DELTA_PATTERN_53\
        );

    \I__685\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8865\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__8865\,
            I => \transmit_module.Y_DELTA_PATTERN_52\
        );

    \I__683\ : InMux
    port map (
            O => \N__8862\,
            I => \N__8859\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__8859\,
            I => \transmit_module.Y_DELTA_PATTERN_74\
        );

    \I__681\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8853\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__8853\,
            I => \transmit_module.Y_DELTA_PATTERN_73\
        );

    \I__679\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8847\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__8847\,
            I => \transmit_module.Y_DELTA_PATTERN_61\
        );

    \I__677\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8841\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__8841\,
            I => \transmit_module.Y_DELTA_PATTERN_65\
        );

    \I__675\ : InMux
    port map (
            O => \N__8838\,
            I => \N__8835\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__8835\,
            I => \transmit_module.Y_DELTA_PATTERN_64\
        );

    \I__673\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8829\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__8829\,
            I => \transmit_module.Y_DELTA_PATTERN_33\
        );

    \I__671\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8823\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__8823\,
            I => \N__8820\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__8820\,
            I => \transmit_module.Y_DELTA_PATTERN_37\
        );

    \I__668\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8814\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__8814\,
            I => \transmit_module.Y_DELTA_PATTERN_36\
        );

    \I__666\ : InMux
    port map (
            O => \N__8811\,
            I => \N__8808\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__8808\,
            I => \transmit_module.Y_DELTA_PATTERN_35\
        );

    \I__664\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8802\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__8802\,
            I => \transmit_module.Y_DELTA_PATTERN_34\
        );

    \I__662\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8796\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__8796\,
            I => \transmit_module.Y_DELTA_PATTERN_81\
        );

    \I__660\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8790\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__8790\,
            I => \transmit_module.Y_DELTA_PATTERN_82\
        );

    \I__658\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8784\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__8784\,
            I => \transmit_module.Y_DELTA_PATTERN_80\
        );

    \I__656\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__8778\,
            I => \transmit_module.Y_DELTA_PATTERN_51\
        );

    \I__654\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8772\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__8772\,
            I => \transmit_module.Y_DELTA_PATTERN_70\
        );

    \I__652\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8766\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__8766\,
            I => \N__8763\
        );

    \I__650\ : Span4Mux_v
    port map (
            O => \N__8763\,
            I => \N__8760\
        );

    \I__649\ : Sp12to4
    port map (
            O => \N__8760\,
            I => \N__8757\
        );

    \I__648\ : Span12Mux_h
    port map (
            O => \N__8757\,
            I => \N__8754\
        );

    \I__647\ : Odrv12
    port map (
            O => \N__8754\,
            I => \line_buffer.n466\
        );

    \I__646\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8748\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__8748\,
            I => \N__8745\
        );

    \I__644\ : Span4Mux_v
    port map (
            O => \N__8745\,
            I => \N__8742\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__8742\,
            I => \N__8739\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__8736\,
            I => \line_buffer.n458\
        );

    \I__640\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8730\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__8730\,
            I => \N__8727\
        );

    \I__638\ : Span4Mux_v
    port map (
            O => \N__8727\,
            I => \N__8724\
        );

    \I__637\ : Span4Mux_h
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__8721\,
            I => \line_buffer.n531\
        );

    \I__635\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__8715\,
            I => \N__8712\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__8712\,
            I => \N__8709\
        );

    \I__632\ : Span4Mux_h
    port map (
            O => \N__8709\,
            I => \N__8706\
        );

    \I__631\ : Sp12to4
    port map (
            O => \N__8706\,
            I => \N__8703\
        );

    \I__630\ : Odrv12
    port map (
            O => \N__8703\,
            I => \line_buffer.n523\
        );

    \I__629\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8697\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__8697\,
            I => \N__8694\
        );

    \I__627\ : Odrv12
    port map (
            O => \N__8694\,
            I => \TVP_VIDEO_c_4\
        );

    \I__626\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8688\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__8688\,
            I => \transmit_module.Y_DELTA_PATTERN_9\
        );

    \I__624\ : InMux
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__8682\,
            I => \transmit_module.Y_DELTA_PATTERN_29\
        );

    \I__622\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8676\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__8676\,
            I => \transmit_module.Y_DELTA_PATTERN_30\
        );

    \I__620\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8670\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__8670\,
            I => \transmit_module.Y_DELTA_PATTERN_32\
        );

    \I__618\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8664\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__8664\,
            I => \transmit_module.Y_DELTA_PATTERN_31\
        );

    \I__616\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8658\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__8658\,
            I => \transmit_module.Y_DELTA_PATTERN_66\
        );

    \I__614\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8652\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__8652\,
            I => \transmit_module.Y_DELTA_PATTERN_44\
        );

    \I__612\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8646\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__8646\,
            I => \transmit_module.Y_DELTA_PATTERN_43\
        );

    \I__610\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8640\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__8640\,
            I => \transmit_module.Y_DELTA_PATTERN_42\
        );

    \I__608\ : InMux
    port map (
            O => \N__8637\,
            I => \N__8634\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__8634\,
            I => \transmit_module.Y_DELTA_PATTERN_41\
        );

    \I__606\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8628\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__8628\,
            I => \transmit_module.Y_DELTA_PATTERN_40\
        );

    \I__604\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__8622\,
            I => \transmit_module.Y_DELTA_PATTERN_60\
        );

    \I__602\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__8616\,
            I => \N__8613\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__8613\,
            I => \transmit_module.Y_DELTA_PATTERN_7\
        );

    \I__599\ : InMux
    port map (
            O => \N__8610\,
            I => \N__8607\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__8607\,
            I => \N__8604\
        );

    \I__597\ : Odrv4
    port map (
            O => \N__8604\,
            I => \transmit_module.Y_DELTA_PATTERN_6\
        );

    \I__596\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8598\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__8598\,
            I => \transmit_module.Y_DELTA_PATTERN_5\
        );

    \I__594\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8592\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__8592\,
            I => \transmit_module.Y_DELTA_PATTERN_4\
        );

    \I__592\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8586\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__8586\,
            I => \transmit_module.Y_DELTA_PATTERN_50\
        );

    \I__590\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8580\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__8580\,
            I => \transmit_module.Y_DELTA_PATTERN_49\
        );

    \I__588\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__8574\,
            I => \transmit_module.Y_DELTA_PATTERN_54\
        );

    \I__586\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8568\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__8568\,
            I => \transmit_module.Y_DELTA_PATTERN_67\
        );

    \I__584\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8562\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__8562\,
            I => \transmit_module.Y_DELTA_PATTERN_77\
        );

    \I__582\ : InMux
    port map (
            O => \N__8559\,
            I => \N__8556\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__8556\,
            I => \transmit_module.Y_DELTA_PATTERN_69\
        );

    \I__580\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8550\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__8550\,
            I => \transmit_module.Y_DELTA_PATTERN_68\
        );

    \I__578\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__8544\,
            I => \transmit_module.Y_DELTA_PATTERN_76\
        );

    \I__576\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8538\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__8538\,
            I => \N__8535\
        );

    \I__574\ : Span4Mux_v
    port map (
            O => \N__8535\,
            I => \N__8532\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__8532\,
            I => \line_buffer.n600\
        );

    \I__572\ : InMux
    port map (
            O => \N__8529\,
            I => \N__8526\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__8526\,
            I => \N__8523\
        );

    \I__570\ : Span4Mux_v
    port map (
            O => \N__8523\,
            I => \N__8520\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__8520\,
            I => \line_buffer.n592\
        );

    \I__568\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__8514\,
            I => \transmit_module.Y_DELTA_PATTERN_28\
        );

    \I__566\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8508\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__8508\,
            I => \transmit_module.Y_DELTA_PATTERN_27\
        );

    \I__564\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__8502\,
            I => \transmit_module.Y_DELTA_PATTERN_8\
        );

    \I__562\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__8496\,
            I => \transmit_module.Y_DELTA_PATTERN_48\
        );

    \I__560\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__8490\,
            I => \transmit_module.Y_DELTA_PATTERN_47\
        );

    \I__558\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__8484\,
            I => \transmit_module.Y_DELTA_PATTERN_55\
        );

    \I__556\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__8478\,
            I => \transmit_module.Y_DELTA_PATTERN_46\
        );

    \I__554\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__8472\,
            I => \transmit_module.Y_DELTA_PATTERN_58\
        );

    \I__552\ : InMux
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__8466\,
            I => \transmit_module.Y_DELTA_PATTERN_59\
        );

    \I__550\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8460\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__8460\,
            I => \transmit_module.Y_DELTA_PATTERN_57\
        );

    \I__548\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8454\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__8454\,
            I => \transmit_module.Y_DELTA_PATTERN_56\
        );

    \I__546\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8448\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__8448\,
            I => \N__8445\
        );

    \I__544\ : Odrv4
    port map (
            O => \N__8445\,
            I => \transmit_module.Y_DELTA_PATTERN_39\
        );

    \I__543\ : InMux
    port map (
            O => \N__8442\,
            I => \N__8439\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__8439\,
            I => \transmit_module.Y_DELTA_PATTERN_45\
        );

    \I__541\ : InMux
    port map (
            O => \N__8436\,
            I => \N__8433\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__8433\,
            I => \N__8430\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__8430\,
            I => \N__8427\
        );

    \I__538\ : Odrv4
    port map (
            O => \N__8427\,
            I => \line_buffer.n599\
        );

    \I__537\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8421\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__8421\,
            I => \N__8418\
        );

    \I__535\ : Span4Mux_v
    port map (
            O => \N__8418\,
            I => \N__8415\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__8415\,
            I => \line_buffer.n591\
        );

    \I__533\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__8409\,
            I => \transmit_module.Y_DELTA_PATTERN_38\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3198\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3187\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.n3166\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3179\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3214\,
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.n3153\,
            carryinitout => \bfn_15_17_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i26_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8511\,
            lcout => \transmit_module.Y_DELTA_PATTERN_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24301\,
            ce => \N__20514\,
            sr => \N__23331\
        );

    \transmit_module.Y_DELTA_PATTERN_i37_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8412\,
            lcout => \transmit_module.Y_DELTA_PATTERN_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24335\,
            ce => \N__9912\,
            sr => \N__23335\
        );

    \transmit_module.Y_DELTA_PATTERN_i46_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8493\,
            lcout => \transmit_module.Y_DELTA_PATTERN_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24312\,
            ce => \N__9900\,
            sr => \N__23274\
        );

    \transmit_module.Y_DELTA_PATTERN_i38_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8451\,
            lcout => \transmit_module.Y_DELTA_PATTERN_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24312\,
            ce => \N__9900\,
            sr => \N__23274\
        );

    \transmit_module.Y_DELTA_PATTERN_i54_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8487\,
            lcout => \transmit_module.Y_DELTA_PATTERN_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24299\,
            ce => \N__9895\,
            sr => \N__23303\
        );

    \transmit_module.Y_DELTA_PATTERN_i55_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8457\,
            lcout => \transmit_module.Y_DELTA_PATTERN_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24299\,
            ce => \N__9895\,
            sr => \N__23303\
        );

    \transmit_module.Y_DELTA_PATTERN_i45_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8481\,
            lcout => \transmit_module.Y_DELTA_PATTERN_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24299\,
            ce => \N__9895\,
            sr => \N__23303\
        );

    \transmit_module.Y_DELTA_PATTERN_i58_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8469\,
            lcout => \transmit_module.Y_DELTA_PATTERN_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24299\,
            ce => \N__9895\,
            sr => \N__23303\
        );

    \transmit_module.Y_DELTA_PATTERN_i57_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8475\,
            lcout => \transmit_module.Y_DELTA_PATTERN_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24299\,
            ce => \N__9895\,
            sr => \N__23303\
        );

    \transmit_module.Y_DELTA_PATTERN_i59_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8625\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24299\,
            ce => \N__9895\,
            sr => \N__23303\
        );

    \transmit_module.Y_DELTA_PATTERN_i56_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8463\,
            lcout => \transmit_module.Y_DELTA_PATTERN_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24299\,
            ce => \N__9895\,
            sr => \N__23303\
        );

    \transmit_module.Y_DELTA_PATTERN_i39_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8631\,
            lcout => \transmit_module.Y_DELTA_PATTERN_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24241\,
            ce => \N__9913\,
            sr => \N__23300\
        );

    \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8442\,
            lcout => \transmit_module.Y_DELTA_PATTERN_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24241\,
            ce => \N__9913\,
            sr => \N__23300\
        );

    \line_buffer.i2203_3_lut_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22827\,
            in1 => \N__8436\,
            in2 => \_gnd_net_\,
            in3 => \N__8424\,
            lcout => \line_buffer.n3540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2191_3_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22826\,
            in1 => \N__8541\,
            in2 => \_gnd_net_\,
            in3 => \N__8529\,
            lcout => \line_buffer.n3528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i28_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8685\,
            lcout => \transmit_module.Y_DELTA_PATTERN_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24334\,
            ce => \N__20517\,
            sr => \N__23333\
        );

    \transmit_module.Y_DELTA_PATTERN_i27_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8517\,
            lcout => \transmit_module.Y_DELTA_PATTERN_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24352\,
            ce => \N__20499\,
            sr => \N__23332\
        );

    \transmit_module.Y_DELTA_PATTERN_i8_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8691\,
            lcout => \transmit_module.Y_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24352\,
            ce => \N__20499\,
            sr => \N__23332\
        );

    \transmit_module.Y_DELTA_PATTERN_i7_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8505\,
            lcout => \transmit_module.Y_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24352\,
            ce => \N__20499\,
            sr => \N__23332\
        );

    \transmit_module.Y_DELTA_PATTERN_i48_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8583\,
            lcout => \transmit_module.Y_DELTA_PATTERN_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24350\,
            ce => \N__9914\,
            sr => \N__23284\
        );

    \transmit_module.Y_DELTA_PATTERN_i69_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8775\,
            lcout => \transmit_module.Y_DELTA_PATTERN_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24350\,
            ce => \N__9914\,
            sr => \N__23284\
        );

    \transmit_module.Y_DELTA_PATTERN_i47_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8499\,
            lcout => \transmit_module.Y_DELTA_PATTERN_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24350\,
            ce => \N__9914\,
            sr => \N__23284\
        );

    \transmit_module.Y_DELTA_PATTERN_i50_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8781\,
            lcout => \transmit_module.Y_DELTA_PATTERN_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24350\,
            ce => \N__9914\,
            sr => \N__23284\
        );

    \transmit_module.Y_DELTA_PATTERN_i49_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8589\,
            lcout => \transmit_module.Y_DELTA_PATTERN_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24350\,
            ce => \N__9914\,
            sr => \N__23284\
        );

    \transmit_module.Y_DELTA_PATTERN_i53_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8577\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24287\,
            ce => \N__9872\,
            sr => \N__23310\
        );

    \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8565\,
            lcout => \transmit_module.Y_DELTA_PATTERN_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24287\,
            ce => \N__9872\,
            sr => \N__23310\
        );

    \transmit_module.Y_DELTA_PATTERN_i67_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8553\,
            lcout => \transmit_module.Y_DELTA_PATTERN_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24287\,
            ce => \N__9872\,
            sr => \N__23310\
        );

    \transmit_module.Y_DELTA_PATTERN_i66_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8571\,
            lcout => \transmit_module.Y_DELTA_PATTERN_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24287\,
            ce => \N__9872\,
            sr => \N__23310\
        );

    \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8892\,
            lcout => \transmit_module.Y_DELTA_PATTERN_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24287\,
            ce => \N__9872\,
            sr => \N__23310\
        );

    \transmit_module.Y_DELTA_PATTERN_i68_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8559\,
            lcout => \transmit_module.Y_DELTA_PATTERN_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24287\,
            ce => \N__9872\,
            sr => \N__23310\
        );

    \transmit_module.Y_DELTA_PATTERN_i75_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8547\,
            lcout => \transmit_module.Y_DELTA_PATTERN_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24287\,
            ce => \N__9872\,
            sr => \N__23310\
        );

    \transmit_module.Y_DELTA_PATTERN_i41_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8643\,
            lcout => \transmit_module.Y_DELTA_PATTERN_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24292\,
            ce => \N__9908\,
            sr => \N__23228\
        );

    \transmit_module.Y_DELTA_PATTERN_i65_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8661\,
            lcout => \transmit_module.Y_DELTA_PATTERN_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24292\,
            ce => \N__9908\,
            sr => \N__23228\
        );

    \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8655\,
            lcout => \transmit_module.Y_DELTA_PATTERN_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24292\,
            ce => \N__9908\,
            sr => \N__23228\
        );

    \transmit_module.Y_DELTA_PATTERN_i42_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8649\,
            lcout => \transmit_module.Y_DELTA_PATTERN_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24292\,
            ce => \N__9908\,
            sr => \N__23228\
        );

    \transmit_module.Y_DELTA_PATTERN_i40_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8637\,
            lcout => \transmit_module.Y_DELTA_PATTERN_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24292\,
            ce => \N__9908\,
            sr => \N__23228\
        );

    \transmit_module.Y_DELTA_PATTERN_i60_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8850\,
            lcout => \transmit_module.Y_DELTA_PATTERN_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24292\,
            ce => \N__9908\,
            sr => \N__23228\
        );

    \transmit_module.Y_DELTA_PATTERN_i6_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8619\,
            lcout => \transmit_module.Y_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24291\,
            ce => \N__20518\,
            sr => \N__23327\
        );

    \transmit_module.Y_DELTA_PATTERN_i5_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8610\,
            lcout => \transmit_module.Y_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24197\,
            ce => \N__20525\,
            sr => \N__23326\
        );

    \transmit_module.Y_DELTA_PATTERN_i4_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8601\,
            lcout => \transmit_module.Y_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24197\,
            ce => \N__20525\,
            sr => \N__23326\
        );

    \transmit_module.Y_DELTA_PATTERN_i3_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8595\,
            lcout => \transmit_module.Y_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24197\,
            ce => \N__20525\,
            sr => \N__23326\
        );

    \line_buffer.i2229_3_lut_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8769\,
            in1 => \N__8751\,
            in2 => \_gnd_net_\,
            in3 => \N__22831\,
            lcout => \line_buffer.n3566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2232_3_lut_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22828\,
            in1 => \N__8733\,
            in2 => \_gnd_net_\,
            in3 => \N__8718\,
            lcout => \line_buffer.n3569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i3_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8700\,
            lcout => \tvp_video_buffer.BUFFER_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i32_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8832\,
            lcout => \transmit_module.Y_DELTA_PATTERN_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24351\,
            ce => \N__20488\,
            sr => \N__23276\
        );

    \transmit_module.Y_DELTA_PATTERN_i9_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9036\,
            lcout => \transmit_module.Y_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24351\,
            ce => \N__20488\,
            sr => \N__23276\
        );

    \transmit_module.Y_DELTA_PATTERN_i29_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8679\,
            lcout => \transmit_module.Y_DELTA_PATTERN_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24351\,
            ce => \N__20488\,
            sr => \N__23276\
        );

    \transmit_module.Y_DELTA_PATTERN_i30_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8667\,
            lcout => \transmit_module.Y_DELTA_PATTERN_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24351\,
            ce => \N__20488\,
            sr => \N__23276\
        );

    \transmit_module.Y_DELTA_PATTERN_i31_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8673\,
            lcout => \transmit_module.Y_DELTA_PATTERN_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24351\,
            ce => \N__20488\,
            sr => \N__23276\
        );

    \transmit_module.Y_DELTA_PATTERN_i35_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8817\,
            lcout => \transmit_module.Y_DELTA_PATTERN_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24353\,
            ce => \N__9915\,
            sr => \N__23334\
        );

    \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8805\,
            lcout => \transmit_module.Y_DELTA_PATTERN_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24353\,
            ce => \N__9915\,
            sr => \N__23334\
        );

    \transmit_module.Y_DELTA_PATTERN_i36_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8826\,
            lcout => \transmit_module.Y_DELTA_PATTERN_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24353\,
            ce => \N__9915\,
            sr => \N__23334\
        );

    \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8811\,
            lcout => \transmit_module.Y_DELTA_PATTERN_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24353\,
            ce => \N__9915\,
            sr => \N__23334\
        );

    \transmit_module.Y_DELTA_PATTERN_i80_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8799\,
            lcout => \transmit_module.Y_DELTA_PATTERN_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24349\,
            ce => \N__9899\,
            sr => \N__23196\
        );

    \transmit_module.Y_DELTA_PATTERN_i81_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8793\,
            lcout => \transmit_module.Y_DELTA_PATTERN_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24349\,
            ce => \N__9899\,
            sr => \N__23196\
        );

    \transmit_module.Y_DELTA_PATTERN_i82_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21135\,
            lcout => \transmit_module.Y_DELTA_PATTERN_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24349\,
            ce => \N__9899\,
            sr => \N__23196\
        );

    \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8787\,
            lcout => \transmit_module.Y_DELTA_PATTERN_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24349\,
            ce => \N__9899\,
            sr => \N__23196\
        );

    \transmit_module.Y_DELTA_PATTERN_i51_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8868\,
            lcout => \transmit_module.Y_DELTA_PATTERN_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24349\,
            ce => \N__9899\,
            sr => \N__23196\
        );

    \transmit_module.Y_DELTA_PATTERN_i70_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8904\,
            lcout => \transmit_module.Y_DELTA_PATTERN_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24271\,
            ce => \N__9894\,
            sr => \N__23323\
        );

    \transmit_module.Y_DELTA_PATTERN_i71_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8886\,
            lcout => \transmit_module.Y_DELTA_PATTERN_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24271\,
            ce => \N__9894\,
            sr => \N__23323\
        );

    \transmit_module.Y_DELTA_PATTERN_i78_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8898\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24271\,
            ce => \N__9894\,
            sr => \N__23323\
        );

    \transmit_module.Y_DELTA_PATTERN_i72_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8856\,
            lcout => \transmit_module.Y_DELTA_PATTERN_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24271\,
            ce => \N__9894\,
            sr => \N__23323\
        );

    \transmit_module.Y_DELTA_PATTERN_i74_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8880\,
            lcout => \transmit_module.Y_DELTA_PATTERN_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24271\,
            ce => \N__9894\,
            sr => \N__23323\
        );

    \transmit_module.Y_DELTA_PATTERN_i52_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8874\,
            lcout => \transmit_module.Y_DELTA_PATTERN_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24271\,
            ce => \N__9894\,
            sr => \N__23323\
        );

    \transmit_module.Y_DELTA_PATTERN_i73_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8862\,
            lcout => \transmit_module.Y_DELTA_PATTERN_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24271\,
            ce => \N__9894\,
            sr => \N__23323\
        );

    \transmit_module.Y_DELTA_PATTERN_i61_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8994\,
            lcout => \transmit_module.Y_DELTA_PATTERN_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24113\,
            ce => \N__9904\,
            sr => \N__23224\
        );

    \transmit_module.Y_DELTA_PATTERN_i63_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8838\,
            lcout => \transmit_module.Y_DELTA_PATTERN_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24113\,
            ce => \N__9904\,
            sr => \N__23224\
        );

    \transmit_module.Y_DELTA_PATTERN_i64_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8844\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24113\,
            ce => \N__9904\,
            sr => \N__23224\
        );

    \transmit_module.Y_DELTA_PATTERN_i62_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9000\,
            lcout => \transmit_module.Y_DELTA_PATTERN_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24113\,
            ce => \N__9904\,
            sr => \N__23224\
        );

    \transmit_module.ADDR_Y_COMPONENT__i11_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22767\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24222\,
            ce => \N__15388\,
            sr => \N__23324\
        );

    \transmit_module.ADDR_Y_COMPONENT__i10_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12369\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23973\,
            ce => \N__15401\,
            sr => \N__23296\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2266_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__21507\,
            in1 => \N__8931\,
            in2 => \N__21306\,
            in3 => \N__8988\,
            lcout => OPEN,
            ltout => \line_buffer.n3599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i2_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__21304\,
            in1 => \N__8976\,
            in2 => \N__8970\,
            in3 => \N__9084\,
            lcout => \TX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2233_3_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8967\,
            in1 => \N__22829\,
            in2 => \_gnd_net_\,
            in3 => \N__8955\,
            lcout => \line_buffer.n3570\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i2_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8925\,
            lcout => \tvp_video_buffer.BUFFER_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i10_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8910\,
            lcout => \tvp_video_buffer.BUFFER_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21931\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i12_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9567\,
            lcout => \transmit_module.Y_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24332\,
            ce => \N__20510\,
            sr => \N__23275\
        );

    \transmit_module.Y_DELTA_PATTERN_i11_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9048\,
            lcout => \transmit_module.Y_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24332\,
            ce => \N__20510\,
            sr => \N__23275\
        );

    \transmit_module.Y_DELTA_PATTERN_i10_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9042\,
            lcout => \transmit_module.Y_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24332\,
            ce => \N__20510\,
            sr => \N__23275\
        );

    \sync_buffer.BUFFER_0__i1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15540\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sync_buffer.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.WIRE_OUT_0__9_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9024\,
            lcout => \RX_TX_SYNC_BUFF\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.BUFFER_0__i2_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9030\,
            lcout => \sync_buffer.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1160_2_lut_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9018\,
            in2 => \_gnd_net_\,
            in3 => \N__11891\,
            lcout => \transmit_module.video_signal_controller.n2395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__9687\,
            in1 => \N__9939\,
            in2 => \N__9786\,
            in3 => \N__9660\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i3_4_lut_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9735\,
            in1 => \N__9759\,
            in2 => \N__9012\,
            in3 => \N__9815\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101000100"
        )
    port map (
            in0 => \N__12193\,
            in1 => \N__9006\,
            in2 => \N__9009\,
            in3 => \N__9711\,
            lcout => \transmit_module.video_signal_controller.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__9734\,
            in1 => \N__9758\,
            in2 => \N__9816\,
            in3 => \N__9785\,
            lcout => \transmit_module.video_signal_controller.n55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2230_3_lut_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9114\,
            in1 => \N__9102\,
            in2 => \_gnd_net_\,
            in3 => \N__22821\,
            lcout => \line_buffer.n3567\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_X_i0_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9937\,
            in2 => \_gnd_net_\,
            in3 => \N__9072\,
            lcout => \transmit_module.video_signal_controller.VGA_X_0\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \transmit_module.video_signal_controller.n3180\,
            clk => \N__24221\,
            ce => 'H',
            sr => \N__11900\
        );

    \transmit_module.video_signal_controller.VGA_X_i1_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9655\,
            in2 => \_gnd_net_\,
            in3 => \N__9069\,
            lcout => \transmit_module.video_signal_controller.VGA_X_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3180\,
            carryout => \transmit_module.video_signal_controller.n3181\,
            clk => \N__24221\,
            ce => 'H',
            sr => \N__11900\
        );

    \transmit_module.video_signal_controller.VGA_X_i2_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9685\,
            in2 => \_gnd_net_\,
            in3 => \N__9066\,
            lcout => \transmit_module.video_signal_controller.VGA_X_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3181\,
            carryout => \transmit_module.video_signal_controller.n3182\,
            clk => \N__24221\,
            ce => 'H',
            sr => \N__11900\
        );

    \transmit_module.video_signal_controller.VGA_X_i3_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9780\,
            in2 => \_gnd_net_\,
            in3 => \N__9063\,
            lcout => \transmit_module.video_signal_controller.VGA_X_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3182\,
            carryout => \transmit_module.video_signal_controller.n3183\,
            clk => \N__24221\,
            ce => 'H',
            sr => \N__11900\
        );

    \transmit_module.video_signal_controller.VGA_X_i4_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9810\,
            in2 => \_gnd_net_\,
            in3 => \N__9060\,
            lcout => \transmit_module.video_signal_controller.VGA_X_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3183\,
            carryout => \transmit_module.video_signal_controller.n3184\,
            clk => \N__24221\,
            ce => 'H',
            sr => \N__11900\
        );

    \transmit_module.video_signal_controller.VGA_X_i5_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9756\,
            in2 => \_gnd_net_\,
            in3 => \N__9057\,
            lcout => \transmit_module.video_signal_controller.VGA_X_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3184\,
            carryout => \transmit_module.video_signal_controller.n3185\,
            clk => \N__24221\,
            ce => 'H',
            sr => \N__11900\
        );

    \transmit_module.video_signal_controller.VGA_X_i6_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9732\,
            in2 => \_gnd_net_\,
            in3 => \N__9054\,
            lcout => \transmit_module.video_signal_controller.VGA_X_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3185\,
            carryout => \transmit_module.video_signal_controller.n3186\,
            clk => \N__24221\,
            ce => 'H',
            sr => \N__11900\
        );

    \transmit_module.video_signal_controller.VGA_X_i7_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9709\,
            in2 => \_gnd_net_\,
            in3 => \N__9051\,
            lcout => \transmit_module.video_signal_controller.VGA_X_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3186\,
            carryout => \transmit_module.video_signal_controller.n3187\,
            clk => \N__24221\,
            ce => 'H',
            sr => \N__11900\
        );

    \transmit_module.video_signal_controller.VGA_X_i8_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11949\,
            in2 => \_gnd_net_\,
            in3 => \N__9189\,
            lcout => \transmit_module.video_signal_controller.VGA_X_8\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \transmit_module.video_signal_controller.n3188\,
            clk => \N__24067\,
            ce => 'H',
            sr => \N__11904\
        );

    \transmit_module.video_signal_controller.VGA_X_i9_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12150\,
            in2 => \_gnd_net_\,
            in3 => \N__9186\,
            lcout => \transmit_module.video_signal_controller.VGA_X_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3188\,
            carryout => \transmit_module.video_signal_controller.n3189\,
            clk => \N__24067\,
            ce => 'H',
            sr => \N__11904\
        );

    \transmit_module.video_signal_controller.VGA_X_i10_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12189\,
            in2 => \_gnd_net_\,
            in3 => \N__9183\,
            lcout => \transmit_module.video_signal_controller.VGA_X_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3189\,
            carryout => \transmit_module.video_signal_controller.n3190\,
            clk => \N__24067\,
            ce => 'H',
            sr => \N__11904\
        );

    \transmit_module.video_signal_controller.VGA_X_i11_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12242\,
            in2 => \_gnd_net_\,
            in3 => \N__9180\,
            lcout => \transmit_module.video_signal_controller.VGA_X_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24067\,
            ce => 'H',
            sr => \N__11904\
        );

    \transmit_module.Y_DELTA_PATTERN_i0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9162\,
            lcout => \transmit_module.Y_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23978\,
            ce => \N__20526\,
            sr => \N__23336\
        );

    \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9177\,
            lcout => \transmit_module.Y_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23978\,
            ce => \N__20526\,
            sr => \N__23336\
        );

    \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9168\,
            lcout => \transmit_module.Y_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23978\,
            ce => \N__20526\,
            sr => \N__23336\
        );

    \line_buffer.i2190_3_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22808\,
            in1 => \N__9156\,
            in2 => \_gnd_net_\,
            in3 => \N__9144\,
            lcout => \line_buffer.n3527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__21498\,
            in1 => \N__9123\,
            in2 => \N__21300\,
            in3 => \N__9432\,
            lcout => \line_buffer.n3617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i3_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9426\,
            lcout => n1816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23951\,
            ce => 'H',
            sr => \N__22424\
        );

    \line_buffer.i2193_3_lut_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9369\,
            in1 => \N__22830\,
            in2 => \_gnd_net_\,
            in3 => \N__9357\,
            lcout => \line_buffer.n3530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i1_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9345\,
            lcout => \RX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i5_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9246\,
            lcout => \RX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i14_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9204\,
            lcout => \tvp_video_buffer.BUFFER_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i6_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9230\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21932\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i11_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9198\,
            lcout => \tvp_video_buffer.BUFFER_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21951\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i16_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9579\,
            lcout => \transmit_module.Y_DELTA_PATTERN_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24300\,
            ce => \N__20503\,
            sr => \N__23198\
        );

    \transmit_module.Y_DELTA_PATTERN_i17_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9549\,
            lcout => \transmit_module.Y_DELTA_PATTERN_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24300\,
            ce => \N__20503\,
            sr => \N__23198\
        );

    \transmit_module.Y_DELTA_PATTERN_i15_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9573\,
            lcout => \transmit_module.Y_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24300\,
            ce => \N__20503\,
            sr => \N__23198\
        );

    \transmit_module.Y_DELTA_PATTERN_i13_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9555\,
            lcout => \transmit_module.Y_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24300\,
            ce => \N__20503\,
            sr => \N__23198\
        );

    \transmit_module.Y_DELTA_PATTERN_i14_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9561\,
            lcout => \transmit_module.Y_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24300\,
            ce => \N__20503\,
            sr => \N__23198\
        );

    \transmit_module.Y_DELTA_PATTERN_i18_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11451\,
            lcout => \transmit_module.Y_DELTA_PATTERN_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24300\,
            ce => \N__20503\,
            sr => \N__23198\
        );

    \tvp_video_buffer.WIRE_OUT_i2_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9543\,
            lcout => \RX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21959\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11972\,
            in2 => \_gnd_net_\,
            in3 => \N__9441\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_0\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \transmit_module.video_signal_controller.n3191\,
            clk => \N__24283\,
            ce => \N__11899\,
            sr => \N__9597\
        );

    \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11993\,
            in2 => \_gnd_net_\,
            in3 => \N__9438\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3191\,
            carryout => \transmit_module.video_signal_controller.n3192\,
            clk => \N__24283\,
            ce => \N__11899\,
            sr => \N__9597\
        );

    \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12026\,
            in2 => \_gnd_net_\,
            in3 => \N__9435\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3192\,
            carryout => \transmit_module.video_signal_controller.n3193\,
            clk => \N__24283\,
            ce => \N__11899\,
            sr => \N__9597\
        );

    \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11760\,
            in2 => \_gnd_net_\,
            in3 => \N__9624\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3193\,
            carryout => \transmit_module.video_signal_controller.n3194\,
            clk => \N__24283\,
            ce => \N__11899\,
            sr => \N__9597\
        );

    \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11742\,
            in2 => \_gnd_net_\,
            in3 => \N__9621\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3194\,
            carryout => \transmit_module.video_signal_controller.n3195\,
            clk => \N__24283\,
            ce => \N__11899\,
            sr => \N__9597\
        );

    \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11703\,
            in2 => \_gnd_net_\,
            in3 => \N__9618\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3195\,
            carryout => \transmit_module.video_signal_controller.n3196\,
            clk => \N__24283\,
            ce => \N__11899\,
            sr => \N__9597\
        );

    \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11718\,
            in2 => \_gnd_net_\,
            in3 => \N__9615\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3196\,
            carryout => \transmit_module.video_signal_controller.n3197\,
            clk => \N__24283\,
            ce => \N__11899\,
            sr => \N__9597\
        );

    \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11664\,
            in2 => \_gnd_net_\,
            in3 => \N__9612\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3197\,
            carryout => \transmit_module.video_signal_controller.n3198\,
            clk => \N__24283\,
            ce => \N__11899\,
            sr => \N__9597\
        );

    \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11676\,
            in2 => \_gnd_net_\,
            in3 => \N__9609\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_8\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \transmit_module.video_signal_controller.n3199\,
            clk => \N__24228\,
            ce => \N__11898\,
            sr => \N__9593\
        );

    \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13694\,
            in2 => \_gnd_net_\,
            in3 => \N__9606\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3199\,
            carryout => \transmit_module.video_signal_controller.n3200\,
            clk => \N__24228\,
            ce => \N__11898\,
            sr => \N__9593\
        );

    \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13737\,
            in2 => \_gnd_net_\,
            in3 => \N__9603\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3200\,
            carryout => \transmit_module.video_signal_controller.n3201\,
            clk => \N__24228\,
            ce => \N__11898\,
            sr => \N__9593\
        );

    \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13757\,
            in2 => \_gnd_net_\,
            in3 => \N__9600\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24228\,
            ce => \N__11898\,
            sr => \N__9593\
        );

    \transmit_module.video_signal_controller.VGA_HS_66_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12159\,
            in1 => \N__11954\,
            in2 => \N__12256\,
            in3 => \N__9945\,
            lcout => \ADV_HSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1712_2_lut_3_lut_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9686\,
            in1 => \N__9659\,
            in2 => \_gnd_net_\,
            in3 => \N__9938\,
            lcout => \transmit_module.video_signal_controller.n2955\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.old_VGA_HS_40_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.old_VGA_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i124_2_lut_4_lut_rep_24_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__11857\,
            in1 => \N__11787\,
            in2 => \N__23174\,
            in3 => \N__11815\,
            lcout => \transmit_module.n3680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9811\,
            in2 => \_gnd_net_\,
            in3 => \N__9781\,
            lcout => \transmit_module.video_signal_controller.n3363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9757\,
            in1 => \N__9733\,
            in2 => \_gnd_net_\,
            in3 => \N__9710\,
            lcout => \transmit_module.video_signal_controller.n2014\,
            ltout => \transmit_module.video_signal_controller.n2014_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1761_4_lut_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__11953\,
            in1 => \N__9630\,
            in2 => \N__9690\,
            in3 => \N__11927\,
            lcout => \transmit_module.video_signal_controller.n3004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1_3_lut_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__16240\,
            in1 => \N__23120\,
            in2 => \_gnd_net_\,
            in3 => \N__20633\,
            lcout => \transmit_module.n2310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i506_2_lut_rep_20_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9684\,
            in2 => \_gnd_net_\,
            in3 => \N__9654\,
            lcout => \transmit_module.video_signal_controller.n3676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i7_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__16241\,
            in1 => \N__23121\,
            in2 => \N__13005\,
            in3 => \N__13020\,
            lcout => \transmit_module.TX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i1_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__16265\,
            in1 => \N__10683\,
            in2 => \N__23240\,
            in3 => \N__10182\,
            lcout => \transmit_module.TX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i2_3_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12460\,
            in1 => \N__14024\,
            in2 => \_gnd_net_\,
            in3 => \N__12117\,
            lcout => \transmit_module.n146\,
            ltout => \transmit_module.n146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1643_4_lut_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__23119\,
            in1 => \N__16239\,
            in2 => \N__10176\,
            in3 => \N__10682\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i10_3_lut_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20626\,
            in1 => \N__12477\,
            in2 => \_gnd_net_\,
            in3 => \N__12500\,
            lcout => \transmit_module.n107\,
            ltout => \transmit_module.n107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i9_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__10428\,
            in1 => \N__23125\,
            in2 => \N__9951\,
            in3 => \N__16317\,
            lcout => \transmit_module.TX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i3_3_lut_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12106\,
            in1 => \N__14027\,
            in2 => \_gnd_net_\,
            in3 => \N__12084\,
            lcout => \transmit_module.n145\,
            ltout => \transmit_module.n145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i2_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__23253\,
            in1 => \N__16314\,
            in2 => \N__9948\,
            in3 => \N__10956\,
            lcout => \transmit_module.TX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i3_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__16315\,
            in1 => \N__10704\,
            in2 => \N__23241\,
            in3 => \N__10941\,
            lcout => \transmit_module.TX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i5_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__16316\,
            in1 => \N__10674\,
            in2 => \N__23242\,
            in3 => \N__10440\,
            lcout => \transmit_module.TX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i2_3_lut_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12461\,
            in1 => \N__12435\,
            in2 => \_gnd_net_\,
            in3 => \N__20627\,
            lcout => \transmit_module.n115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i6_3_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14029\,
            in2 => \N__12327\,
            in3 => \N__12396\,
            lcout => \transmit_module.n142\,
            ltout => \transmit_module.n142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1647_4_lut_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__23212\,
            in1 => \N__16304\,
            in2 => \N__10668\,
            in3 => \N__10439\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i8_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__16307\,
            in1 => \N__11439\,
            in2 => \N__23299\,
            in3 => \N__11445\,
            lcout => \transmit_module.TX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i6_3_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12397\,
            in1 => \N__20592\,
            in2 => \_gnd_net_\,
            in3 => \N__12375\,
            lcout => \transmit_module.n111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i10_3_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12499\,
            in1 => \N__14028\,
            in2 => \_gnd_net_\,
            in3 => \N__12294\,
            lcout => \transmit_module.n138\,
            ltout => \transmit_module.n138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1651_4_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__23213\,
            in1 => \N__16305\,
            in2 => \N__10422\,
            in3 => \N__10419\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i10_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__16306\,
            in1 => \N__12756\,
            in2 => \N__23298\,
            in3 => \N__12744\,
            lcout => \transmit_module.TX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i9_3_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12427\,
            in1 => \N__20580\,
            in2 => \_gnd_net_\,
            in3 => \N__12405\,
            lcout => \transmit_module.n108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i9_3_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14041\,
            in1 => \N__12426\,
            in2 => \_gnd_net_\,
            in3 => \N__12306\,
            lcout => \transmit_module.n139\,
            ltout => \transmit_module.n139_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1650_4_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__11438\,
            in1 => \N__23234\,
            in2 => \N__11427\,
            in3 => \N__16308\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i11_3_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20579\,
            in1 => \N__11202\,
            in2 => \_gnd_net_\,
            in3 => \N__12362\,
            lcout => \transmit_module.n106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1644_4_lut_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__16322\,
            in1 => \N__10952\,
            in2 => \N__23302\,
            in3 => \N__11190\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i3_3_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20590\,
            in1 => \N__10689\,
            in2 => \_gnd_net_\,
            in3 => \N__12107\,
            lcout => \transmit_module.n114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i4_3_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12075\,
            in1 => \N__14042\,
            in2 => \_gnd_net_\,
            in3 => \N__12048\,
            lcout => \transmit_module.n144\,
            ltout => \transmit_module.n144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1645_4_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__23286\,
            in1 => \N__16323\,
            in2 => \N__10932\,
            in3 => \N__10700\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i4_3_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20591\,
            in1 => \N__11586\,
            in2 => \_gnd_net_\,
            in3 => \N__12073\,
            lcout => \transmit_module.n113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i2_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12108\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23852\,
            ce => \N__15390\,
            sr => \N__23238\
        );

    \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12074\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23852\,
            ce => \N__15390\,
            sr => \N__23238\
        );

    \line_buffer.i2194_3_lut_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11580\,
            in1 => \N__11565\,
            in2 => \_gnd_net_\,
            in3 => \N__22832\,
            lcout => OPEN,
            ltout => \line_buffer.n3531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i7_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__21294\,
            in1 => \N__11547\,
            in2 => \N__11535\,
            in3 => \N__11532\,
            lcout => \TX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i8_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11526\,
            lcout => \ADV_B_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23835\,
            ce => 'H',
            sr => \N__22414\
        );

    \transmit_module.X_DELTA_PATTERN_i6_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13866\,
            lcout => \transmit_module.X_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24333\,
            ce => \N__18663\,
            sr => \N__20492\
        );

    \transmit_module.X_DELTA_PATTERN_i12_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11622\,
            lcout => \transmit_module.X_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24333\,
            ce => \N__18663\,
            sr => \N__20492\
        );

    \transmit_module.Y_DELTA_PATTERN_i24_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11457\,
            lcout => \transmit_module.Y_DELTA_PATTERN_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24331\,
            ce => \N__20487\,
            sr => \N__23197\
        );

    \transmit_module.Y_DELTA_PATTERN_i25_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11469\,
            lcout => \transmit_module.Y_DELTA_PATTERN_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24331\,
            ce => \N__20487\,
            sr => \N__23197\
        );

    \transmit_module.Y_DELTA_PATTERN_i19_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11652\,
            lcout => \transmit_module.Y_DELTA_PATTERN_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24331\,
            ce => \N__20487\,
            sr => \N__23197\
        );

    \transmit_module.Y_DELTA_PATTERN_i20_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11646\,
            lcout => \transmit_module.Y_DELTA_PATTERN_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24331\,
            ce => \N__20487\,
            sr => \N__23197\
        );

    \transmit_module.Y_DELTA_PATTERN_i21_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11640\,
            lcout => \transmit_module.Y_DELTA_PATTERN_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24331\,
            ce => \N__20487\,
            sr => \N__23197\
        );

    \transmit_module.Y_DELTA_PATTERN_i22_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11628\,
            lcout => \transmit_module.Y_DELTA_PATTERN_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24331\,
            ce => \N__20487\,
            sr => \N__23197\
        );

    \transmit_module.Y_DELTA_PATTERN_i23_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11634\,
            lcout => \transmit_module.Y_DELTA_PATTERN_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24331\,
            ce => \N__20487\,
            sr => \N__23197\
        );

    \transmit_module.X_DELTA_PATTERN_i13_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11613\,
            lcout => \transmit_module.X_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24273\,
            ce => \N__18655\,
            sr => \N__20486\
        );

    \transmit_module.X_DELTA_PATTERN_i14_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18675\,
            lcout => \transmit_module.X_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24273\,
            ce => \N__18655\,
            sr => \N__20486\
        );

    \transmit_module.X_DELTA_PATTERN_i3_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11592\,
            lcout => \transmit_module.X_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24273\,
            ce => \N__18655\,
            sr => \N__20486\
        );

    \transmit_module.X_DELTA_PATTERN_i5_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11607\,
            lcout => \transmit_module.X_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24273\,
            ce => \N__18655\,
            sr => \N__20486\
        );

    \transmit_module.X_DELTA_PATTERN_i4_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24273\,
            ce => \N__18655\,
            sr => \N__20486\
        );

    \transmit_module.video_signal_controller.i480_2_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11992\,
            in2 => \_gnd_net_\,
            in3 => \N__12025\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n6_adj_622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__11739\,
            in1 => \N__11758\,
            in2 => \N__11763\,
            in3 => \N__11684\,
            lcout => \transmit_module.video_signal_controller.VGA_VISIBLE_N_588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2180_3_lut_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__11740\,
            in1 => \N__11759\,
            in2 => \_gnd_net_\,
            in3 => \N__11685\,
            lcout => \transmit_module.video_signal_controller.n3517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11757\,
            in1 => \N__11991\,
            in2 => \_gnd_net_\,
            in3 => \N__12024\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__11717\,
            in1 => \N__11741\,
            in2 => \N__11721\,
            in3 => \N__11702\,
            lcout => \transmit_module.video_signal_controller.n3461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13753\,
            in1 => \N__13729\,
            in2 => \_gnd_net_\,
            in3 => \N__11716\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i4_4_lut_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13690\,
            in1 => \N__11701\,
            in2 => \N__11688\,
            in3 => \N__13709\,
            lcout => \transmit_module.video_signal_controller.n2016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12272\,
            in2 => \_gnd_net_\,
            in3 => \N__13673\,
            lcout => \transmit_module.VGA_VISIBLE_Y\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11675\,
            in2 => \_gnd_net_\,
            in3 => \N__11663\,
            lcout => \transmit_module.video_signal_controller.n3375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i124_2_lut_4_lut_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__11786\,
            in1 => \N__23025\,
            in2 => \N__11859\,
            in3 => \N__11814\,
            lcout => \transmit_module.n2206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VS_67_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__12033\,
            in1 => \N__12006\,
            in2 => \N__12000\,
            in3 => \N__11973\,
            lcout => \ADV_VSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i124_2_lut_4_lut_rep_23_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__11785\,
            in1 => \N__23024\,
            in2 => \N__11858\,
            in3 => \N__11813\,
            lcout => \transmit_module.n3679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1729_4_lut_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__11961\,
            in1 => \N__11955\,
            in2 => \N__11928\,
            in3 => \N__11913\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2972_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1735_4_lut_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__12255\,
            in1 => \N__12199\,
            in2 => \N__11907\,
            in3 => \N__12162\,
            lcout => \transmit_module.video_signal_controller.n2047\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i1_3_lut_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20628\,
            in1 => \N__12471\,
            in2 => \_gnd_net_\,
            in3 => \N__13909\,
            lcout => \transmit_module.n116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i2_3_lut_rep_19_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11850\,
            in1 => \N__11812\,
            in2 => \_gnd_net_\,
            in3 => \N__11784\,
            lcout => \transmit_module.n3675\,
            ltout => \transmit_module.n3675_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i2_3_lut_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__23091\,
            in1 => \_gnd_net_\,
            in2 => \N__11766\,
            in3 => \N__14026\,
            lcout => \transmit_module.n2084\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_2_lut_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12257\,
            in2 => \_gnd_net_\,
            in3 => \N__12160\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n6_adj_623_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__12201\,
            in1 => \N__12210\,
            in2 => \N__12276\,
            in3 => \N__12273\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n7_adj_624_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__12258\,
            in1 => \N__13674\,
            in2 => \N__12213\,
            in3 => \N__12123\,
            lcout => \transmit_module.VGA_VISIBLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1696_4_lut_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110100"
        )
    port map (
            in0 => \N__20629\,
            in1 => \N__16264\,
            in2 => \N__23223\,
            in3 => \N__14025\,
            lcout => \transmit_module.n2070\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1771_3_lut_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__12209\,
            in1 => \N__12200\,
            in2 => \_gnd_net_\,
            in3 => \N__12161\,
            lcout => \transmit_module.video_signal_controller.n3014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_2_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18686\,
            in2 => \N__13913\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n132\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \transmit_module.n3159\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_3_lut_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12453\,
            in2 => \_gnd_net_\,
            in3 => \N__12111\,
            lcout => \transmit_module.n131\,
            ltout => OPEN,
            carryin => \transmit_module.n3159\,
            carryout => \transmit_module.n3160\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_4_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12100\,
            in2 => \_gnd_net_\,
            in3 => \N__12078\,
            lcout => \transmit_module.n130\,
            ltout => OPEN,
            carryin => \transmit_module.n3160\,
            carryout => \transmit_module.n3161\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_5_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12064\,
            in2 => \_gnd_net_\,
            in3 => \N__12036\,
            lcout => \transmit_module.n129\,
            ltout => OPEN,
            carryin => \transmit_module.n3161\,
            carryout => \transmit_module.n3162\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_6_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15513\,
            in2 => \_gnd_net_\,
            in3 => \N__12330\,
            lcout => \transmit_module.n128\,
            ltout => OPEN,
            carryin => \transmit_module.n3162\,
            carryout => \transmit_module.n3163\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_7_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12399\,
            in3 => \N__12315\,
            lcout => \transmit_module.n127\,
            ltout => OPEN,
            carryin => \transmit_module.n3163\,
            carryout => \transmit_module.n3164\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_8_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15439\,
            in3 => \N__12312\,
            lcout => \transmit_module.n126\,
            ltout => OPEN,
            carryin => \transmit_module.n3164\,
            carryout => \transmit_module.n3165\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_9_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15477\,
            in3 => \N__12309\,
            lcout => \transmit_module.n125\,
            ltout => OPEN,
            carryin => \transmit_module.n3165\,
            carryout => \transmit_module.n3166\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_10_lut_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12429\,
            in3 => \N__12297\,
            lcout => \transmit_module.n124\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \transmit_module.n3167\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_11_lut_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12501\,
            in3 => \N__12288\,
            lcout => \transmit_module.n123\,
            ltout => OPEN,
            carryin => \transmit_module.n3167\,
            carryout => \transmit_module.n3168\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_12_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12360\,
            in2 => \_gnd_net_\,
            in3 => \N__12285\,
            lcout => \transmit_module.n122\,
            ltout => OPEN,
            carryin => \transmit_module.n3168\,
            carryout => \transmit_module.n3169\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_13_lut_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22763\,
            in2 => \_gnd_net_\,
            in3 => \N__12282\,
            lcout => \transmit_module.n121\,
            ltout => OPEN,
            carryin => \transmit_module.n3169\,
            carryout => \transmit_module.n3170\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_14_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21439\,
            in2 => \_gnd_net_\,
            in3 => \N__12279\,
            lcout => \transmit_module.n120\,
            ltout => OPEN,
            carryin => \transmit_module.n3170\,
            carryout => \transmit_module.n3171\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_15_lut_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21228\,
            in2 => \_gnd_net_\,
            in3 => \N__12504\,
            lcout => \transmit_module.n119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i9_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12498\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24146\,
            ce => \N__15397\,
            sr => \N__23140\
        );

    \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13914\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24066\,
            ce => \N__15389\,
            sr => \N__23239\
        );

    \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12462\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24066\,
            ce => \N__15389\,
            sr => \N__23239\
        );

    \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12428\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24066\,
            ce => \N__15389\,
            sr => \N__23239\
        );

    \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21484\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24066\,
            ce => \N__15389\,
            sr => \N__23239\
        );

    \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21270\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24066\,
            ce => \N__15389\,
            sr => \N__23239\
        );

    \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12398\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24066\,
            ce => \N__15389\,
            sr => \N__23239\
        );

    \transmit_module.mux_14_i11_3_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14039\,
            in1 => \N__12361\,
            in2 => \_gnd_net_\,
            in3 => \N__12339\,
            lcout => \transmit_module.n137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i7_3_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20604\,
            in1 => \N__15408\,
            in2 => \_gnd_net_\,
            in3 => \N__15444\,
            lcout => \transmit_module.n110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i8_3_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20605\,
            in1 => \N__15450\,
            in2 => \_gnd_net_\,
            in3 => \N__15488\,
            lcout => \transmit_module.n109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1648_4_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__16299\,
            in1 => \N__13778\,
            in2 => \N__23297\,
            in3 => \N__13797\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i5_3_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20625\,
            in1 => \N__15495\,
            in2 => \_gnd_net_\,
            in3 => \N__15525\,
            lcout => \transmit_module.n112\,
            ltout => \transmit_module.n112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1646_4_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__16298\,
            in1 => \N__23233\,
            in2 => \N__13242\,
            in3 => \N__13956\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i8_3_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14040\,
            in1 => \N__15487\,
            in2 => \_gnd_net_\,
            in3 => \N__13029\,
            lcout => \transmit_module.n140\,
            ltout => \transmit_module.n140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1649_4_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__16300\,
            in1 => \N__23229\,
            in2 => \N__13008\,
            in3 => \N__12995\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1652_4_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__16321\,
            in1 => \N__12755\,
            in2 => \N__23301\,
            in3 => \N__12743\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1141_1_lut_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14043\,
            lcout => \transmit_module.n2385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i4_LC_15_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_vs_buffer.BUFFER_0__i1_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13610\,
            lcout => \tvp_vs_buffer.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21933\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_vs_buffer.BUFFER_0__i2_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13593\,
            lcout => \tvp_vs_buffer.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21933\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_vs_buffer.BUFFER_0__i3_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13587\,
            lcout => \tvp_vs_buffer.BUFFER_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.sync_wd.i2_2_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19873\,
            in2 => \_gnd_net_\,
            in3 => \N__21007\,
            lcout => OPEN,
            ltout => \receive_module.sync_wd.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.sync_wd.i1_4_lut_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__21692\,
            in1 => \N__13549\,
            in2 => \N__13476\,
            in3 => \N__19668\,
            lcout => OPEN,
            ltout => \receive_module.sync_wd.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.sync_wd.SYNC_BAD_16_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__13470\,
            in1 => \N__18163\,
            in2 => \N__13473\,
            in3 => \N__20096\,
            lcout => \DEBUG_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.sync_wd.old_visible_17_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19669\,
            lcout => \receive_module.sync_wd.old_visible\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.X_243__i0_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15705\,
            in2 => \_gnd_net_\,
            in3 => \N__13464\,
            lcout => \receive_module.rx_counter.X_0\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \receive_module.rx_counter.n3207\,
            clk => \N__21947\,
            ce => 'H',
            sr => \N__15746\
        );

    \receive_module.rx_counter.X_243__i1_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15729\,
            in2 => \_gnd_net_\,
            in3 => \N__13662\,
            lcout => \receive_module.rx_counter.X_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3207\,
            carryout => \receive_module.rx_counter.n3208\,
            clk => \N__21947\,
            ce => 'H',
            sr => \N__15746\
        );

    \receive_module.rx_counter.X_243__i2_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15717\,
            in2 => \_gnd_net_\,
            in3 => \N__13659\,
            lcout => \receive_module.rx_counter.X_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3208\,
            carryout => \receive_module.rx_counter.n3209\,
            clk => \N__21947\,
            ce => 'H',
            sr => \N__15746\
        );

    \receive_module.rx_counter.X_243__i3_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16003\,
            in2 => \_gnd_net_\,
            in3 => \N__13656\,
            lcout => \receive_module.rx_counter.X_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3209\,
            carryout => \receive_module.rx_counter.n3210\,
            clk => \N__21947\,
            ce => 'H',
            sr => \N__15746\
        );

    \receive_module.rx_counter.X_243__i4_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15946\,
            in2 => \_gnd_net_\,
            in3 => \N__13653\,
            lcout => \receive_module.rx_counter.X_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3210\,
            carryout => \receive_module.rx_counter.n3211\,
            clk => \N__21947\,
            ce => 'H',
            sr => \N__15746\
        );

    \receive_module.rx_counter.X_243__i5_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15976\,
            in2 => \_gnd_net_\,
            in3 => \N__13650\,
            lcout => \receive_module.rx_counter.X_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3211\,
            carryout => \receive_module.rx_counter.n3212\,
            clk => \N__21947\,
            ce => 'H',
            sr => \N__15746\
        );

    \receive_module.rx_counter.X_243__i6_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15871\,
            in2 => \_gnd_net_\,
            in3 => \N__13647\,
            lcout => \receive_module.rx_counter.X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3212\,
            carryout => \receive_module.rx_counter.n3213\,
            clk => \N__21947\,
            ce => 'H',
            sr => \N__15746\
        );

    \receive_module.rx_counter.X_243__i7_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15901\,
            in2 => \_gnd_net_\,
            in3 => \N__13644\,
            lcout => \receive_module.rx_counter.X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3213\,
            carryout => \receive_module.rx_counter.n3214\,
            clk => \N__21947\,
            ce => 'H',
            sr => \N__15746\
        );

    \receive_module.rx_counter.X_243__i8_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15842\,
            in2 => \_gnd_net_\,
            in3 => \N__13641\,
            lcout => \receive_module.rx_counter.X_8\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \receive_module.rx_counter.n3215\,
            clk => \N__21952\,
            ce => 'H',
            sr => \N__15750\
        );

    \receive_module.rx_counter.X_243__i9_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15824\,
            in2 => \_gnd_net_\,
            in3 => \N__13638\,
            lcout => \receive_module.rx_counter.X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21952\,
            ce => 'H',
            sr => \N__15750\
        );

    \receive_module.rx_counter.old_VS_52_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20067\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.rx_counter.old_VS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21955\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_adj_25_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16004\,
            in2 => \_gnd_net_\,
            in3 => \N__15977\,
            lcout => \receive_module.rx_counter.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i131_2_lut_rep_16_2_lut_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18998\,
            in2 => \_gnd_net_\,
            in3 => \N__20066\,
            lcout => \receive_module.rx_counter.n3672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13767\,
            lcout => \TVP_VSYNC_buff\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21955\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_24_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15950\,
            in2 => \_gnd_net_\,
            in3 => \N__15872\,
            lcout => \receive_module.rx_counter.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20056\,
            lcout => \receive_module.n3674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13758\,
            in2 => \_gnd_net_\,
            in3 => \N__13736\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3673_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__13716\,
            in1 => \N__13710\,
            in2 => \N__13698\,
            in3 => \N__13695\,
            lcout => \transmit_module.video_signal_controller.n3379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13809\,
            lcout => \transmit_module.X_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24250\,
            ce => \N__18645\,
            sr => \N__20419\
        );

    \transmit_module.X_DELTA_PATTERN_i8_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13845\,
            lcout => \transmit_module.X_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24250\,
            ce => \N__18645\,
            sr => \N__20419\
        );

    \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13872\,
            lcout => \transmit_module.X_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24250\,
            ce => \N__18645\,
            sr => \N__20419\
        );

    \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13854\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24250\,
            ce => \N__18645\,
            sr => \N__20419\
        );

    \transmit_module.X_DELTA_PATTERN_i9_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13839\,
            lcout => \transmit_module.X_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24250\,
            ce => \N__18645\,
            sr => \N__20419\
        );

    \transmit_module.X_DELTA_PATTERN_i10_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13821\,
            lcout => \transmit_module.X_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24250\,
            ce => \N__18645\,
            sr => \N__20419\
        );

    \transmit_module.X_DELTA_PATTERN_i11_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13833\,
            lcout => \transmit_module.X_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24250\,
            ce => \N__18645\,
            sr => \N__20419\
        );

    \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13815\,
            lcout => \transmit_module.X_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24250\,
            ce => \N__18645\,
            sr => \N__20419\
        );

    \transmit_module.mux_14_i7_3_lut_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14001\,
            in1 => \N__15432\,
            in2 => \_gnd_net_\,
            in3 => \N__13803\,
            lcout => \transmit_module.n141\,
            ltout => \transmit_module.n141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i6_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__23143\,
            in1 => \N__16238\,
            in2 => \N__13785\,
            in3 => \N__13782\,
            lcout => \transmit_module.TX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i1_3_lut_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14002\,
            in1 => \N__14274\,
            in2 => \_gnd_net_\,
            in3 => \N__13908\,
            lcout => \transmit_module.n147\,
            ltout => \transmit_module.n147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1637_4_lut_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__23141\,
            in1 => \N__16233\,
            in2 => \N__14268\,
            in3 => \N__13928\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i5_3_lut_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14000\,
            in1 => \N__15514\,
            in2 => \_gnd_net_\,
            in3 => \N__13962\,
            lcout => \transmit_module.n143\,
            ltout => \transmit_module.n143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i4_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__23142\,
            in1 => \N__13944\,
            in2 => \N__13932\,
            in3 => \N__16237\,
            lcout => \transmit_module.TX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i0_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__13929\,
            in1 => \N__23144\,
            in2 => \N__16266\,
            in3 => \N__13920\,
            lcout => \transmit_module.TX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_2_lut_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14637\,
            in2 => \_gnd_net_\,
            in3 => \N__13884\,
            lcout => \receive_module.n137\,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \receive_module.n3146\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_3_lut_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15123\,
            in2 => \_gnd_net_\,
            in3 => \N__13881\,
            lcout => \receive_module.n136\,
            ltout => OPEN,
            carryin => \receive_module.n3146\,
            carryout => \receive_module.n3147\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_4_lut_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14356\,
            in2 => \_gnd_net_\,
            in3 => \N__13878\,
            lcout => \receive_module.n135\,
            ltout => OPEN,
            carryin => \receive_module.n3147\,
            carryout => \receive_module.n3148\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_5_lut_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17617\,
            in2 => \_gnd_net_\,
            in3 => \N__13875\,
            lcout => \receive_module.n134\,
            ltout => OPEN,
            carryin => \receive_module.n3148\,
            carryout => \receive_module.n3149\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_6_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17362\,
            in3 => \N__14301\,
            lcout => \receive_module.n133\,
            ltout => OPEN,
            carryin => \receive_module.n3149\,
            carryout => \receive_module.n3150\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_7_lut_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19348\,
            in2 => \_gnd_net_\,
            in3 => \N__14298\,
            lcout => \receive_module.n132\,
            ltout => OPEN,
            carryin => \receive_module.n3150\,
            carryout => \receive_module.n3151\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_8_lut_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16864\,
            in2 => \_gnd_net_\,
            in3 => \N__14295\,
            lcout => \receive_module.n131\,
            ltout => OPEN,
            carryin => \receive_module.n3151\,
            carryout => \receive_module.n3152\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_9_lut_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16618\,
            in2 => \_gnd_net_\,
            in3 => \N__14292\,
            lcout => \receive_module.n130\,
            ltout => OPEN,
            carryin => \receive_module.n3152\,
            carryout => \receive_module.n3153\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_10_lut_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17116\,
            in2 => \_gnd_net_\,
            in3 => \N__14289\,
            lcout => \receive_module.n129\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \receive_module.n3154\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_11_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17853\,
            in2 => \_gnd_net_\,
            in3 => \N__14286\,
            lcout => \receive_module.n128\,
            ltout => OPEN,
            carryin => \receive_module.n3154\,
            carryout => \receive_module.n3155\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_12_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14880\,
            in2 => \_gnd_net_\,
            in3 => \N__14283\,
            lcout => \receive_module.n127\,
            ltout => OPEN,
            carryin => \receive_module.n3155\,
            carryout => \receive_module.n3156\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i11_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18762\,
            in2 => \_gnd_net_\,
            in3 => \N__14280\,
            lcout => \RX_ADDR_11\,
            ltout => OPEN,
            carryin => \receive_module.n3156\,
            carryout => \receive_module.n3157\,
            clk => \N__21966\,
            ce => \N__16164\,
            sr => \N__19272\
        );

    \receive_module.BRAM_ADDR__i12_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18919\,
            in2 => \_gnd_net_\,
            in3 => \N__14277\,
            lcout => \RX_ADDR_12\,
            ltout => OPEN,
            carryin => \receive_module.n3157\,
            carryout => \receive_module.n3158\,
            clk => \N__21966\,
            ce => \N__16164\,
            sr => \N__19272\
        );

    \receive_module.BRAM_ADDR__i13_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18834\,
            in2 => \_gnd_net_\,
            in3 => \N__15528\,
            lcout => \RX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21966\,
            ce => \N__16164\,
            sr => \N__19272\
        );

    \transmit_module.ADDR_Y_COMPONENT__i4_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15524\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23977\,
            ce => \N__15402\,
            sr => \N__23252\
        );

    \transmit_module.ADDR_Y_COMPONENT__i7_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15489\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23977\,
            ce => \N__15402\,
            sr => \N__23252\
        );

    \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15443\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23977\,
            ce => \N__15402\,
            sr => \N__23252\
        );

    \receive_module.BRAM_ADDR__i1_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__20132\,
            in1 => \N__15327\,
            in2 => \N__15124\,
            in3 => \N__19672\,
            lcout => \RX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21971\,
            ce => 'H',
            sr => \N__19291\
        );

    \receive_module.BRAM_ADDR__i10_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__19671\,
            in1 => \N__20131\,
            in2 => \N__14881\,
            in3 => \N__15090\,
            lcout => \RX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21971\,
            ce => 'H',
            sr => \N__19291\
        );

    \receive_module.BRAM_ADDR__i0_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__20130\,
            in1 => \N__14844\,
            in2 => \N__14638\,
            in3 => \N__19670\,
            lcout => \RX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21971\,
            ce => 'H',
            sr => \N__19291\
        );

    \transmit_module.VGA_R__i1_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20919\,
            lcout => n1818,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23845\,
            ce => 'H',
            sr => \N__22397\
        );

    \receive_module.BRAM_ADDR__i2_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__20139\,
            in1 => \N__14553\,
            in2 => \N__19697\,
            in3 => \N__14328\,
            lcout => \RX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__19302\
        );

    \tvp_video_buffer.BUFFER_0__i12_LC_16_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15681\,
            lcout => \tvp_video_buffer.BUFFER_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21927\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__18621\,
            in1 => \N__18544\,
            in2 => \N__18600\,
            in3 => \N__18570\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_4_lut_adj_22_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__18521\,
            in1 => \N__18461\,
            in2 => \N__15672\,
            in3 => \N__15761\,
            lcout => \receive_module.rx_counter.n4_adj_612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__18520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18460\,
            lcout => \receive_module.rx_counter.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i3_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15669\,
            lcout => \RX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_27_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18519\,
            in2 => \_gnd_net_\,
            in3 => \N__18543\,
            lcout => \receive_module.rx_counter.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__18594\,
            in1 => \N__18622\,
            in2 => \_gnd_net_\,
            in3 => \N__18571\,
            lcout => \receive_module.rx_counter.n3450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i6_4_lut_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__18572\,
            in1 => \N__18595\,
            in2 => \N__18549\,
            in3 => \N__19179\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.SYNC_46_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15552\,
            in1 => \N__18623\,
            in2 => \N__15543\,
            in3 => \N__15762\,
            lcout => \RX_TX_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_3_lut_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__18500\,
            in1 => \N__18459\,
            in2 => \_gnd_net_\,
            in3 => \N__18482\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_adj_21_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__19180\,
            in1 => \N__15780\,
            in2 => \N__15771\,
            in3 => \N__15768\,
            lcout => \receive_module.rx_counter.n3478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i606_2_lut_rep_21_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18481\,
            in2 => \_gnd_net_\,
            in3 => \N__18499\,
            lcout => \receive_module.rx_counter.n3677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_1_lut_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20001\,
            lcout => \receive_module.rx_counter.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_adj_23_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15728\,
            in1 => \N__15716\,
            in2 => \_gnd_net_\,
            in3 => \N__15704\,
            lcout => \receive_module.rx_counter.n3222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19032\,
            in2 => \_gnd_net_\,
            in3 => \N__15693\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_0\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \receive_module.rx_counter.n3202\,
            clk => \N__21953\,
            ce => \N__18947\,
            sr => \N__18981\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16020\,
            in2 => \_gnd_net_\,
            in3 => \N__15690\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3202\,
            carryout => \receive_module.rx_counter.n3203\,
            clk => \N__21953\,
            ce => \N__18947\,
            sr => \N__18981\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19044\,
            in2 => \_gnd_net_\,
            in3 => \N__15687\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3203\,
            carryout => \receive_module.rx_counter.n3204\,
            clk => \N__21953\,
            ce => \N__18947\,
            sr => \N__18981\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19020\,
            in2 => \_gnd_net_\,
            in3 => \N__15684\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3204\,
            carryout => \receive_module.rx_counter.n3205\,
            clk => \N__21953\,
            ce => \N__18947\,
            sr => \N__18981\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19056\,
            in2 => \_gnd_net_\,
            in3 => \N__16050\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3205\,
            carryout => \receive_module.rx_counter.n3206\,
            clk => \N__21953\,
            ce => \N__18947\,
            sr => \N__18981\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16032\,
            in2 => \_gnd_net_\,
            in3 => \N__16047\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21953\,
            ce => \N__18947\,
            sr => \N__18981\
        );

    \receive_module.rx_counter.i2089_4_lut_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__16044\,
            in1 => \N__16038\,
            in2 => \N__15909\,
            in3 => \N__15924\,
            lcout => \receive_module.rx_counter.n3426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2182_2_lut_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16031\,
            in2 => \_gnd_net_\,
            in3 => \N__16019\,
            lcout => \receive_module.rx_counter.n3519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16008\,
            in1 => \N__15981\,
            in2 => \N__15954\,
            in3 => \N__15923\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_4_lut_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__15908\,
            in1 => \N__15848\,
            in2 => \N__15879\,
            in3 => \N__15876\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i58_4_lut_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__15849\,
            in1 => \N__15828\,
            in2 => \N__15810\,
            in3 => \N__15807\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.O_VISIBLE_53_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__19191\,
            in1 => \N__15801\,
            in2 => \N__15792\,
            in3 => \N__15789\,
            lcout => \DEBUG_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21960\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__18920\,
            in1 => \N__19592\,
            in2 => \N__18866\,
            in3 => \N__18779\,
            lcout => \line_buffer.n473\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__18921\,
            in1 => \N__19591\,
            in2 => \N__18867\,
            in3 => \N__18780\,
            lcout => \line_buffer.n570\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__18781\,
            in1 => \N__18922\,
            in2 => \N__18871\,
            in3 => \N__19593\,
            lcout => \line_buffer.n571\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__rep_1_i0_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16377\,
            in1 => \N__16320\,
            in2 => \_gnd_net_\,
            in3 => \N__16365\,
            lcout => \TX_ADDR_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24102\,
            ce => \N__16179\,
            sr => \N__23243\
        );

    \transmit_module.BRAM_ADDR__i13_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16319\,
            in1 => \N__16356\,
            in2 => \_gnd_net_\,
            in3 => \N__16344\,
            lcout => \TX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24102\,
            ce => \N__16179\,
            sr => \N__23243\
        );

    \transmit_module.BRAM_ADDR__i12_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16335\,
            in1 => \N__16318\,
            in2 => \_gnd_net_\,
            in3 => \N__16188\,
            lcout => \TX_ADDR_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24102\,
            ce => \N__16179\,
            sr => \N__23243\
        );

    \receive_module.rx_counter.i246_2_lut_rep_15_2_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19645\,
            in2 => \_gnd_net_\,
            in3 => \N__20104\,
            lcout => \receive_module.n3671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18777\,
            in1 => \N__18833\,
            in2 => \N__19676\,
            in3 => \N__18918\,
            lcout => \line_buffer.n603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__18917\,
            in1 => \N__19641\,
            in2 => \N__18850\,
            in3 => \N__18776\,
            lcout => \line_buffer.n539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__18916\,
            in1 => \N__19649\,
            in2 => \N__18849\,
            in3 => \N__18778\,
            lcout => \line_buffer.n474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i9_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__20135\,
            in1 => \N__19667\,
            in2 => \N__17854\,
            in3 => \N__18069\,
            lcout => \RX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21968\,
            ce => 'H',
            sr => \N__19300\
        );

    \receive_module.BRAM_ADDR__i3_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__17817\,
            in1 => \N__20133\,
            in2 => \N__19684\,
            in3 => \N__17598\,
            lcout => \RX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21968\,
            ce => 'H',
            sr => \N__19300\
        );

    \receive_module.BRAM_ADDR__i4_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__17571\,
            in1 => \N__20136\,
            in2 => \N__17361\,
            in3 => \N__19659\,
            lcout => \RX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21968\,
            ce => 'H',
            sr => \N__19300\
        );

    \receive_module.BRAM_ADDR__i8_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__20138\,
            in1 => \N__17100\,
            in2 => \N__19686\,
            in3 => \N__17319\,
            lcout => \RX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21968\,
            ce => 'H',
            sr => \N__19300\
        );

    \receive_module.BRAM_ADDR__i6_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__20134\,
            in1 => \N__19660\,
            in2 => \N__16857\,
            in3 => \N__17073\,
            lcout => \RX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21968\,
            ce => 'H',
            sr => \N__19300\
        );

    \receive_module.BRAM_ADDR__i7_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__20137\,
            in1 => \N__16599\,
            in2 => \N__19685\,
            in3 => \N__16818\,
            lcout => \RX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21968\,
            ce => 'H',
            sr => \N__19300\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2257_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22754\,
            in1 => \N__16572\,
            in2 => \N__21497\,
            in3 => \N__16551\,
            lcout => \line_buffer.n3587\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3623_bdd_4_lut_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__21458\,
            in1 => \N__18438\,
            in2 => \N__18414\,
            in3 => \N__19200\,
            lcout => \line_buffer.n3626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3587_bdd_4_lut_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__18393\,
            in1 => \N__21459\,
            in2 => \N__18381\,
            in3 => \N__18360\,
            lcout => OPEN,
            ltout => \line_buffer.n3590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i3_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21293\,
            in2 => \N__18354\,
            in3 => \N__18351\,
            lcout => \TX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23771\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i4_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18345\,
            lcout => n1815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23653\,
            ce => 'H',
            sr => \N__22426\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18930\,
            in1 => \N__19680\,
            in2 => \N__18872\,
            in3 => \N__18789\,
            lcout => \line_buffer.n602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21999\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_DEBUG_c_3_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PULSE_1HZ_I_0_2_lut_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18176\,
            in2 => \_gnd_net_\,
            in3 => \N__18966\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i1_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i9_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18114\,
            lcout => \tvp_video_buffer.BUFFER_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.Y__i0_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18624\,
            in2 => \_gnd_net_\,
            in3 => \N__18603\,
            lcout => \receive_module.rx_counter.Y_0\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \receive_module.rx_counter.n3172\,
            clk => \N__21930\,
            ce => \N__20022\,
            sr => \N__19299\
        );

    \receive_module.rx_counter.Y__i1_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18599\,
            in2 => \_gnd_net_\,
            in3 => \N__18576\,
            lcout => \receive_module.rx_counter.Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3172\,
            carryout => \receive_module.rx_counter.n3173\,
            clk => \N__21930\,
            ce => \N__20022\,
            sr => \N__19299\
        );

    \receive_module.rx_counter.Y__i2_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18573\,
            in2 => \_gnd_net_\,
            in3 => \N__18552\,
            lcout => \receive_module.rx_counter.Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3173\,
            carryout => \receive_module.rx_counter.n3174\,
            clk => \N__21930\,
            ce => \N__20022\,
            sr => \N__19299\
        );

    \receive_module.rx_counter.Y__i3_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18545\,
            in2 => \_gnd_net_\,
            in3 => \N__18525\,
            lcout => \receive_module.rx_counter.Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3174\,
            carryout => \receive_module.rx_counter.n3175\,
            clk => \N__21930\,
            ce => \N__20022\,
            sr => \N__19299\
        );

    \receive_module.rx_counter.Y__i4_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18522\,
            in2 => \_gnd_net_\,
            in3 => \N__18504\,
            lcout => \receive_module.rx_counter.Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3175\,
            carryout => \receive_module.rx_counter.n3176\,
            clk => \N__21930\,
            ce => \N__20022\,
            sr => \N__19299\
        );

    \receive_module.rx_counter.Y__i5_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18501\,
            in2 => \_gnd_net_\,
            in3 => \N__18486\,
            lcout => \receive_module.rx_counter.Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3176\,
            carryout => \receive_module.rx_counter.n3177\,
            clk => \N__21930\,
            ce => \N__20022\,
            sr => \N__19299\
        );

    \receive_module.rx_counter.Y__i6_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18483\,
            in2 => \_gnd_net_\,
            in3 => \N__18465\,
            lcout => \receive_module.rx_counter.Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3177\,
            carryout => \receive_module.rx_counter.n3178\,
            clk => \N__21930\,
            ce => \N__20022\,
            sr => \N__19299\
        );

    \receive_module.rx_counter.Y__i7_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18462\,
            in2 => \_gnd_net_\,
            in3 => \N__18441\,
            lcout => \receive_module.rx_counter.Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3178\,
            carryout => \receive_module.rx_counter.n3179\,
            clk => \N__21930\,
            ce => \N__20022\,
            sr => \N__19299\
        );

    \receive_module.rx_counter.Y__i8_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19190\,
            in2 => \_gnd_net_\,
            in3 => \N__19194\,
            lcout => \receive_module.rx_counter.Y_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21935\,
            ce => \N__20018\,
            sr => \N__19298\
        );

    \tvp_video_buffer.WIRE_OUT_i0_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19164\,
            lcout => \RX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_26_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19055\,
            in2 => \_gnd_net_\,
            in3 => \N__19043\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n7_adj_619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_4_lut_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__19031\,
            in1 => \N__19019\,
            in2 => \N__19008\,
            in3 => \N__19005\,
            lcout => \receive_module.rx_counter.n11\,
            ltout => \receive_module.rx_counter.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1304_2_lut_3_lut_3_lut_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__18999\,
            in1 => \_gnd_net_\,
            in2 => \N__18984\,
            in3 => \N__20079\,
            lcout => \receive_module.rx_counter.n2547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.PULSE_1HZ_49_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__18972\,
            in1 => \N__18959\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PULSE_1HZ\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__18948\,
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18929\,
            in1 => \N__19594\,
            in2 => \N__18873\,
            in3 => \N__18788\,
            lcout => \line_buffer.n538\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18690\,
            lcout => \transmit_module.X_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24251\,
            ce => \N__18662\,
            sr => \N__20515\
        );

    \tvp_video_buffer.BUFFER_0__i7_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i6_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19812\,
            lcout => \RX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i15_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19818\,
            lcout => \tvp_video_buffer.BUFFER_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2281_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22707\,
            in1 => \N__19806\,
            in2 => \N__21464\,
            in3 => \N__19791\,
            lcout => OPEN,
            ltout => \line_buffer.n3593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3593_bdd_4_lut_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__19779\,
            in1 => \N__19764\,
            in2 => \N__19743\,
            in3 => \N__21414\,
            lcout => \line_buffer.n3596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2291_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__22633\,
            in1 => \N__19740\,
            in2 => \N__21463\,
            in3 => \N__19731\,
            lcout => \line_buffer.n3629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i5_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__20129\,
            in1 => \N__19713\,
            in2 => \N__19690\,
            in3 => \N__19329\,
            lcout => \RX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21965\,
            ce => 'H',
            sr => \N__19301\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2286_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22753\,
            in1 => \N__19227\,
            in2 => \N__21499\,
            in3 => \N__19212\,
            lcout => \line_buffer.n3623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_hs_buffer.BUFFER_0__i2_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20151\,
            lcout => \tvp_hs_buffer.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20168\,
            lcout => \tvp_hs_buffer.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_hs_buffer.WIRE_OUT_0__9_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20145\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \TVP_HSYNC_buff\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i249_3_lut_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__19983\,
            in1 => \N__19999\,
            in2 => \_gnd_net_\,
            in3 => \N__20100\,
            lcout => \receive_module.rx_counter.n2078\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_HS_51_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20000\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.rx_counter.old_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i92_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21141\,
            lcout => \transmit_module.Y_DELTA_PATTERN_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24314\,
            ce => \N__23395\,
            sr => \N__23283\
        );

    \transmit_module.Y_DELTA_PATTERN_i97_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19977\,
            lcout => \transmit_module.Y_DELTA_PATTERN_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24220\,
            ce => \N__23387\,
            sr => \N__23285\
        );

    \transmit_module.Y_DELTA_PATTERN_i98_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24220\,
            ce => \N__23387\,
            sr => \N__23285\
        );

    \transmit_module.Y_DELTA_PATTERN_i89_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20640\,
            lcout => \transmit_module.Y_DELTA_PATTERN_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24220\,
            ce => \N__23387\,
            sr => \N__23285\
        );

    \transmit_module.Y_DELTA_PATTERN_i88_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19971\,
            lcout => \transmit_module.Y_DELTA_PATTERN_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24220\,
            ce => \N__23387\,
            sr => \N__23285\
        );

    \transmit_module.Y_DELTA_PATTERN_i91_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20652\,
            lcout => \transmit_module.Y_DELTA_PATTERN_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24220\,
            ce => \N__23387\,
            sr => \N__23285\
        );

    \transmit_module.Y_DELTA_PATTERN_i90_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20646\,
            lcout => \transmit_module.Y_DELTA_PATTERN_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24220\,
            ce => \N__23387\,
            sr => \N__23285\
        );

    \transmit_module.Y_DELTA_PATTERN_i99_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20634\,
            lcout => \transmit_module.Y_DELTA_PATTERN_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24227\,
            ce => \N__20516\,
            sr => \N__23282\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22755\,
            in1 => \N__20370\,
            in2 => \N__21505\,
            in3 => \N__20352\,
            lcout => \line_buffer.n3653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3629_bdd_4_lut_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__20337\,
            in1 => \N__21478\,
            in2 => \N__20319\,
            in3 => \N__20301\,
            lcout => \line_buffer.n3632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2296_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22723\,
            in1 => \N__20295\,
            in2 => \N__21502\,
            in3 => \N__20277\,
            lcout => OPEN,
            ltout => \line_buffer.n3635_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3635_bdd_4_lut_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__20262\,
            in1 => \N__20241\,
            in2 => \N__20223\,
            in3 => \N__21479\,
            lcout => \line_buffer.n3638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3653_bdd_4_lut_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001100"
        )
    port map (
            in0 => \N__20220\,
            in1 => \N__20205\,
            in2 => \N__21503\,
            in3 => \N__20190\,
            lcout => OPEN,
            ltout => \line_buffer.n3656_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i5_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21267\,
            in2 => \N__20934\,
            in3 => \N__20931\,
            lcout => \TX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i0_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21268\,
            in1 => \N__20781\,
            in2 => \_gnd_net_\,
            in3 => \N__20925\,
            lcout => \TX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3647_bdd_4_lut_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__20907\,
            in1 => \N__20829\,
            in2 => \N__20886\,
            in3 => \N__21483\,
            lcout => OPEN,
            ltout => \line_buffer.n3650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i1_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20865\,
            in2 => \N__20859\,
            in3 => \N__21269\,
            lcout => \TX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2306_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22759\,
            in1 => \N__20856\,
            in2 => \N__21501\,
            in3 => \N__20844\,
            lcout => \line_buffer.n3647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3641_bdd_4_lut_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__21474\,
            in1 => \N__20823\,
            in2 => \N__20805\,
            in3 => \N__21090\,
            lcout => \line_buffer.n3644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i6_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20775\,
            lcout => n1813,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23772\,
            ce => 'H',
            sr => \N__22425\
        );

    \transmit_module.VGA_R__i2_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20709\,
            lcout => n1817,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23815\,
            ce => 'H',
            sr => \N__22427\
        );

    \transmit_module.Y_DELTA_PATTERN_i96_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20658\,
            lcout => \transmit_module.Y_DELTA_PATTERN_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24213\,
            ce => \N__23391\,
            sr => \N__23280\
        );

    \transmit_module.Y_DELTA_PATTERN_i94_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21153\,
            lcout => \transmit_module.Y_DELTA_PATTERN_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24213\,
            ce => \N__23391\,
            sr => \N__23280\
        );

    \transmit_module.Y_DELTA_PATTERN_i95_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21159\,
            lcout => \transmit_module.Y_DELTA_PATTERN_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24213\,
            ce => \N__23391\,
            sr => \N__23280\
        );

    \transmit_module.Y_DELTA_PATTERN_i93_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21147\,
            lcout => \transmit_module.Y_DELTA_PATTERN_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24213\,
            ce => \N__23391\,
            sr => \N__23280\
        );

    \transmit_module.Y_DELTA_PATTERN_i83_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21774\,
            lcout => \transmit_module.Y_DELTA_PATTERN_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24213\,
            ce => \N__23391\,
            sr => \N__23280\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2301_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22769\,
            in1 => \N__21126\,
            in2 => \N__21504\,
            in3 => \N__21111\,
            lcout => \line_buffer.n3641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2196_3_lut_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22833\,
            in1 => \N__21084\,
            in2 => \_gnd_net_\,
            in3 => \N__21072\,
            lcout => \line_buffer.n3533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i7_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22005\,
            lcout => \RX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2212_3_lut_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20961\,
            in1 => \N__20949\,
            in2 => \_gnd_net_\,
            in3 => \N__22825\,
            lcout => \line_buffer.n3549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2276_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__21506\,
            in1 => \N__22839\,
            in2 => \N__21299\,
            in3 => \N__21762\,
            lcout => OPEN,
            ltout => \line_buffer.n3611_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i4_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__21283\,
            in1 => \N__21750\,
            in2 => \N__21741\,
            in3 => \N__21549\,
            lcout => \TX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i4_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21633\,
            lcout => \RX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i13_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21585\,
            lcout => \tvp_video_buffer.BUFFER_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i5_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21623\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2211_3_lut_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21579\,
            in1 => \N__21564\,
            in2 => \_gnd_net_\,
            in3 => \N__22771\,
            lcout => \line_buffer.n3548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2236_3_lut_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21540\,
            in1 => \N__21528\,
            in2 => \_gnd_net_\,
            in3 => \N__22770\,
            lcout => \line_buffer.n3573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2271_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__21500\,
            in1 => \N__21324\,
            in2 => \N__21295\,
            in3 => \N__22566\,
            lcout => \line_buffer.n3605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i6_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__22335\,
            in1 => \N__21312\,
            in2 => \N__21305\,
            in3 => \N__21165\,
            lcout => \TX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i5_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22560\,
            lcout => n1814,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23957\,
            ce => 'H',
            sr => \N__22431\
        );

    \transmit_module.VGA_R__i7_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22494\,
            lcout => n1812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23957\,
            ce => 'H',
            sr => \N__22431\
        );

    \line_buffer.i2235_3_lut_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22362\,
            in1 => \N__22347\,
            in2 => \_gnd_net_\,
            in3 => \N__22807\,
            lcout => \line_buffer.n3572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_20_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i8_LC_21_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22026\,
            lcout => \tvp_video_buffer.BUFFER_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i16_LC_21_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22011\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21949\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i87_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21783\,
            lcout => \transmit_module.Y_DELTA_PATTERN_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24295\,
            ce => \N__23396\,
            sr => \N__23281\
        );

    \transmit_module.Y_DELTA_PATTERN_i84_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24381\,
            lcout => \transmit_module.Y_DELTA_PATTERN_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24315\,
            ce => \N__23397\,
            sr => \N__23325\
        );

    \transmit_module.Y_DELTA_PATTERN_i85_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24369\,
            lcout => \transmit_module.Y_DELTA_PATTERN_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24315\,
            ce => \N__23397\,
            sr => \N__23325\
        );

    \transmit_module.Y_DELTA_PATTERN_i86_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24315\,
            ce => \N__23397\,
            sr => \N__23325\
        );

    \line_buffer.i2197_3_lut_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22768\,
            in1 => \N__22869\,
            in2 => \_gnd_net_\,
            in3 => \N__22854\,
            lcout => \line_buffer.n3534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2202_3_lut_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22798\,
            in1 => \N__22602\,
            in2 => \_gnd_net_\,
            in3 => \N__22587\,
            lcout => \line_buffer.n3539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
