// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 14 2018 01:24:34

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "main" view "INTERFACE"

module main (
    TVP_VIDEO,
    ADV_B,
    ADV_G,
    ADV_R,
    DEBUG,
    TVP_CLK,
    ADV_CLK,
    TVP_HSYNC,
    ADV_HSYNC,
    TVP_VSYNC,
    ADV_VSYNC,
    ADV_BLANK_N,
    LED,
    ADV_SYNC_N);

    input [9:0] TVP_VIDEO;
    output [7:0] ADV_B;
    output [7:0] ADV_G;
    output [7:0] ADV_R;
    inout [7:0] DEBUG;
    input TVP_CLK;
    output ADV_CLK;
    input TVP_HSYNC;
    output ADV_HSYNC;
    input TVP_VSYNC;
    output ADV_VSYNC;
    output ADV_BLANK_N;
    output LED;
    output ADV_SYNC_N;

    wire N__18943;
    wire N__18942;
    wire N__18941;
    wire N__18932;
    wire N__18931;
    wire N__18930;
    wire N__18923;
    wire N__18922;
    wire N__18921;
    wire N__18914;
    wire N__18913;
    wire N__18912;
    wire N__18905;
    wire N__18904;
    wire N__18903;
    wire N__18896;
    wire N__18895;
    wire N__18894;
    wire N__18887;
    wire N__18886;
    wire N__18885;
    wire N__18878;
    wire N__18877;
    wire N__18876;
    wire N__18869;
    wire N__18868;
    wire N__18867;
    wire N__18860;
    wire N__18859;
    wire N__18858;
    wire N__18851;
    wire N__18850;
    wire N__18849;
    wire N__18842;
    wire N__18841;
    wire N__18840;
    wire N__18833;
    wire N__18832;
    wire N__18831;
    wire N__18824;
    wire N__18823;
    wire N__18822;
    wire N__18815;
    wire N__18814;
    wire N__18813;
    wire N__18806;
    wire N__18805;
    wire N__18804;
    wire N__18797;
    wire N__18796;
    wire N__18795;
    wire N__18788;
    wire N__18787;
    wire N__18786;
    wire N__18779;
    wire N__18778;
    wire N__18777;
    wire N__18770;
    wire N__18769;
    wire N__18768;
    wire N__18761;
    wire N__18760;
    wire N__18759;
    wire N__18752;
    wire N__18751;
    wire N__18750;
    wire N__18743;
    wire N__18742;
    wire N__18741;
    wire N__18734;
    wire N__18733;
    wire N__18732;
    wire N__18725;
    wire N__18724;
    wire N__18723;
    wire N__18716;
    wire N__18715;
    wire N__18714;
    wire N__18707;
    wire N__18706;
    wire N__18705;
    wire N__18698;
    wire N__18697;
    wire N__18696;
    wire N__18689;
    wire N__18688;
    wire N__18687;
    wire N__18680;
    wire N__18679;
    wire N__18678;
    wire N__18671;
    wire N__18670;
    wire N__18669;
    wire N__18662;
    wire N__18661;
    wire N__18660;
    wire N__18653;
    wire N__18652;
    wire N__18651;
    wire N__18644;
    wire N__18643;
    wire N__18642;
    wire N__18635;
    wire N__18634;
    wire N__18633;
    wire N__18626;
    wire N__18625;
    wire N__18624;
    wire N__18617;
    wire N__18616;
    wire N__18615;
    wire N__18608;
    wire N__18607;
    wire N__18606;
    wire N__18599;
    wire N__18598;
    wire N__18597;
    wire N__18590;
    wire N__18589;
    wire N__18588;
    wire N__18581;
    wire N__18580;
    wire N__18579;
    wire N__18572;
    wire N__18571;
    wire N__18570;
    wire N__18563;
    wire N__18562;
    wire N__18561;
    wire N__18554;
    wire N__18553;
    wire N__18552;
    wire N__18545;
    wire N__18544;
    wire N__18543;
    wire N__18536;
    wire N__18535;
    wire N__18534;
    wire N__18527;
    wire N__18526;
    wire N__18525;
    wire N__18518;
    wire N__18517;
    wire N__18516;
    wire N__18509;
    wire N__18508;
    wire N__18507;
    wire N__18490;
    wire N__18489;
    wire N__18488;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18477;
    wire N__18476;
    wire N__18475;
    wire N__18474;
    wire N__18473;
    wire N__18472;
    wire N__18471;
    wire N__18470;
    wire N__18469;
    wire N__18466;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18451;
    wire N__18450;
    wire N__18449;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18441;
    wire N__18440;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18386;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18368;
    wire N__18363;
    wire N__18360;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18322;
    wire N__18317;
    wire N__18310;
    wire N__18303;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18236;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18192;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18184;
    wire N__18181;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18156;
    wire N__18151;
    wire N__18150;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18139;
    wire N__18138;
    wire N__18137;
    wire N__18136;
    wire N__18135;
    wire N__18130;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18108;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18084;
    wire N__18077;
    wire N__18070;
    wire N__18069;
    wire N__18068;
    wire N__18067;
    wire N__18064;
    wire N__18059;
    wire N__18056;
    wire N__18055;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18007;
    wire N__18004;
    wire N__17999;
    wire N__17992;
    wire N__17989;
    wire N__17980;
    wire N__17979;
    wire N__17976;
    wire N__17975;
    wire N__17974;
    wire N__17973;
    wire N__17972;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17943;
    wire N__17940;
    wire N__17937;
    wire N__17934;
    wire N__17931;
    wire N__17926;
    wire N__17925;
    wire N__17922;
    wire N__17919;
    wire N__17916;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17897;
    wire N__17892;
    wire N__17887;
    wire N__17878;
    wire N__17877;
    wire N__17876;
    wire N__17875;
    wire N__17874;
    wire N__17873;
    wire N__17872;
    wire N__17871;
    wire N__17870;
    wire N__17869;
    wire N__17868;
    wire N__17867;
    wire N__17866;
    wire N__17865;
    wire N__17862;
    wire N__17861;
    wire N__17858;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17846;
    wire N__17839;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17806;
    wire N__17803;
    wire N__17796;
    wire N__17789;
    wire N__17784;
    wire N__17781;
    wire N__17780;
    wire N__17777;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17754;
    wire N__17749;
    wire N__17746;
    wire N__17737;
    wire N__17736;
    wire N__17733;
    wire N__17730;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17713;
    wire N__17712;
    wire N__17709;
    wire N__17706;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17694;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17686;
    wire N__17685;
    wire N__17684;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17672;
    wire N__17669;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17657;
    wire N__17652;
    wire N__17651;
    wire N__17650;
    wire N__17649;
    wire N__17646;
    wire N__17641;
    wire N__17636;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17589;
    wire N__17588;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17580;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17559;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17548;
    wire N__17541;
    wire N__17538;
    wire N__17535;
    wire N__17532;
    wire N__17531;
    wire N__17530;
    wire N__17529;
    wire N__17522;
    wire N__17519;
    wire N__17518;
    wire N__17517;
    wire N__17516;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17499;
    wire N__17498;
    wire N__17497;
    wire N__17496;
    wire N__17495;
    wire N__17492;
    wire N__17491;
    wire N__17490;
    wire N__17485;
    wire N__17482;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17474;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17457;
    wire N__17454;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17436;
    wire N__17435;
    wire N__17434;
    wire N__17429;
    wire N__17426;
    wire N__17425;
    wire N__17424;
    wire N__17423;
    wire N__17420;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17412;
    wire N__17411;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17397;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17385;
    wire N__17382;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17341;
    wire N__17338;
    wire N__17337;
    wire N__17334;
    wire N__17333;
    wire N__17332;
    wire N__17331;
    wire N__17330;
    wire N__17329;
    wire N__17328;
    wire N__17327;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17313;
    wire N__17312;
    wire N__17311;
    wire N__17306;
    wire N__17301;
    wire N__17292;
    wire N__17287;
    wire N__17282;
    wire N__17277;
    wire N__17272;
    wire N__17269;
    wire N__17268;
    wire N__17265;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17250;
    wire N__17249;
    wire N__17246;
    wire N__17245;
    wire N__17242;
    wire N__17241;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17226;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17214;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17200;
    wire N__17197;
    wire N__17196;
    wire N__17195;
    wire N__17190;
    wire N__17187;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17140;
    wire N__17137;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17085;
    wire N__17080;
    wire N__17075;
    wire N__17068;
    wire N__17065;
    wire N__17060;
    wire N__17055;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17033;
    wire N__17030;
    wire N__17023;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16962;
    wire N__16959;
    wire N__16956;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16944;
    wire N__16941;
    wire N__16938;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16770;
    wire N__16767;
    wire N__16764;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16736;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16686;
    wire N__16683;
    wire N__16680;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16644;
    wire N__16641;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16513;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16482;
    wire N__16481;
    wire N__16480;
    wire N__16479;
    wire N__16476;
    wire N__16475;
    wire N__16472;
    wire N__16471;
    wire N__16470;
    wire N__16467;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16452;
    wire N__16449;
    wire N__16446;
    wire N__16445;
    wire N__16444;
    wire N__16443;
    wire N__16440;
    wire N__16433;
    wire N__16432;
    wire N__16427;
    wire N__16424;
    wire N__16415;
    wire N__16410;
    wire N__16407;
    wire N__16406;
    wire N__16405;
    wire N__16402;
    wire N__16399;
    wire N__16392;
    wire N__16387;
    wire N__16386;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16354;
    wire N__16353;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16317;
    wire N__16314;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16272;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16260;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16151;
    wire N__16150;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16129;
    wire N__16126;
    wire N__16125;
    wire N__16124;
    wire N__16123;
    wire N__16122;
    wire N__16121;
    wire N__16120;
    wire N__16119;
    wire N__16118;
    wire N__16115;
    wire N__16114;
    wire N__16113;
    wire N__16112;
    wire N__16111;
    wire N__16110;
    wire N__16109;
    wire N__16108;
    wire N__16107;
    wire N__16106;
    wire N__16105;
    wire N__16104;
    wire N__16103;
    wire N__16102;
    wire N__16101;
    wire N__16100;
    wire N__16099;
    wire N__16098;
    wire N__16097;
    wire N__16096;
    wire N__16095;
    wire N__16094;
    wire N__16093;
    wire N__16092;
    wire N__16091;
    wire N__16090;
    wire N__16089;
    wire N__16088;
    wire N__16087;
    wire N__16086;
    wire N__16085;
    wire N__16084;
    wire N__16083;
    wire N__16082;
    wire N__16081;
    wire N__16080;
    wire N__16079;
    wire N__16078;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15978;
    wire N__15975;
    wire N__15972;
    wire N__15969;
    wire N__15968;
    wire N__15967;
    wire N__15966;
    wire N__15965;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15933;
    wire N__15928;
    wire N__15925;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15853;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15837;
    wire N__15836;
    wire N__15835;
    wire N__15834;
    wire N__15831;
    wire N__15830;
    wire N__15827;
    wire N__15826;
    wire N__15825;
    wire N__15822;
    wire N__15819;
    wire N__15814;
    wire N__15813;
    wire N__15812;
    wire N__15811;
    wire N__15810;
    wire N__15809;
    wire N__15808;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15794;
    wire N__15789;
    wire N__15786;
    wire N__15785;
    wire N__15782;
    wire N__15781;
    wire N__15778;
    wire N__15777;
    wire N__15776;
    wire N__15773;
    wire N__15772;
    wire N__15769;
    wire N__15768;
    wire N__15761;
    wire N__15756;
    wire N__15751;
    wire N__15746;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15723;
    wire N__15720;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15708;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15670;
    wire N__15665;
    wire N__15656;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15567;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15453;
    wire N__15450;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15357;
    wire N__15356;
    wire N__15355;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15325;
    wire N__15322;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15213;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15119;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14973;
    wire N__14970;
    wire N__14967;
    wire N__14964;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14952;
    wire N__14949;
    wire N__14946;
    wire N__14943;
    wire N__14940;
    wire N__14937;
    wire N__14934;
    wire N__14931;
    wire N__14928;
    wire N__14925;
    wire N__14922;
    wire N__14919;
    wire N__14916;
    wire N__14913;
    wire N__14910;
    wire N__14907;
    wire N__14904;
    wire N__14901;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14873;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14855;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14830;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14749;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14682;
    wire N__14679;
    wire N__14676;
    wire N__14673;
    wire N__14670;
    wire N__14667;
    wire N__14664;
    wire N__14661;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14649;
    wire N__14646;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14513;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14466;
    wire N__14463;
    wire N__14460;
    wire N__14457;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14445;
    wire N__14444;
    wire N__14443;
    wire N__14442;
    wire N__14441;
    wire N__14440;
    wire N__14437;
    wire N__14436;
    wire N__14435;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14427;
    wire N__14426;
    wire N__14425;
    wire N__14424;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14413;
    wire N__14412;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14404;
    wire N__14403;
    wire N__14402;
    wire N__14399;
    wire N__14398;
    wire N__14397;
    wire N__14394;
    wire N__14391;
    wire N__14388;
    wire N__14385;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14362;
    wire N__14361;
    wire N__14360;
    wire N__14357;
    wire N__14352;
    wire N__14349;
    wire N__14348;
    wire N__14345;
    wire N__14342;
    wire N__14335;
    wire N__14332;
    wire N__14325;
    wire N__14320;
    wire N__14311;
    wire N__14308;
    wire N__14303;
    wire N__14300;
    wire N__14297;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14279;
    wire N__14264;
    wire N__14257;
    wire N__14254;
    wire N__14247;
    wire N__14242;
    wire N__14233;
    wire N__14230;
    wire N__14229;
    wire N__14226;
    wire N__14223;
    wire N__14220;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14185;
    wire N__14184;
    wire N__14183;
    wire N__14182;
    wire N__14181;
    wire N__14180;
    wire N__14179;
    wire N__14178;
    wire N__14177;
    wire N__14176;
    wire N__14175;
    wire N__14174;
    wire N__14173;
    wire N__14172;
    wire N__14171;
    wire N__14168;
    wire N__14167;
    wire N__14166;
    wire N__14165;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14149;
    wire N__14142;
    wire N__14141;
    wire N__14140;
    wire N__14139;
    wire N__14132;
    wire N__14131;
    wire N__14130;
    wire N__14125;
    wire N__14122;
    wire N__14113;
    wire N__14110;
    wire N__14103;
    wire N__14102;
    wire N__14101;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14050;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13911;
    wire N__13908;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13896;
    wire N__13893;
    wire N__13890;
    wire N__13887;
    wire N__13884;
    wire N__13881;
    wire N__13878;
    wire N__13875;
    wire N__13872;
    wire N__13869;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13834;
    wire N__13831;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13704;
    wire N__13701;
    wire N__13698;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13566;
    wire N__13563;
    wire N__13560;
    wire N__13557;
    wire N__13554;
    wire N__13551;
    wire N__13548;
    wire N__13545;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13507;
    wire N__13504;
    wire N__13501;
    wire N__13498;
    wire N__13495;
    wire N__13492;
    wire N__13489;
    wire N__13486;
    wire N__13485;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13473;
    wire N__13470;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13458;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13398;
    wire N__13395;
    wire N__13392;
    wire N__13389;
    wire N__13386;
    wire N__13383;
    wire N__13380;
    wire N__13377;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13353;
    wire N__13350;
    wire N__13347;
    wire N__13344;
    wire N__13341;
    wire N__13338;
    wire N__13335;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13274;
    wire N__13269;
    wire N__13266;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13227;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13149;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13022;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13004;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12988;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12816;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12776;
    wire N__12775;
    wire N__12772;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12758;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12739;
    wire N__12736;
    wire N__12733;
    wire N__12730;
    wire N__12727;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12643;
    wire N__12640;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12627;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12616;
    wire N__12615;
    wire N__12614;
    wire N__12607;
    wire N__12604;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12596;
    wire N__12595;
    wire N__12594;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12580;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12569;
    wire N__12568;
    wire N__12561;
    wire N__12558;
    wire N__12555;
    wire N__12554;
    wire N__12553;
    wire N__12546;
    wire N__12543;
    wire N__12540;
    wire N__12539;
    wire N__12538;
    wire N__12537;
    wire N__12536;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12522;
    wire N__12521;
    wire N__12514;
    wire N__12511;
    wire N__12508;
    wire N__12507;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12493;
    wire N__12490;
    wire N__12487;
    wire N__12486;
    wire N__12485;
    wire N__12478;
    wire N__12475;
    wire N__12472;
    wire N__12471;
    wire N__12470;
    wire N__12465;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12451;
    wire N__12444;
    wire N__12441;
    wire N__12438;
    wire N__12437;
    wire N__12436;
    wire N__12433;
    wire N__12426;
    wire N__12423;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12409;
    wire N__12408;
    wire N__12407;
    wire N__12404;
    wire N__12399;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12356;
    wire N__12353;
    wire N__12348;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12165;
    wire N__12162;
    wire N__12161;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12118;
    wire N__12115;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12086;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12064;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11967;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11854;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11835;
    wire N__11834;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11812;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11658;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11541;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11509;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10915;
    wire N__10912;
    wire N__10911;
    wire N__10906;
    wire N__10903;
    wire N__10902;
    wire N__10899;
    wire N__10898;
    wire N__10895;
    wire N__10890;
    wire N__10887;
    wire N__10882;
    wire N__10881;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10864;
    wire N__10861;
    wire N__10860;
    wire N__10857;
    wire N__10854;
    wire N__10849;
    wire N__10846;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10788;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10656;
    wire N__10653;
    wire N__10650;
    wire N__10647;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10635;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10612;
    wire N__10609;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10597;
    wire N__10594;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10500;
    wire N__10497;
    wire N__10494;
    wire N__10491;
    wire N__10488;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10345;
    wire N__10342;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10311;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10257;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10197;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10146;
    wire N__10143;
    wire N__10138;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10084;
    wire N__10081;
    wire N__10078;
    wire N__10077;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10026;
    wire N__10021;
    wire N__10020;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9960;
    wire N__9957;
    wire N__9956;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9934;
    wire N__9931;
    wire N__9930;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9898;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9883;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9873;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9759;
    wire N__9756;
    wire N__9753;
    wire N__9750;
    wire N__9747;
    wire N__9744;
    wire N__9741;
    wire N__9738;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9723;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9702;
    wire N__9699;
    wire N__9696;
    wire N__9693;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9658;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9630;
    wire N__9627;
    wire N__9626;
    wire N__9623;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9601;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9384;
    wire N__9381;
    wire N__9378;
    wire N__9375;
    wire N__9370;
    wire N__9367;
    wire N__9366;
    wire N__9363;
    wire N__9362;
    wire N__9359;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9337;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9092;
    wire N__9089;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9030;
    wire N__9027;
    wire N__9024;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8851;
    wire N__8848;
    wire N__8847;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8820;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8751;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8691;
    wire N__8688;
    wire N__8687;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8671;
    wire N__8668;
    wire N__8665;
    wire N__8656;
    wire N__8655;
    wire N__8654;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8636;
    wire N__8633;
    wire N__8626;
    wire N__8623;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8572;
    wire N__8569;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8557;
    wire N__8554;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8542;
    wire N__8539;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8502;
    wire N__8499;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8433;
    wire N__8430;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8394;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8262;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8245;
    wire N__8244;
    wire N__8243;
    wire N__8240;
    wire N__8235;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8157;
    wire N__8154;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8113;
    wire N__8110;
    wire N__8109;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8101;
    wire N__8098;
    wire N__8093;
    wire N__8090;
    wire N__8083;
    wire N__8082;
    wire N__8081;
    wire N__8080;
    wire N__8079;
    wire N__8076;
    wire N__8073;
    wire N__8068;
    wire N__8065;
    wire N__8056;
    wire N__8053;
    wire N__8052;
    wire N__8051;
    wire N__8050;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8036;
    wire N__8033;
    wire N__8026;
    wire N__8025;
    wire N__8024;
    wire N__8023;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8011;
    wire N__8008;
    wire N__7999;
    wire N__7998;
    wire N__7997;
    wire N__7994;
    wire N__7989;
    wire N__7984;
    wire N__7983;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7966;
    wire N__7963;
    wire N__7960;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7942;
    wire N__7939;
    wire N__7936;
    wire N__7933;
    wire N__7930;
    wire N__7927;
    wire N__7924;
    wire N__7921;
    wire N__7918;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7882;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7831;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7756;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7741;
    wire N__7738;
    wire N__7737;
    wire N__7734;
    wire N__7733;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7708;
    wire N__7705;
    wire N__7704;
    wire N__7703;
    wire N__7702;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7690;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7660;
    wire N__7657;
    wire N__7656;
    wire N__7653;
    wire N__7650;
    wire N__7645;
    wire N__7642;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7630;
    wire N__7627;
    wire N__7626;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7609;
    wire N__7606;
    wire N__7605;
    wire N__7604;
    wire N__7603;
    wire N__7600;
    wire N__7593;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7528;
    wire N__7525;
    wire N__7524;
    wire N__7523;
    wire N__7520;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7476;
    wire N__7475;
    wire N__7474;
    wire N__7471;
    wire N__7468;
    wire N__7463;
    wire N__7460;
    wire N__7453;
    wire N__7450;
    wire N__7449;
    wire N__7448;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7436;
    wire N__7433;
    wire N__7426;
    wire N__7425;
    wire N__7424;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7412;
    wire N__7409;
    wire N__7402;
    wire N__7401;
    wire N__7400;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7378;
    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7361;
    wire N__7358;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7251;
    wire N__7250;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7238;
    wire N__7231;
    wire N__7230;
    wire N__7229;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7217;
    wire N__7214;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7153;
    wire N__7150;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7138;
    wire N__7135;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7123;
    wire N__7120;
    wire N__7119;
    wire N__7118;
    wire N__7115;
    wire N__7110;
    wire N__7105;
    wire N__7102;
    wire N__7101;
    wire N__7100;
    wire N__7095;
    wire N__7092;
    wire N__7089;
    wire N__7084;
    wire N__7081;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7045;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7026;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6993;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6985;
    wire N__6982;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6889;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6881;
    wire N__6876;
    wire N__6873;
    wire N__6868;
    wire N__6867;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6852;
    wire N__6849;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6818;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6796;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6764;
    wire N__6759;
    wire N__6756;
    wire N__6751;
    wire N__6748;
    wire N__6747;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6736;
    wire N__6733;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6700;
    wire N__6697;
    wire N__6696;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6671;
    wire N__6668;
    wire N__6663;
    wire N__6660;
    wire N__6655;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6647;
    wire N__6646;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6634;
    wire N__6627;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6609;
    wire N__6608;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6544;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6536;
    wire N__6531;
    wire N__6528;
    wire N__6523;
    wire N__6522;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6514;
    wire N__6511;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6442;
    wire N__6441;
    wire N__6440;
    wire N__6437;
    wire N__6436;
    wire N__6433;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6403;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6389;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6359;
    wire N__6356;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6335;
    wire N__6332;
    wire N__6325;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6315;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6304;
    wire N__6301;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6289;
    wire N__6284;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6265;
    wire N__6262;
    wire N__6257;
    wire N__6252;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6223;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6195;
    wire N__6192;
    wire N__6191;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6171;
    wire N__6168;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6140;
    wire N__6137;
    wire N__6130;
    wire N__6127;
    wire N__6122;
    wire N__6117;
    wire N__6112;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6088;
    wire N__6083;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6069;
    wire N__6064;
    wire N__6063;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6044;
    wire N__6039;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6003;
    wire N__6002;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5994;
    wire N__5991;
    wire N__5990;
    wire N__5987;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire VCCG0;
    wire TVP_VIDEO_c_4;
    wire GNDG0;
    wire TVP_VIDEO_c_5;
    wire TVP_VIDEO_c_3;
    wire TVP_VIDEO_c_7;
    wire TVP_VIDEO_c_6;
    wire TVP_VIDEO_c_8;
    wire TVP_VIDEO_c_9;
    wire TVP_VIDEO_c_2;
    wire \line_buffer.n730 ;
    wire \line_buffer.n632 ;
    wire \line_buffer.n762 ;
    wire \line_buffer.n759 ;
    wire \line_buffer.n751 ;
    wire \receive_module.rx_counter.n2975_cascade_ ;
    wire \line_buffer.n698 ;
    wire \receive_module.rx_counter.n2900 ;
    wire \receive_module.rx_counter.n2900_cascade_ ;
    wire \receive_module.rx_counter.n2943 ;
    wire \receive_module.rx_counter.n10 ;
    wire bfn_10_14_0_;
    wire \receive_module.rx_counter.n9 ;
    wire \receive_module.rx_counter.n2782 ;
    wire \receive_module.rx_counter.n8 ;
    wire \receive_module.rx_counter.n2783 ;
    wire \receive_module.rx_counter.X_3 ;
    wire \receive_module.rx_counter.n2784 ;
    wire \receive_module.rx_counter.X_4 ;
    wire \receive_module.rx_counter.n2785 ;
    wire \receive_module.rx_counter.X_5 ;
    wire \receive_module.rx_counter.n2786 ;
    wire \receive_module.rx_counter.X_6 ;
    wire \receive_module.rx_counter.n2787 ;
    wire \receive_module.rx_counter.X_7 ;
    wire \receive_module.rx_counter.n2788 ;
    wire \receive_module.rx_counter.n2789 ;
    wire \receive_module.rx_counter.X_8 ;
    wire bfn_10_15_0_;
    wire \receive_module.rx_counter.n2790 ;
    wire \receive_module.rx_counter.X_9 ;
    wire n3184;
    wire \receive_module.rx_counter.n4_cascade_ ;
    wire \receive_module.rx_counter.n2986_cascade_ ;
    wire \receive_module.rx_counter.n2989_cascade_ ;
    wire \receive_module.rx_counter.n31_adj_572 ;
    wire \receive_module.rx_counter.n7 ;
    wire \receive_module.rx_counter.n3166 ;
    wire \receive_module.rx_counter.n2978_cascade_ ;
    wire \receive_module.rx_counter.n4_adj_571 ;
    wire bfn_12_12_0_;
    wire \receive_module.rx_counter.n2758 ;
    wire \receive_module.rx_counter.n2759 ;
    wire \receive_module.rx_counter.n2760 ;
    wire \receive_module.rx_counter.n2761 ;
    wire \receive_module.rx_counter.n2762 ;
    wire \receive_module.rx_counter.n2763 ;
    wire \receive_module.rx_counter.n2764 ;
    wire \receive_module.rx_counter.n2765 ;
    wire bfn_12_13_0_;
    wire \receive_module.rx_counter.Y_7 ;
    wire \receive_module.rx_counter.Y_4 ;
    wire \receive_module.rx_counter.Y_2 ;
    wire \receive_module.rx_counter.Y_8 ;
    wire \receive_module.rx_counter.n6_cascade_ ;
    wire \receive_module.rx_counter.Y_3 ;
    wire \line_buffer.n723 ;
    wire \line_buffer.n715 ;
    wire \transmit_module.video_signal_controller.n2972 ;
    wire \transmit_module.video_signal_controller.n3014 ;
    wire \transmit_module.video_signal_controller.n3186_cascade_ ;
    wire ADV_HSYNC_c;
    wire \transmit_module.video_signal_controller.n12 ;
    wire \transmit_module.video_signal_controller.n3182_cascade_ ;
    wire \transmit_module.video_signal_controller.n8 ;
    wire \transmit_module.X_DELTA_PATTERN_9 ;
    wire \transmit_module.X_DELTA_PATTERN_8 ;
    wire \line_buffer.n758 ;
    wire \line_buffer.n750 ;
    wire \receive_module.n2152 ;
    wire TVP_HSYNC_c;
    wire \receive_module.old_HS ;
    wire \transmit_module.video_signal_controller.n2484 ;
    wire \receive_module.rx_counter.Y_5 ;
    wire n2147_cascade_;
    wire \receive_module.rx_counter.Y_6 ;
    wire Y_0;
    wire Y_1;
    wire n5_cascade_;
    wire n3009;
    wire \transmit_module.video_signal_controller.VGA_X_0 ;
    wire bfn_13_15_0_;
    wire \transmit_module.video_signal_controller.VGA_X_1 ;
    wire \transmit_module.video_signal_controller.n2766 ;
    wire \transmit_module.video_signal_controller.VGA_X_2 ;
    wire \transmit_module.video_signal_controller.n2767 ;
    wire \transmit_module.video_signal_controller.VGA_X_3 ;
    wire \transmit_module.video_signal_controller.n2768 ;
    wire \transmit_module.video_signal_controller.VGA_X_4 ;
    wire \transmit_module.video_signal_controller.n2769 ;
    wire \transmit_module.video_signal_controller.n2770 ;
    wire \transmit_module.video_signal_controller.n2771 ;
    wire \transmit_module.video_signal_controller.n2772 ;
    wire \transmit_module.video_signal_controller.n2773 ;
    wire bfn_13_16_0_;
    wire \transmit_module.video_signal_controller.n2774 ;
    wire \transmit_module.video_signal_controller.n2775 ;
    wire \transmit_module.X_DELTA_PATTERN_13 ;
    wire \transmit_module.X_DELTA_PATTERN_10 ;
    wire \transmit_module.X_DELTA_PATTERN_12 ;
    wire \transmit_module.X_DELTA_PATTERN_11 ;
    wire \transmit_module.X_DELTA_PATTERN_7 ;
    wire \transmit_module.X_DELTA_PATTERN_15 ;
    wire \transmit_module.X_DELTA_PATTERN_14 ;
    wire \line_buffer.n754 ;
    wire \line_buffer.n746 ;
    wire \line_buffer.n682 ;
    wire \line_buffer.n3143_cascade_ ;
    wire \line_buffer.n690 ;
    wire \line_buffer.n694 ;
    wire \line_buffer.n686 ;
    wire \line_buffer.n3101 ;
    wire \line_buffer.n691 ;
    wire \line_buffer.n683 ;
    wire \line_buffer.n722 ;
    wire \line_buffer.n714 ;
    wire bfn_14_14_0_;
    wire \transmit_module.video_signal_controller.n2776 ;
    wire \transmit_module.video_signal_controller.n2777 ;
    wire \transmit_module.video_signal_controller.n2778 ;
    wire \transmit_module.video_signal_controller.n2779 ;
    wire \transmit_module.video_signal_controller.n2780 ;
    wire \transmit_module.video_signal_controller.n2781 ;
    wire n2147;
    wire \transmit_module.video_signal_controller.n2262 ;
    wire \transmit_module.video_signal_controller.VGA_Y_0 ;
    wire \transmit_module.video_signal_controller.n3022_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_8 ;
    wire \transmit_module.video_signal_controller.VGA_X_6 ;
    wire \transmit_module.video_signal_controller.VGA_X_5 ;
    wire \transmit_module.video_signal_controller.VGA_X_7 ;
    wire \transmit_module.video_signal_controller.VGA_Y_1 ;
    wire \transmit_module.video_signal_controller.VGA_Y_2 ;
    wire \transmit_module.video_signal_controller.VGA_Y_5 ;
    wire \transmit_module.video_signal_controller.VGA_Y_6 ;
    wire \transmit_module.X_DELTA_PATTERN_1 ;
    wire \transmit_module.X_DELTA_PATTERN_2 ;
    wire \transmit_module.X_DELTA_PATTERN_6 ;
    wire \transmit_module.X_DELTA_PATTERN_5 ;
    wire \transmit_module.X_DELTA_PATTERN_4 ;
    wire \transmit_module.X_DELTA_PATTERN_3 ;
    wire \line_buffer.n755 ;
    wire \line_buffer.n747 ;
    wire \line_buffer.n3031_cascade_ ;
    wire \line_buffer.n3030 ;
    wire \line_buffer.n3095_cascade_ ;
    wire \line_buffer.n3040 ;
    wire \line_buffer.n625 ;
    wire \line_buffer.n617 ;
    wire \line_buffer.n3089 ;
    wire \line_buffer.n3092_cascade_ ;
    wire \line_buffer.n3146 ;
    wire \line_buffer.n626 ;
    wire \line_buffer.n618 ;
    wire \line_buffer.n3039 ;
    wire \receive_module.rx_counter.n10_adj_570_cascade_ ;
    wire bfn_15_11_0_;
    wire \receive_module.rx_counter.FRAME_COUNTER_1 ;
    wire \receive_module.rx_counter.n2753 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_2 ;
    wire \receive_module.rx_counter.n2754 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_3 ;
    wire \receive_module.rx_counter.n2755 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_4 ;
    wire \receive_module.rx_counter.n2756 ;
    wire \receive_module.rx_counter.n2757 ;
    wire \receive_module.rx_counter.n2227 ;
    wire n1955;
    wire INVADV_R__i1C_net;
    wire TX_DATA_2;
    wire n1953;
    wire INVADV_R__i3C_net;
    wire \transmit_module.video_signal_controller.VGA_Y_4 ;
    wire \transmit_module.video_signal_controller.n3183 ;
    wire \transmit_module.video_signal_controller.VGA_Y_3 ;
    wire \transmit_module.video_signal_controller.n6 ;
    wire \transmit_module.video_signal_controller.VGA_X_9 ;
    wire \transmit_module.video_signal_controller.VGA_X_10 ;
    wire \transmit_module.video_signal_controller.VGA_VISIBLE_N_558_cascade_ ;
    wire \transmit_module.video_signal_controller.n18 ;
    wire VGA_VISIBLE_cascade_;
    wire \transmit_module.X_DELTA_PATTERN_0 ;
    wire bfn_15_17_0_;
    wire \transmit_module.n2740 ;
    wire \transmit_module.n2741 ;
    wire \transmit_module.n2742 ;
    wire \transmit_module.n2743 ;
    wire \transmit_module.n2744 ;
    wire \transmit_module.n2745 ;
    wire \transmit_module.n2746 ;
    wire \transmit_module.n2747 ;
    wire bfn_15_18_0_;
    wire \transmit_module.n2748 ;
    wire \transmit_module.n2749 ;
    wire \transmit_module.n2750 ;
    wire \transmit_module.n2751 ;
    wire \transmit_module.n2752 ;
    wire \transmit_module.n2200 ;
    wire DEBUG_c_6;
    wire \transmit_module.n382 ;
    wire n22;
    wire \transmit_module.n383 ;
    wire DEBUG_c_5;
    wire n23;
    wire \transmit_module.n384 ;
    wire DEBUG_c_4;
    wire n24;
    wire \transmit_module.n386 ;
    wire DEBUG_c_2;
    wire n26;
    wire \receive_module.rx_counter.FRAME_COUNTER_5 ;
    wire \receive_module.rx_counter.n10_adj_570 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_0 ;
    wire LED_c;
    wire \receive_module.old_VS ;
    wire \receive_module.n252 ;
    wire n1950;
    wire INVADV_R__i6C_net;
    wire n1954;
    wire TX_DATA_3;
    wire n1952;
    wire n1951;
    wire n1949;
    wire ADV_B_c;
    wire INVADV_R__i2C_net;
    wire n19;
    wire \transmit_module.n379 ;
    wire \transmit_module.TX_ADDR_9 ;
    wire \transmit_module.TX_ADDR_8 ;
    wire \transmit_module.n380 ;
    wire n20;
    wire \transmit_module.TX_ADDR_10 ;
    wire \transmit_module.n378 ;
    wire n18;
    wire \line_buffer.n3104 ;
    wire TX_DATA_6;
    wire GB_BUFFER_TVP_CLK_c_THRU_CO;
    wire \line_buffer.n689 ;
    wire \line_buffer.n681 ;
    wire \line_buffer.n3140_cascade_ ;
    wire TX_DATA_1;
    wire \line_buffer.n713 ;
    wire \line_buffer.n721 ;
    wire \line_buffer.n624 ;
    wire \line_buffer.n616 ;
    wire \line_buffer.n3107_cascade_ ;
    wire \line_buffer.n3110 ;
    wire \line_buffer.n745 ;
    wire \line_buffer.n753 ;
    wire \line_buffer.n3137 ;
    wire \line_buffer.n761 ;
    wire \transmit_module.n387 ;
    wire DEBUG_c_1;
    wire n27;
    wire DEBUG_c_7;
    wire \transmit_module.n381 ;
    wire n21;
    wire \transmit_module.n385 ;
    wire DEBUG_c_3;
    wire n25_adj_573;
    wire \line_buffer.n3028 ;
    wire \line_buffer.n3125_cascade_ ;
    wire TX_DATA_7;
    wire \line_buffer.n727 ;
    wire \line_buffer.n719 ;
    wire \line_buffer.n3043 ;
    wire \line_buffer.n726 ;
    wire \line_buffer.n718 ;
    wire \line_buffer.n629 ;
    wire \line_buffer.n621 ;
    wire \line_buffer.n3161_cascade_ ;
    wire \line_buffer.n3164 ;
    wire \line_buffer.n630 ;
    wire \line_buffer.n622 ;
    wire \line_buffer.n3042 ;
    wire CONSTANT_ONE_NET;
    wire \line_buffer.n623 ;
    wire \line_buffer.n615 ;
    wire \line_buffer.n720 ;
    wire \line_buffer.n712 ;
    wire \line_buffer.n3113 ;
    wire \line_buffer.n688 ;
    wire \line_buffer.n680 ;
    wire \line_buffer.n3122_cascade_ ;
    wire \line_buffer.n3116 ;
    wire TX_DATA_0;
    wire RX_ADDR_0;
    wire \receive_module.n136 ;
    wire bfn_18_14_0_;
    wire \receive_module.n2727 ;
    wire \receive_module.n2728 ;
    wire \receive_module.n2729 ;
    wire \receive_module.n2730 ;
    wire RX_ADDR_5;
    wire \receive_module.n131 ;
    wire \receive_module.n2731 ;
    wire \receive_module.n2732 ;
    wire RX_ADDR_7;
    wire \receive_module.n129 ;
    wire \receive_module.n2733 ;
    wire \receive_module.n2734 ;
    wire RX_ADDR_8;
    wire \receive_module.n128 ;
    wire bfn_18_15_0_;
    wire RX_ADDR_9;
    wire \receive_module.n127 ;
    wire \receive_module.n2735 ;
    wire \receive_module.n2736 ;
    wire \receive_module.n2737 ;
    wire \receive_module.n2738 ;
    wire \receive_module.n2739 ;
    wire \receive_module.n3181 ;
    wire \transmit_module.n388 ;
    wire ADV_VSYNC_c;
    wire DEBUG_c_0;
    wire VGA_VISIBLE;
    wire n28;
    wire \line_buffer.n744 ;
    wire \line_buffer.n752 ;
    wire \line_buffer.n3119 ;
    wire \line_buffer.n695 ;
    wire \line_buffer.n687 ;
    wire \line_buffer.n3027 ;
    wire \line_buffer.n725 ;
    wire \line_buffer.n717 ;
    wire \receive_module.n133 ;
    wire RX_ADDR_3;
    wire \receive_module.n134 ;
    wire RX_ADDR_2;
    wire \receive_module.n135 ;
    wire RX_ADDR_1;
    wire \line_buffer.n628 ;
    wire \line_buffer.n620 ;
    wire \line_buffer.n3149 ;
    wire \line_buffer.n3152_cascade_ ;
    wire TX_DATA_5;
    wire \line_buffer.n692 ;
    wire \line_buffer.n684 ;
    wire \line_buffer.n3024 ;
    wire \line_buffer.n3131_cascade_ ;
    wire TX_ADDR_13;
    wire TX_DATA_4;
    wire ADV_CLK_c;
    wire \line_buffer.n716 ;
    wire \line_buffer.n724 ;
    wire \line_buffer.n3046 ;
    wire \receive_module.n132 ;
    wire RX_ADDR_4;
    wire \receive_module.n130 ;
    wire RX_ADDR_6;
    wire \receive_module.n126 ;
    wire TVP_VSYNC_c;
    wire RX_ADDR_10;
    wire TVP_CLK_c;
    wire \receive_module.n3185 ;
    wire \line_buffer.n757 ;
    wire \line_buffer.n749 ;
    wire \line_buffer.n685 ;
    wire \line_buffer.n693 ;
    wire \line_buffer.n3155_cascade_ ;
    wire TX_ADDR_12;
    wire \line_buffer.n3158 ;
    wire \line_buffer.n627 ;
    wire \line_buffer.n619 ;
    wire \line_buffer.n3045 ;
    wire TX_ADDR_11;
    wire \line_buffer.n756 ;
    wire \line_buffer.n748 ;
    wire \line_buffer.n3025 ;
    wire \line_buffer.n729 ;
    wire \line_buffer.n697 ;
    wire RX_ADDR_12;
    wire RX_ADDR_11;
    wire RX_ADDR_13;
    wire n25;
    wire \line_buffer.n633 ;
    wire _gnd_net_;

    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \tx_pll.TX_PLL_inst .TEST_MODE=1'b0;
    defparam \tx_pll.TX_PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \tx_pll.TX_PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \tx_pll.TX_PLL_inst .FILTER_RANGE=3'b010;
    defparam \tx_pll.TX_PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \tx_pll.TX_PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \tx_pll.TX_PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \tx_pll.TX_PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \tx_pll.TX_PLL_inst .DIVR=4'b0000;
    defparam \tx_pll.TX_PLL_inst .DIVQ=3'b100;
    defparam \tx_pll.TX_PLL_inst .DIVF=7'b0100110;
    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \tx_pll.TX_PLL_inst  (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(ADV_CLK_c),
            .REFERENCECLK(N__10366),
            .RESETB(N__12536),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .PLLOUTGLOBAL());
    defparam \line_buffer.mem2_physical .WRITE_MODE=3;
    defparam \line_buffer.mem2_physical .READ_MODE=3;
    defparam \line_buffer.mem2_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem2_physical  (
            .RDATA({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,\line_buffer.n630 ,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,\line_buffer.n629 ,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .RADDR({N__10449,N__10983,N__10710,N__11640,N__9738,N__9459,N__9195,N__11364,N__8931,N__11919,N__13905}),
            .WADDR({N__16212,N__14607,N__12846,N__13098,N__16575,N__13341,N__16827,N__15426,N__15177,N__14943,N__13602}),
            .MASK({dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37}),
            .WDATA({dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,N__6514,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,N__6634,dangling_wire_49,dangling_wire_50,dangling_wire_51}),
            .RCLKE(),
            .RCLK(N__17397),
            .RE(N__12569),
            .WCLKE(),
            .WCLK(N__16118),
            .WE(N__17737));
    defparam \line_buffer.mem14_physical .WRITE_MODE=3;
    defparam \line_buffer.mem14_physical .READ_MODE=3;
    defparam \line_buffer.mem14_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem14_physical  (
            .RDATA({dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,\line_buffer.n717 ,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,\line_buffer.n716 ,dangling_wire_63,dangling_wire_64,dangling_wire_65}),
            .RADDR({N__10521,N__11055,N__10782,N__11712,N__9810,N__9531,N__9267,N__11436,N__9003,N__11991,N__13977}),
            .WADDR({N__16284,N__14679,N__12918,N__13170,N__16647,N__13413,N__16899,N__15498,N__15249,N__15015,N__13674}),
            .MASK({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .WDATA({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,N__6432,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,N__6304,dangling_wire_93,dangling_wire_94,dangling_wire_95}),
            .RCLKE(),
            .RCLK(N__17531),
            .RE(N__12471),
            .WCLKE(),
            .WCLK(N__16102),
            .WE(N__18235));
    defparam \line_buffer.mem8_physical .WRITE_MODE=3;
    defparam \line_buffer.mem8_physical .READ_MODE=3;
    defparam \line_buffer.mem8_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem8_physical  (
            .RDATA({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,\line_buffer.n620 ,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\line_buffer.n619 ,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .RADDR({N__10434,N__10962,N__10677,N__11631,N__9717,N__9432,N__9168,N__11343,N__8892,N__11898,N__13884}),
            .WADDR({N__16185,N__14580,N__12819,N__13059,N__16548,N__13320,N__16794,N__15399,N__15162,N__14916,N__13581}),
            .MASK({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .WDATA({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,N__6442,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,N__6324,dangling_wire_137,dangling_wire_138,dangling_wire_139}),
            .RCLKE(),
            .RCLK(N__17245),
            .RE(N__12627),
            .WCLKE(),
            .WCLK(N__16123),
            .WE(N__6746));
    defparam \line_buffer.mem28_physical .WRITE_MODE=3;
    defparam \line_buffer.mem28_physical .READ_MODE=3;
    defparam \line_buffer.mem28_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem28_physical  (
            .RDATA({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,\line_buffer.n721 ,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,\line_buffer.n720 ,dangling_wire_151,dangling_wire_152,dangling_wire_153}),
            .RADDR({N__10542,N__11070,N__10785,N__11739,N__9825,N__9540,N__9276,N__11451,N__9000,N__12006,N__13992}),
            .WADDR({N__16293,N__14688,N__12927,N__13167,N__16656,N__13428,N__16902,N__15507,N__15270,N__15024,N__13689}),
            .MASK({dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169}),
            .WDATA({dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,N__6171,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,N__6848,dangling_wire_181,dangling_wire_182,dangling_wire_183}),
            .RCLKE(),
            .RCLK(N__17268),
            .RE(N__12553),
            .WCLKE(),
            .WCLK(N__16100),
            .WE(N__6764));
    defparam \line_buffer.mem5_physical .WRITE_MODE=3;
    defparam \line_buffer.mem5_physical .READ_MODE=3;
    defparam \line_buffer.mem5_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem5_physical  (
            .RDATA({dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,\line_buffer.n727 ,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,\line_buffer.n726 ,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .RADDR({N__10470,N__10998,N__10713,N__11667,N__9753,N__9468,N__9204,N__11379,N__8928,N__11934,N__13920}),
            .WADDR({N__16221,N__14616,N__12855,N__13095,N__16584,N__13356,N__16830,N__15435,N__15198,N__14952,N__13617}),
            .MASK({dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213}),
            .WDATA({dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,N__6536,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,N__6647,dangling_wire_225,dangling_wire_226,dangling_wire_227}),
            .RCLKE(),
            .RCLK(N__17213),
            .RE(N__12615),
            .WCLKE(),
            .WCLK(N__16114),
            .WE(N__6796));
    defparam \line_buffer.mem11_physical .WRITE_MODE=3;
    defparam \line_buffer.mem11_physical .READ_MODE=3;
    defparam \line_buffer.mem11_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem11_physical  (
            .RDATA({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,\line_buffer.n685 ,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,\line_buffer.n684 ,dangling_wire_239,dangling_wire_240,dangling_wire_241}),
            .RADDR({N__10557,N__11091,N__10818,N__11748,N__9846,N__9567,N__9303,N__11472,N__9039,N__12027,N__14013}),
            .WADDR({N__16320,N__14715,N__12954,N__13206,N__16683,N__13449,N__16935,N__15534,N__15285,N__15051,N__13710}),
            .MASK({dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .WDATA({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,N__6389,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,N__6283,dangling_wire_269,dangling_wire_270,dangling_wire_271}),
            .RCLKE(),
            .RCLK(N__17579),
            .RE(N__12436),
            .WCLKE(),
            .WCLK(N__16088),
            .WE(N__18192));
    defparam \line_buffer.mem21_physical .WRITE_MODE=3;
    defparam \line_buffer.mem21_physical .READ_MODE=3;
    defparam \line_buffer.mem21_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem21_physical  (
            .RDATA({dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,\line_buffer.n747 ,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,\line_buffer.n746 ,dangling_wire_283,dangling_wire_284,dangling_wire_285}),
            .RADDR({N__10425,N__10959,N__10686,N__11616,N__9714,N__9435,N__9171,N__11340,N__8907,N__11895,N__13881}),
            .WADDR({N__16188,N__14583,N__12822,N__13074,N__16551,N__13317,N__16803,N__15402,N__15153,N__14919,N__13578}),
            .MASK({dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301}),
            .WDATA({dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,N__6112,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,N__6010,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .RCLKE(),
            .RCLK(N__17313),
            .RE(N__12595),
            .WCLKE(),
            .WCLK(N__16122),
            .WE(N__12161));
    defparam \line_buffer.mem12_physical .WRITE_MODE=3;
    defparam \line_buffer.mem12_physical .READ_MODE=3;
    defparam \line_buffer.mem12_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem12_physical  (
            .RDATA({dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,\line_buffer.n683 ,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,\line_buffer.n682 ,dangling_wire_327,dangling_wire_328,dangling_wire_329}),
            .RADDR({N__10545,N__11079,N__10806,N__11736,N__9834,N__9555,N__9291,N__11460,N__9027,N__12015,N__14001}),
            .WADDR({N__16308,N__14703,N__12942,N__13194,N__16671,N__13437,N__16923,N__15522,N__15273,N__15039,N__13698}),
            .MASK({dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345}),
            .WDATA({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,N__6069,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,N__6002,dangling_wire_357,dangling_wire_358,dangling_wire_359}),
            .RCLKE(),
            .RCLK(N__17559),
            .RE(N__12437),
            .WCLKE(),
            .WCLK(N__16095),
            .WE(N__18191));
    defparam \line_buffer.mem18_physical .WRITE_MODE=3;
    defparam \line_buffer.mem18_physical .READ_MODE=3;
    defparam \line_buffer.mem18_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem18_physical  (
            .RDATA({dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,\line_buffer.n626 ,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,\line_buffer.n625 ,dangling_wire_371,dangling_wire_372,dangling_wire_373}),
            .RADDR({N__10473,N__11007,N__10734,N__11664,N__9762,N__9483,N__9219,N__11388,N__8955,N__11943,N__13929}),
            .WADDR({N__16236,N__14631,N__12870,N__13122,N__16599,N__13365,N__16851,N__15450,N__15201,N__14967,N__13626}),
            .MASK({dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389}),
            .WDATA({dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,N__6101,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,N__6003,dangling_wire_401,dangling_wire_402,dangling_wire_403}),
            .RCLKE(),
            .RCLK(N__17457),
            .RE(N__12539),
            .WCLKE(),
            .WCLK(N__16111),
            .WE(N__17729));
    defparam \line_buffer.mem24_physical .WRITE_MODE=3;
    defparam \line_buffer.mem24_physical .READ_MODE=3;
    defparam \line_buffer.mem24_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem24_physical  (
            .RDATA({dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,\line_buffer.n691 ,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,\line_buffer.n690 ,dangling_wire_415,dangling_wire_416,dangling_wire_417}),
            .RADDR({N__10590,N__11118,N__10833,N__11785,N__9873,N__9588,N__9324,N__11499,N__9048,N__12054,N__14040}),
            .WADDR({N__16341,N__14736,N__12975,N__13215,N__16704,N__13476,N__16950,N__15555,N__15318,N__15072,N__13737}),
            .MASK({dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .WDATA({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,N__6038,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,N__5927,dangling_wire_445,dangling_wire_446,dangling_wire_447}),
            .RCLKE(),
            .RCLK(N__17587),
            .RE(N__12485),
            .WCLKE(),
            .WCLK(N__16083),
            .WE(N__6993));
    defparam \line_buffer.mem1_physical .WRITE_MODE=3;
    defparam \line_buffer.mem1_physical .READ_MODE=3;
    defparam \line_buffer.mem1_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem1_physical  (
            .RDATA({dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,\line_buffer.n719 ,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,\line_buffer.n718 ,dangling_wire_459,dangling_wire_460,dangling_wire_461}),
            .RADDR({N__10581,N__11115,N__10842,N__11772,N__9870,N__9591,N__9327,N__11496,N__9061,N__12051,N__14037}),
            .WADDR({N__16344,N__14739,N__12978,N__13228,N__16707,N__13473,N__16959,N__15558,N__15309,N__15075,N__13734}),
            .MASK({dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477}),
            .WDATA({dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,N__6493,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,N__6608,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .RCLKE(),
            .RCLK(N__17589),
            .RE(N__12408),
            .WCLKE(),
            .WCLK(N__16081),
            .WE(N__18244));
    defparam \line_buffer.mem15_physical .WRITE_MODE=3;
    defparam \line_buffer.mem15_physical .READ_MODE=3;
    defparam \line_buffer.mem15_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem15_physical  (
            .RDATA({dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,\line_buffer.n715 ,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,\line_buffer.n714 ,dangling_wire_503,dangling_wire_504,dangling_wire_505}),
            .RADDR({N__10509,N__11043,N__10770,N__11700,N__9798,N__9519,N__9255,N__11424,N__8991,N__11979,N__13965}),
            .WADDR({N__16272,N__14667,N__12906,N__13158,N__16635,N__13401,N__16887,N__15486,N__15237,N__15003,N__13662}),
            .MASK({dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521}),
            .WDATA({dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,N__6082,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,N__5994,dangling_wire_533,dangling_wire_534,dangling_wire_535}),
            .RCLKE(),
            .RCLK(N__17530),
            .RE(N__12506),
            .WCLKE(),
            .WCLK(N__16105),
            .WE(N__18236));
    defparam \line_buffer.mem27_physical .WRITE_MODE=3;
    defparam \line_buffer.mem27_physical .READ_MODE=3;
    defparam \line_buffer.mem27_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem27_physical  (
            .RDATA({dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,\line_buffer.n723 ,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,\line_buffer.n722 ,dangling_wire_547,dangling_wire_548,dangling_wire_549}),
            .RADDR({N__10554,N__11082,N__10797,N__11751,N__9837,N__9552,N__9288,N__11463,N__9012,N__12018,N__14004}),
            .WADDR({N__16305,N__14700,N__12939,N__13179,N__16668,N__13440,N__16914,N__15519,N__15282,N__15036,N__13701}),
            .MASK({dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565}),
            .WDATA({dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,N__6063,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,N__5958,dangling_wire_577,dangling_wire_578,dangling_wire_579}),
            .RCLKE(),
            .RCLK(N__17548),
            .RE(N__12522),
            .WCLKE(),
            .WCLK(N__16098),
            .WE(N__6788));
    defparam \line_buffer.mem22_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .WRITE_MODE=3;
    defparam \line_buffer.mem22_physical .READ_MODE=3;
    defparam \line_buffer.mem22_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem22_physical  (
            .RDATA({dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,\line_buffer.n745 ,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,\line_buffer.n744 ,dangling_wire_591,dangling_wire_592,dangling_wire_593}),
            .RADDR({N__10413,N__10947,N__10674,N__11604,N__9702,N__9423,N__9159,N__11328,N__8895,N__11883,N__13869}),
            .WADDR({N__16176,N__14571,N__12810,N__13062,N__16539,N__13305,N__16791,N__15390,N__15141,N__14907,N__13566}),
            .MASK({dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609}),
            .WDATA({dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,N__6223,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,N__6907,dangling_wire_621,dangling_wire_622,dangling_wire_623}),
            .RCLKE(),
            .RCLK(N__17226),
            .RE(N__12614),
            .WCLKE(),
            .WCLK(N__16124),
            .WE(N__12166));
    defparam \line_buffer.mem4_physical .WRITE_MODE=3;
    defparam \line_buffer.mem4_physical .READ_MODE=3;
    defparam \line_buffer.mem4_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem4_physical  (
            .RDATA({dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,\line_buffer.n695 ,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,\line_buffer.n694 ,dangling_wire_635,dangling_wire_636,dangling_wire_637}),
            .RADDR({N__10482,N__11010,N__10725,N__11679,N__9765,N__9480,N__9216,N__11391,N__8940,N__11946,N__13932}),
            .WADDR({N__16233,N__14628,N__12867,N__13107,N__16596,N__13368,N__16842,N__15447,N__15210,N__14964,N__13629}),
            .MASK({dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653}),
            .WDATA({dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,N__6521,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,N__6646,dangling_wire_665,dangling_wire_666,dangling_wire_667}),
            .RCLKE(),
            .RCLK(N__17425),
            .RE(N__12600),
            .WCLKE(),
            .WCLK(N__16112),
            .WE(N__6992));
    defparam \line_buffer.mem16_physical .WRITE_MODE=3;
    defparam \line_buffer.mem16_physical .READ_MODE=3;
    defparam \line_buffer.mem16_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem16_physical  (
            .RDATA({dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,\line_buffer.n713 ,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,\line_buffer.n712 ,dangling_wire_679,dangling_wire_680,dangling_wire_681}),
            .RADDR({N__10497,N__11031,N__10758,N__11688,N__9786,N__9507,N__9243,N__11412,N__8979,N__11967,N__13953}),
            .WADDR({N__16260,N__14655,N__12894,N__13146,N__16623,N__13389,N__16875,N__15474,N__15225,N__14991,N__13650}),
            .MASK({dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697}),
            .WDATA({dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,N__6222,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,N__6888,dangling_wire_709,dangling_wire_710,dangling_wire_711}),
            .RCLKE(),
            .RCLK(N__17499),
            .RE(N__12507),
            .WCLKE(),
            .WCLK(N__16107),
            .WE(N__18243));
    defparam \line_buffer.mem30_physical .WRITE_MODE=3;
    defparam \line_buffer.mem30_physical .READ_MODE=3;
    defparam \line_buffer.mem30_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem30_physical  (
            .RDATA({dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,\line_buffer.n755 ,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,\line_buffer.n754 ,dangling_wire_723,dangling_wire_724,dangling_wire_725}),
            .RADDR({N__10506,N__11034,N__10749,N__11703,N__9789,N__9504,N__9240,N__11415,N__8964,N__11970,N__13956}),
            .WADDR({N__16257,N__14652,N__12891,N__13131,N__16620,N__13392,N__16866,N__15471,N__15234,N__14988,N__13653}),
            .MASK({dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741}),
            .WDATA({dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,N__6088,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,N__5990,dangling_wire_753,dangling_wire_754,dangling_wire_755}),
            .RCLKE(),
            .RCLK(N__17481),
            .RE(N__12580),
            .WCLKE(),
            .WCLK(N__16108),
            .WE(N__6691));
    defparam \line_buffer.mem25_physical .WRITE_MODE=3;
    defparam \line_buffer.mem25_physical .READ_MODE=3;
    defparam \line_buffer.mem25_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem25_physical  (
            .RDATA({dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,\line_buffer.n689 ,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,\line_buffer.n688 ,dangling_wire_767,dangling_wire_768,dangling_wire_769}),
            .RADDR({N__10578,N__11106,N__10821,N__11775,N__9861,N__9576,N__9312,N__11487,N__9036,N__12042,N__14028}),
            .WADDR({N__16329,N__14724,N__12963,N__13203,N__16692,N__13464,N__16938,N__15543,N__15306,N__15060,N__13725}),
            .MASK({dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785}),
            .WDATA({dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,N__6190,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,N__6835,dangling_wire_797,dangling_wire_798,dangling_wire_799}),
            .RCLKE(),
            .RCLK(N__17572),
            .RE(N__12486),
            .WCLKE(),
            .WCLK(N__16086),
            .WE(N__6985));
    defparam \line_buffer.mem7_physical .WRITE_MODE=3;
    defparam \line_buffer.mem7_physical .READ_MODE=3;
    defparam \line_buffer.mem7_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem7_physical  (
            .RDATA({dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,\line_buffer.n622 ,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,\line_buffer.n621 ,dangling_wire_811,dangling_wire_812,dangling_wire_813}),
            .RADDR({N__10446,N__10974,N__10689,N__11643,N__9729,N__9444,N__9180,N__11355,N__8904,N__11910,N__13896}),
            .WADDR({N__16197,N__14592,N__12831,N__13071,N__16560,N__13332,N__16806,N__15411,N__15174,N__14928,N__13593}),
            .MASK({dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829}),
            .WDATA({dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,N__6544,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,N__6655,dangling_wire_841,dangling_wire_842,dangling_wire_843}),
            .RCLKE(),
            .RCLK(N__17225),
            .RE(N__12626),
            .WCLKE(),
            .WCLK(N__16121),
            .WE(N__6736));
    defparam \line_buffer.mem20_physical .WRITE_MODE=3;
    defparam \line_buffer.mem20_physical .READ_MODE=3;
    defparam \line_buffer.mem20_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem20_physical  (
            .RDATA({dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,\line_buffer.n749 ,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,\line_buffer.n748 ,dangling_wire_855,dangling_wire_856,dangling_wire_857}),
            .RADDR({N__10437,N__10971,N__10698,N__11628,N__9726,N__9447,N__9183,N__11352,N__8919,N__11907,N__13893}),
            .WADDR({N__16200,N__14595,N__12834,N__13086,N__16563,N__13329,N__16815,N__15414,N__15165,N__14931,N__13590}),
            .MASK({dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873}),
            .WDATA({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,N__6440,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,N__6325,dangling_wire_885,dangling_wire_886,dangling_wire_887}),
            .RCLKE(),
            .RCLK(N__17396),
            .RE(N__12594),
            .WCLKE(),
            .WCLK(N__16120),
            .WE(N__12160));
    defparam \line_buffer.mem13_physical .WRITE_MODE=3;
    defparam \line_buffer.mem13_physical .READ_MODE=3;
    defparam \line_buffer.mem13_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem13_physical  (
            .RDATA({dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,\line_buffer.n681 ,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,\line_buffer.n680 ,dangling_wire_899,dangling_wire_900,dangling_wire_901}),
            .RADDR({N__10533,N__11067,N__10794,N__11724,N__9822,N__9543,N__9279,N__11448,N__9015,N__12003,N__13989}),
            .WADDR({N__16296,N__14691,N__12930,N__13182,N__16659,N__13425,N__16911,N__15510,N__15261,N__15027,N__13686}),
            .MASK({dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917}),
            .WDATA({dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,N__6191,dangling_wire_922,dangling_wire_923,dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,dangling_wire_928,N__6881,dangling_wire_929,dangling_wire_930,dangling_wire_931}),
            .RCLKE(),
            .RCLK(N__17558),
            .RE(N__12470),
            .WCLKE(),
            .WCLK(N__16099),
            .WE(N__18184));
    defparam \line_buffer.mem19_physical .WRITE_MODE=3;
    defparam \line_buffer.mem19_physical .READ_MODE=3;
    defparam \line_buffer.mem19_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem19_physical  (
            .RDATA({dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,\line_buffer.n624 ,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,\line_buffer.n623 ,dangling_wire_943,dangling_wire_944,dangling_wire_945}),
            .RADDR({N__10461,N__10995,N__10722,N__11652,N__9750,N__9471,N__9207,N__11376,N__8943,N__11931,N__13917}),
            .WADDR({N__16224,N__14619,N__12858,N__13110,N__16587,N__13353,N__16839,N__15438,N__15189,N__14955,N__13614}),
            .MASK({dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961}),
            .WDATA({dangling_wire_962,dangling_wire_963,dangling_wire_964,dangling_wire_965,N__6205,dangling_wire_966,dangling_wire_967,dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,dangling_wire_972,N__6900,dangling_wire_973,dangling_wire_974,dangling_wire_975}),
            .RCLKE(),
            .RCLK(N__17311),
            .RE(N__12568),
            .WCLKE(),
            .WCLK(N__16113),
            .WE(N__17736));
    defparam \line_buffer.mem23_physical .WRITE_MODE=3;
    defparam \line_buffer.mem23_physical .READ_MODE=3;
    defparam \line_buffer.mem23_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem23_physical  (
            .RDATA({dangling_wire_976,dangling_wire_977,dangling_wire_978,dangling_wire_979,\line_buffer.n693 ,dangling_wire_980,dangling_wire_981,dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,\line_buffer.n692 ,dangling_wire_987,dangling_wire_988,dangling_wire_989}),
            .RADDR({N__10597,N__11128,N__10845,N__11791,N__9883,N__9600,N__9336,N__11509,N__9060,N__12064,N__14050}),
            .WADDR({N__16353,N__14748,N__12987,N__13227,N__16716,N__13486,N__16962,N__15567,N__15325,N__15084,N__13747}),
            .MASK({dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997,dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005}),
            .WDATA({dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,dangling_wire_1009,N__6402,dangling_wire_1010,dangling_wire_1011,dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,dangling_wire_1016,N__6251,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019}),
            .RCLKE(),
            .RCLK(N__17588),
            .RE(N__12451),
            .WCLKE(),
            .WCLK(N__16079),
            .WE(N__6994));
    defparam \line_buffer.mem0_physical .WRITE_MODE=3;
    defparam \line_buffer.mem0_physical .READ_MODE=3;
    defparam \line_buffer.mem0_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem0_physical  (
            .RDATA({dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,dangling_wire_1023,\line_buffer.n687 ,dangling_wire_1024,dangling_wire_1025,dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,\line_buffer.n686 ,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033}),
            .RADDR({N__10593,N__11127,N__10849,N__11784,N__9882,N__9601,N__9337,N__11508,N__9067,N__12063,N__14049}),
            .WADDR({N__16354,N__14749,N__12988,N__13234,N__16717,N__13485,N__16966,N__15568,N__15321,N__15085,N__13746}),
            .MASK({dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041,dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049}),
            .WDATA({dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,dangling_wire_1053,N__6468,dangling_wire_1054,dangling_wire_1055,dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,dangling_wire_1060,N__6607,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063}),
            .RCLKE(),
            .RCLK(N__17590),
            .RE(N__12407),
            .WCLKE(),
            .WCLK(N__16078),
            .WE(N__18199));
    defparam \line_buffer.mem26_physical .WRITE_MODE=3;
    defparam \line_buffer.mem26_physical .READ_MODE=3;
    defparam \line_buffer.mem26_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem26_physical  (
            .RDATA({dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,dangling_wire_1067,\line_buffer.n725 ,dangling_wire_1068,dangling_wire_1069,dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,\line_buffer.n724 ,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077}),
            .RADDR({N__10566,N__11094,N__10809,N__11763,N__9849,N__9564,N__9300,N__11475,N__9024,N__12030,N__14016}),
            .WADDR({N__16317,N__14712,N__12951,N__13191,N__16680,N__13452,N__16926,N__15531,N__15294,N__15048,N__13713}),
            .MASK({dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085,dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093}),
            .WDATA({dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,dangling_wire_1097,N__6388,dangling_wire_1098,dangling_wire_1099,dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,dangling_wire_1104,N__6276,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107}),
            .RCLKE(),
            .RCLK(N__17327),
            .RE(N__12521),
            .WCLKE(),
            .WCLK(N__16091),
            .WE(N__6795));
    defparam \line_buffer.mem3_physical .WRITE_MODE=3;
    defparam \line_buffer.mem3_physical .READ_MODE=3;
    defparam \line_buffer.mem3_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem3_physical  (
            .RDATA({dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,dangling_wire_1111,\line_buffer.n751 ,dangling_wire_1112,dangling_wire_1113,dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,\line_buffer.n750 ,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121}),
            .RADDR({N__10518,N__11046,N__10761,N__11715,N__9801,N__9516,N__9252,N__11427,N__8976,N__11982,N__13968}),
            .WADDR({N__16269,N__14664,N__12903,N__13143,N__16632,N__13404,N__16878,N__15483,N__15246,N__15000,N__13665}),
            .MASK({dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129,dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137}),
            .WDATA({dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,dangling_wire_1141,N__6522,dangling_wire_1142,dangling_wire_1143,dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,dangling_wire_1148,N__6626,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151}),
            .RCLKE(),
            .RCLK(N__17529),
            .RE(N__12579),
            .WCLKE(),
            .WCLK(N__16106),
            .WE(N__12165));
    defparam \line_buffer.mem17_physical .WRITE_MODE=3;
    defparam \line_buffer.mem17_physical .READ_MODE=3;
    defparam \line_buffer.mem17_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem17_physical  (
            .RDATA({dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,dangling_wire_1155,\line_buffer.n628 ,dangling_wire_1156,dangling_wire_1157,dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,\line_buffer.n627 ,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165}),
            .RADDR({N__10485,N__11019,N__10746,N__11676,N__9774,N__9495,N__9231,N__11400,N__8967,N__11955,N__13941}),
            .WADDR({N__16248,N__14643,N__12882,N__13134,N__16611,N__13377,N__16863,N__15462,N__15213,N__14979,N__13638}),
            .MASK({dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173,dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181}),
            .WDATA({dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,dangling_wire_1185,N__6441,dangling_wire_1186,dangling_wire_1187,dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,dangling_wire_1192,N__6314,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195}),
            .RCLKE(),
            .RCLK(N__17498),
            .RE(N__12538),
            .WCLKE(),
            .WCLK(N__16109),
            .WE(N__17712));
    defparam \line_buffer.mem31_physical .WRITE_MODE=3;
    defparam \line_buffer.mem31_physical .READ_MODE=3;
    defparam \line_buffer.mem31_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem31_physical  (
            .RDATA({dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,dangling_wire_1199,\line_buffer.n753 ,dangling_wire_1200,dangling_wire_1201,dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,\line_buffer.n752 ,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209}),
            .RADDR({N__10494,N__11022,N__10737,N__11691,N__9777,N__9492,N__9228,N__11403,N__8952,N__11958,N__13944}),
            .WADDR({N__16245,N__14640,N__12879,N__13119,N__16608,N__13380,N__16854,N__15459,N__15222,N__14976,N__13641}),
            .MASK({dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217,dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225}),
            .WDATA({dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,dangling_wire_1229,N__6195,dangling_wire_1230,dangling_wire_1231,dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,dangling_wire_1236,N__6866,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239}),
            .RCLKE(),
            .RCLK(N__17241),
            .RE(N__12599),
            .WCLKE(),
            .WCLK(N__16110),
            .WE(N__6692));
    defparam \line_buffer.mem9_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .WRITE_MODE=3;
    defparam \line_buffer.mem9_physical .READ_MODE=3;
    defparam \line_buffer.mem9_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem9_physical  (
            .RDATA({dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,dangling_wire_1243,\line_buffer.n618 ,dangling_wire_1244,dangling_wire_1245,dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,\line_buffer.n617 ,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253}),
            .RADDR({N__10422,N__10950,N__10665,N__11619,N__9705,N__9420,N__9156,N__11331,N__8880,N__11886,N__13872}),
            .WADDR({N__16173,N__14568,N__12807,N__13047,N__16536,N__13308,N__16782,N__15387,N__15150,N__14904,N__13569}),
            .MASK({dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261,dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269}),
            .WDATA({dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,dangling_wire_1273,N__6111,dangling_wire_1274,dangling_wire_1275,dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,dangling_wire_1280,N__6001,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283}),
            .RCLKE(),
            .RCLK(N__17151),
            .RE(N__12631),
            .WCLKE(),
            .WCLK(N__16125),
            .WE(N__6747));
    defparam \line_buffer.mem29_physical .WRITE_MODE=3;
    defparam \line_buffer.mem29_physical .READ_MODE=3;
    defparam \line_buffer.mem29_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem29_physical  (
            .RDATA({dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,dangling_wire_1287,\line_buffer.n757 ,dangling_wire_1288,dangling_wire_1289,dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,\line_buffer.n756 ,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297}),
            .RADDR({N__10530,N__11058,N__10773,N__11727,N__9813,N__9528,N__9264,N__11439,N__8988,N__11994,N__13980}),
            .WADDR({N__16281,N__14676,N__12915,N__13155,N__16644,N__13416,N__16890,N__15495,N__15258,N__15012,N__13677}),
            .MASK({dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305,dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313}),
            .WDATA({dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,dangling_wire_1317,N__6436,dangling_wire_1318,dangling_wire_1319,dangling_wire_1320,dangling_wire_1321,dangling_wire_1322,dangling_wire_1323,dangling_wire_1324,N__6289,dangling_wire_1325,dangling_wire_1326,dangling_wire_1327}),
            .RCLKE(),
            .RCLK(N__17518),
            .RE(N__12554),
            .WCLKE(),
            .WCLK(N__16104),
            .WE(N__6696));
    defparam \line_buffer.mem6_physical .WRITE_MODE=3;
    defparam \line_buffer.mem6_physical .READ_MODE=3;
    defparam \line_buffer.mem6_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem6_physical  (
            .RDATA({dangling_wire_1328,dangling_wire_1329,dangling_wire_1330,dangling_wire_1331,\line_buffer.n759 ,dangling_wire_1332,dangling_wire_1333,dangling_wire_1334,dangling_wire_1335,dangling_wire_1336,dangling_wire_1337,dangling_wire_1338,\line_buffer.n758 ,dangling_wire_1339,dangling_wire_1340,dangling_wire_1341}),
            .RADDR({N__10458,N__10986,N__10701,N__11655,N__9741,N__9456,N__9192,N__11367,N__8916,N__11922,N__13908}),
            .WADDR({N__16209,N__14604,N__12843,N__13083,N__16572,N__13344,N__16818,N__15423,N__15186,N__14940,N__13605}),
            .MASK({dangling_wire_1342,dangling_wire_1343,dangling_wire_1344,dangling_wire_1345,dangling_wire_1346,dangling_wire_1347,dangling_wire_1348,dangling_wire_1349,dangling_wire_1350,dangling_wire_1351,dangling_wire_1352,dangling_wire_1353,dangling_wire_1354,dangling_wire_1355,dangling_wire_1356,dangling_wire_1357}),
            .WDATA({dangling_wire_1358,dangling_wire_1359,dangling_wire_1360,dangling_wire_1361,N__6543,dangling_wire_1362,dangling_wire_1363,dangling_wire_1364,dangling_wire_1365,dangling_wire_1366,dangling_wire_1367,dangling_wire_1368,N__6654,dangling_wire_1369,dangling_wire_1370,dangling_wire_1371}),
            .RCLKE(),
            .RCLK(N__17328),
            .RE(N__12616),
            .WCLKE(),
            .WCLK(N__16119),
            .WE(N__6700));
    defparam \line_buffer.mem10_physical .WRITE_MODE=3;
    defparam \line_buffer.mem10_physical .READ_MODE=3;
    defparam \line_buffer.mem10_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem10_physical  (
            .RDATA({dangling_wire_1372,dangling_wire_1373,dangling_wire_1374,dangling_wire_1375,\line_buffer.n616 ,dangling_wire_1376,dangling_wire_1377,dangling_wire_1378,dangling_wire_1379,dangling_wire_1380,dangling_wire_1381,dangling_wire_1382,\line_buffer.n615 ,dangling_wire_1383,dangling_wire_1384,dangling_wire_1385}),
            .RADDR({N__10569,N__11103,N__10830,N__11760,N__9858,N__9579,N__9315,N__11484,N__9051,N__12039,N__14025}),
            .WADDR({N__16332,N__14727,N__12966,N__13218,N__16695,N__13461,N__16947,N__15546,N__15297,N__15063,N__13722}),
            .MASK({dangling_wire_1386,dangling_wire_1387,dangling_wire_1388,dangling_wire_1389,dangling_wire_1390,dangling_wire_1391,dangling_wire_1392,dangling_wire_1393,dangling_wire_1394,dangling_wire_1395,dangling_wire_1396,dangling_wire_1397,dangling_wire_1398,dangling_wire_1399,dangling_wire_1400,dangling_wire_1401}),
            .WDATA({dangling_wire_1402,dangling_wire_1403,dangling_wire_1404,dangling_wire_1405,N__6215,dangling_wire_1406,dangling_wire_1407,dangling_wire_1408,dangling_wire_1409,dangling_wire_1410,dangling_wire_1411,dangling_wire_1412,N__6867,dangling_wire_1413,dangling_wire_1414,dangling_wire_1415}),
            .RCLKE(),
            .RCLK(N__17580),
            .RE(N__12409),
            .WCLKE(),
            .WCLK(N__16085),
            .WE(N__6751));
    PRE_IO_GBUF TVP_CLK_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__18941),
            .GLOBALBUFFEROUTPUT(TVP_CLK_c));
    defparam TVP_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_CLK_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_CLK_pad_iopad (
            .OE(N__18943),
            .DIN(N__18942),
            .DOUT(N__18941),
            .PACKAGEPIN(TVP_CLK));
    defparam TVP_CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_CLK_pad_preio (
            .PADOEN(N__18943),
            .PADOUT(N__18942),
            .PADIN(N__18941),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_CLK_pad_iopad (
            .OE(N__18932),
            .DIN(N__18931),
            .DOUT(N__18930),
            .PACKAGEPIN(ADV_CLK));
    defparam ADV_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_CLK_pad_preio (
            .PADOEN(N__18932),
            .PADOUT(N__18931),
            .PADIN(N__18930),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17312),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_3_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_3_iopad (
            .OE(N__18923),
            .DIN(N__18922),
            .DOUT(N__18921),
            .PACKAGEPIN(DEBUG[3]));
    defparam DEBUG_pad_3_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_3_preio (
            .PADOEN(N__18923),
            .PADOUT(N__18922),
            .PADIN(N__18921),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11557),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_2_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_2_iopad (
            .OE(N__18914),
            .DIN(N__18913),
            .DOUT(N__18912),
            .PACKAGEPIN(TVP_VIDEO[2]));
    defparam TVP_VIDEO_pad_2_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_2_preio (
            .PADOEN(N__18914),
            .PADOUT(N__18913),
            .PADIN(N__18912),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_5_iopad (
            .OE(N__18905),
            .DIN(N__18904),
            .DOUT(N__18903),
            .PACKAGEPIN(ADV_G[5]));
    defparam ADV_G_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_5_preio (
            .PADOEN(N__18905),
            .PADOUT(N__18904),
            .PADIN(N__18903),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10311),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_3_iopad (
            .OE(N__18896),
            .DIN(N__18895),
            .DOUT(N__18894),
            .PACKAGEPIN(ADV_B[3]));
    defparam ADV_B_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_3_preio (
            .PADOEN(N__18896),
            .PADOUT(N__18895),
            .PADIN(N__18894),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10197),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_4_iopad (
            .OE(N__18887),
            .DIN(N__18886),
            .DOUT(N__18885),
            .PACKAGEPIN(ADV_R[4]));
    defparam ADV_R_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_4_preio (
            .PADOEN(N__18887),
            .PADOUT(N__18886),
            .PADIN(N__18885),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10127),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_8_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_8_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_8_iopad (
            .OE(N__18878),
            .DIN(N__18877),
            .DOUT(N__18876),
            .PACKAGEPIN(TVP_VIDEO[8]));
    defparam TVP_VIDEO_pad_8_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_8_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_8_preio (
            .PADOEN(N__18878),
            .PADOUT(N__18877),
            .PADIN(N__18876),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_0_iopad (
            .OE(N__18869),
            .DIN(N__18868),
            .DOUT(N__18867),
            .PACKAGEPIN(ADV_B[0]));
    defparam ADV_B_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_0_preio (
            .PADOEN(N__18869),
            .PADOUT(N__18868),
            .PADIN(N__18867),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8502),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_5_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_5_iopad (
            .OE(N__18860),
            .DIN(N__18859),
            .DOUT(N__18858),
            .PACKAGEPIN(TVP_VIDEO[5]));
    defparam TVP_VIDEO_pad_5_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_5_preio (
            .PADOEN(N__18860),
            .PADOUT(N__18859),
            .PADIN(N__18858),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_2_iopad (
            .OE(N__18851),
            .DIN(N__18850),
            .DOUT(N__18849),
            .PACKAGEPIN(ADV_G[2]));
    defparam ADV_G_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_2_preio (
            .PADOEN(N__18851),
            .PADOUT(N__18850),
            .PADIN(N__18849),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8433),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_VSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_VSYNC_pad_iopad (
            .OE(N__18842),
            .DIN(N__18841),
            .DOUT(N__18840),
            .PACKAGEPIN(ADV_VSYNC));
    defparam ADV_VSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_VSYNC_pad_preio (
            .PADOEN(N__18842),
            .PADOUT(N__18841),
            .PADIN(N__18840),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14452),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_3_iopad (
            .OE(N__18833),
            .DIN(N__18832),
            .DOUT(N__18831),
            .PACKAGEPIN(ADV_R[3]));
    defparam ADV_R_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_3_preio (
            .PADOEN(N__18833),
            .PADOUT(N__18832),
            .PADIN(N__18831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10196),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_5_iopad (
            .OE(N__18824),
            .DIN(N__18823),
            .DOUT(N__18822),
            .PACKAGEPIN(ADV_B[5]));
    defparam ADV_B_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_5_preio (
            .PADOEN(N__18824),
            .PADOUT(N__18823),
            .PADIN(N__18822),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10310),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_7_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_7_iopad (
            .OE(N__18815),
            .DIN(N__18814),
            .DOUT(N__18813),
            .PACKAGEPIN(DEBUG[7]));
    defparam DEBUG_pad_7_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_7_preio (
            .PADOEN(N__18815),
            .PADOUT(N__18814),
            .PADIN(N__18813),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11851),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_6_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_6_iopad (
            .OE(N__18806),
            .DIN(N__18805),
            .DOUT(N__18804),
            .PACKAGEPIN(TVP_VIDEO[6]));
    defparam TVP_VIDEO_pad_6_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_6_preio (
            .PADOEN(N__18806),
            .PADOUT(N__18805),
            .PADIN(N__18804),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_1_iopad (
            .OE(N__18797),
            .DIN(N__18796),
            .DOUT(N__18795),
            .PACKAGEPIN(ADV_G[1]));
    defparam ADV_G_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_1_preio (
            .PADOEN(N__18797),
            .PADOUT(N__18796),
            .PADIN(N__18795),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10264),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_0_iopad (
            .OE(N__18788),
            .DIN(N__18787),
            .DOUT(N__18786),
            .PACKAGEPIN(ADV_R[0]));
    defparam ADV_R_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_0_preio (
            .PADOEN(N__18788),
            .PADOUT(N__18787),
            .PADIN(N__18786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8498),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_2_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_2_iopad (
            .OE(N__18779),
            .DIN(N__18778),
            .DOUT(N__18777),
            .PACKAGEPIN(DEBUG[2]));
    defparam DEBUG_pad_2_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_2_preio (
            .PADOEN(N__18779),
            .PADOUT(N__18778),
            .PADIN(N__18777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9112),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_3_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_3_iopad (
            .OE(N__18770),
            .DIN(N__18769),
            .DOUT(N__18768),
            .PACKAGEPIN(TVP_VIDEO[3]));
    defparam TVP_VIDEO_pad_3_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_3_preio (
            .PADOEN(N__18770),
            .PADOUT(N__18769),
            .PADIN(N__18768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_4_iopad (
            .OE(N__18761),
            .DIN(N__18760),
            .DOUT(N__18759),
            .PACKAGEPIN(ADV_G[4]));
    defparam ADV_G_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_4_preio (
            .PADOEN(N__18761),
            .PADOUT(N__18760),
            .PADIN(N__18759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10138),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_5_iopad (
            .OE(N__18752),
            .DIN(N__18751),
            .DOUT(N__18750),
            .PACKAGEPIN(ADV_R[5]));
    defparam ADV_R_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_5_preio (
            .PADOEN(N__18752),
            .PADOUT(N__18751),
            .PADIN(N__18750),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10318),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_9_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_9_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_9_iopad (
            .OE(N__18743),
            .DIN(N__18742),
            .DOUT(N__18741),
            .PACKAGEPIN(TVP_VIDEO[9]));
    defparam TVP_VIDEO_pad_9_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_9_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_9_preio (
            .PADOEN(N__18743),
            .PADOUT(N__18742),
            .PADIN(N__18741),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_3_iopad (
            .OE(N__18734),
            .DIN(N__18733),
            .DOUT(N__18732),
            .PACKAGEPIN(ADV_G[3]));
    defparam ADV_G_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_3_preio (
            .PADOEN(N__18734),
            .PADOUT(N__18733),
            .PADIN(N__18732),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10198),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_HSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_HSYNC_pad_iopad (
            .OE(N__18725),
            .DIN(N__18724),
            .DOUT(N__18723),
            .PACKAGEPIN(ADV_HSYNC));
    defparam ADV_HSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_HSYNC_pad_preio (
            .PADOEN(N__18725),
            .PADOUT(N__18724),
            .PADIN(N__18723),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7309),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_2_iopad (
            .OE(N__18716),
            .DIN(N__18715),
            .DOUT(N__18714),
            .PACKAGEPIN(ADV_R[2]));
    defparam ADV_R_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_2_preio (
            .PADOEN(N__18716),
            .PADOUT(N__18715),
            .PADIN(N__18714),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8429),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_1_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_1_iopad (
            .OE(N__18707),
            .DIN(N__18706),
            .DOUT(N__18705),
            .PACKAGEPIN(DEBUG[1]));
    defparam DEBUG_pad_1_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_1_preio (
            .PADOEN(N__18707),
            .PADOUT(N__18706),
            .PADIN(N__18705),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12100),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_4_iopad (
            .OE(N__18698),
            .DIN(N__18697),
            .DOUT(N__18696),
            .PACKAGEPIN(ADV_B[4]));
    defparam ADV_B_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_4_preio (
            .PADOEN(N__18698),
            .PADOUT(N__18697),
            .PADIN(N__18696),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10137),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_4_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_4_iopad (
            .OE(N__18689),
            .DIN(N__18688),
            .DOUT(N__18687),
            .PACKAGEPIN(DEBUG[4]));
    defparam DEBUG_pad_4_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_4_preio (
            .PADOEN(N__18689),
            .PADOUT(N__18688),
            .PADIN(N__18687),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9370),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_1_iopad (
            .OE(N__18680),
            .DIN(N__18679),
            .DOUT(N__18678),
            .PACKAGEPIN(ADV_B[1]));
    defparam ADV_B_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_1_preio (
            .PADOEN(N__18680),
            .PADOUT(N__18679),
            .PADIN(N__18678),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10256),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_6_iopad (
            .OE(N__18671),
            .DIN(N__18670),
            .DOUT(N__18669),
            .PACKAGEPIN(ADV_G[6]));
    defparam ADV_G_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_6_preio (
            .PADOEN(N__18671),
            .PADOUT(N__18670),
            .PADIN(N__18669),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10077),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_SYNC_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_SYNC_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_SYNC_N_pad_iopad (
            .OE(N__18662),
            .DIN(N__18661),
            .DOUT(N__18660),
            .PACKAGEPIN(ADV_SYNC_N));
    defparam ADV_SYNC_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_SYNC_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_SYNC_N_pad_preio (
            .PADOEN(N__18662),
            .PADOUT(N__18661),
            .PADIN(N__18660),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_7_iopad (
            .OE(N__18653),
            .DIN(N__18652),
            .DOUT(N__18651),
            .PACKAGEPIN(ADV_R[7]));
    defparam ADV_R_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_7_preio (
            .PADOEN(N__18653),
            .PADOUT(N__18652),
            .PADIN(N__18651),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10020),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_6_iopad (
            .OE(N__18644),
            .DIN(N__18643),
            .DOUT(N__18642),
            .PACKAGEPIN(ADV_B[6]));
    defparam ADV_B_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_6_preio (
            .PADOEN(N__18644),
            .PADOUT(N__18643),
            .PADIN(N__18642),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10076),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_6_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_6_iopad (
            .OE(N__18635),
            .DIN(N__18634),
            .DOUT(N__18633),
            .PACKAGEPIN(DEBUG[6]));
    defparam DEBUG_pad_6_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_6_preio (
            .PADOEN(N__18635),
            .PADOUT(N__18634),
            .PADIN(N__18633),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9934),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_7_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_7_iopad (
            .OE(N__18626),
            .DIN(N__18625),
            .DOUT(N__18624),
            .PACKAGEPIN(TVP_VIDEO[7]));
    defparam TVP_VIDEO_pad_7_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_7_preio (
            .PADOEN(N__18626),
            .PADOUT(N__18625),
            .PADIN(N__18624),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_0_iopad (
            .OE(N__18617),
            .DIN(N__18616),
            .DOUT(N__18615),
            .PACKAGEPIN(ADV_G[0]));
    defparam ADV_G_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_0_preio (
            .PADOEN(N__18617),
            .PADOUT(N__18616),
            .PADIN(N__18615),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8509),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_1_iopad (
            .OE(N__18608),
            .DIN(N__18607),
            .DOUT(N__18606),
            .PACKAGEPIN(ADV_R[1]));
    defparam ADV_R_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_1_preio (
            .PADOEN(N__18608),
            .PADOUT(N__18607),
            .PADIN(N__18606),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10257),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_5_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_5_iopad (
            .OE(N__18599),
            .DIN(N__18598),
            .DOUT(N__18597),
            .PACKAGEPIN(DEBUG[5]));
    defparam DEBUG_pad_5_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_5_preio (
            .PADOEN(N__18599),
            .PADOUT(N__18598),
            .PADIN(N__18597),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9643),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_HSYNC_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_HSYNC_pad_iopad (
            .OE(N__18590),
            .DIN(N__18589),
            .DOUT(N__18588),
            .PACKAGEPIN(TVP_HSYNC));
    defparam TVP_HSYNC_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_HSYNC_pad_preio (
            .PADOEN(N__18590),
            .PADOUT(N__18589),
            .PADIN(N__18588),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_HSYNC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_7_iopad (
            .OE(N__18581),
            .DIN(N__18580),
            .DOUT(N__18579),
            .PACKAGEPIN(ADV_G[7]));
    defparam ADV_G_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_7_preio (
            .PADOEN(N__18581),
            .PADOUT(N__18580),
            .PADIN(N__18579),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10019),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_6_iopad (
            .OE(N__18572),
            .DIN(N__18571),
            .DOUT(N__18570),
            .PACKAGEPIN(ADV_R[6]));
    defparam ADV_R_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_6_preio (
            .PADOEN(N__18572),
            .PADOUT(N__18571),
            .PADIN(N__18570),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10081),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VSYNC_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_VSYNC_pad_iopad (
            .OE(N__18563),
            .DIN(N__18562),
            .DOUT(N__18561),
            .PACKAGEPIN(TVP_VSYNC));
    defparam TVP_VSYNC_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VSYNC_pad_preio (
            .PADOEN(N__18563),
            .PADOUT(N__18562),
            .PADIN(N__18561),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VSYNC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_BLANK_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_BLANK_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_BLANK_N_pad_iopad (
            .OE(N__18554),
            .DIN(N__18553),
            .DOUT(N__18552),
            .PACKAGEPIN(ADV_BLANK_N));
    defparam ADV_BLANK_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_BLANK_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_BLANK_N_pad_preio (
            .PADOEN(N__18554),
            .PADOUT(N__18553),
            .PADIN(N__18552),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12537),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_0_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_0_iopad (
            .OE(N__18545),
            .DIN(N__18544),
            .DOUT(N__18543),
            .PACKAGEPIN(DEBUG[0]));
    defparam DEBUG_pad_0_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_0_preio (
            .PADOEN(N__18545),
            .PADOUT(N__18544),
            .PADIN(N__18543),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14233),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_2_iopad (
            .OE(N__18536),
            .DIN(N__18535),
            .DOUT(N__18534),
            .PACKAGEPIN(ADV_B[2]));
    defparam ADV_B_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_2_preio (
            .PADOEN(N__18536),
            .PADOUT(N__18535),
            .PADIN(N__18534),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8440),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_7_iopad (
            .OE(N__18527),
            .DIN(N__18526),
            .DOUT(N__18525),
            .PACKAGEPIN(ADV_B[7]));
    defparam ADV_B_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_7_preio (
            .PADOEN(N__18527),
            .PADOUT(N__18526),
            .PADIN(N__18525),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10021),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__18518),
            .DIN(N__18517),
            .DOUT(N__18516),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__18518),
            .PADOUT(N__18517),
            .PADIN(N__18516),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8803),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_4_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_4_iopad (
            .OE(N__18509),
            .DIN(N__18508),
            .DOUT(N__18507),
            .PACKAGEPIN(TVP_VIDEO[4]));
    defparam TVP_VIDEO_pad_4_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_4_preio (
            .PADOEN(N__18509),
            .PADOUT(N__18508),
            .PADIN(N__18507),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__4528 (
            .O(N__18490),
            .I(N__18484));
    InMux I__4527 (
            .O(N__18489),
            .I(N__18481));
    InMux I__4526 (
            .O(N__18488),
            .I(N__18478));
    InMux I__4525 (
            .O(N__18487),
            .I(N__18466));
    LocalMux I__4524 (
            .O(N__18484),
            .I(N__18461));
    LocalMux I__4523 (
            .O(N__18481),
            .I(N__18461));
    LocalMux I__4522 (
            .O(N__18478),
            .I(N__18458));
    InMux I__4521 (
            .O(N__18477),
            .I(N__18455));
    InMux I__4520 (
            .O(N__18476),
            .I(N__18452));
    InMux I__4519 (
            .O(N__18475),
            .I(N__18445));
    InMux I__4518 (
            .O(N__18474),
            .I(N__18442));
    InMux I__4517 (
            .O(N__18473),
            .I(N__18436));
    InMux I__4516 (
            .O(N__18472),
            .I(N__18433));
    InMux I__4515 (
            .O(N__18471),
            .I(N__18430));
    InMux I__4514 (
            .O(N__18470),
            .I(N__18427));
    InMux I__4513 (
            .O(N__18469),
            .I(N__18424));
    LocalMux I__4512 (
            .O(N__18466),
            .I(N__18421));
    Span4Mux_h I__4511 (
            .O(N__18461),
            .I(N__18412));
    Span4Mux_v I__4510 (
            .O(N__18458),
            .I(N__18412));
    LocalMux I__4509 (
            .O(N__18455),
            .I(N__18412));
    LocalMux I__4508 (
            .O(N__18452),
            .I(N__18412));
    InMux I__4507 (
            .O(N__18451),
            .I(N__18409));
    InMux I__4506 (
            .O(N__18450),
            .I(N__18406));
    InMux I__4505 (
            .O(N__18449),
            .I(N__18403));
    InMux I__4504 (
            .O(N__18448),
            .I(N__18400));
    LocalMux I__4503 (
            .O(N__18445),
            .I(N__18397));
    LocalMux I__4502 (
            .O(N__18442),
            .I(N__18394));
    InMux I__4501 (
            .O(N__18441),
            .I(N__18390));
    InMux I__4500 (
            .O(N__18440),
            .I(N__18387));
    InMux I__4499 (
            .O(N__18439),
            .I(N__18382));
    LocalMux I__4498 (
            .O(N__18436),
            .I(N__18379));
    LocalMux I__4497 (
            .O(N__18433),
            .I(N__18376));
    LocalMux I__4496 (
            .O(N__18430),
            .I(N__18373));
    LocalMux I__4495 (
            .O(N__18427),
            .I(N__18368));
    LocalMux I__4494 (
            .O(N__18424),
            .I(N__18368));
    Span4Mux_h I__4493 (
            .O(N__18421),
            .I(N__18363));
    Span4Mux_h I__4492 (
            .O(N__18412),
            .I(N__18363));
    LocalMux I__4491 (
            .O(N__18409),
            .I(N__18360));
    LocalMux I__4490 (
            .O(N__18406),
            .I(N__18351));
    LocalMux I__4489 (
            .O(N__18403),
            .I(N__18351));
    LocalMux I__4488 (
            .O(N__18400),
            .I(N__18351));
    Span4Mux_v I__4487 (
            .O(N__18397),
            .I(N__18351));
    Span4Mux_v I__4486 (
            .O(N__18394),
            .I(N__18348));
    InMux I__4485 (
            .O(N__18393),
            .I(N__18345));
    LocalMux I__4484 (
            .O(N__18390),
            .I(N__18342));
    LocalMux I__4483 (
            .O(N__18387),
            .I(N__18339));
    InMux I__4482 (
            .O(N__18386),
            .I(N__18336));
    InMux I__4481 (
            .O(N__18385),
            .I(N__18333));
    LocalMux I__4480 (
            .O(N__18382),
            .I(N__18330));
    Span12Mux_v I__4479 (
            .O(N__18379),
            .I(N__18327));
    Span12Mux_h I__4478 (
            .O(N__18376),
            .I(N__18322));
    Span12Mux_h I__4477 (
            .O(N__18373),
            .I(N__18322));
    Span4Mux_h I__4476 (
            .O(N__18368),
            .I(N__18317));
    Span4Mux_v I__4475 (
            .O(N__18363),
            .I(N__18317));
    Span4Mux_v I__4474 (
            .O(N__18360),
            .I(N__18310));
    Span4Mux_v I__4473 (
            .O(N__18351),
            .I(N__18310));
    Span4Mux_h I__4472 (
            .O(N__18348),
            .I(N__18310));
    LocalMux I__4471 (
            .O(N__18345),
            .I(N__18303));
    Span4Mux_v I__4470 (
            .O(N__18342),
            .I(N__18303));
    Span4Mux_v I__4469 (
            .O(N__18339),
            .I(N__18303));
    LocalMux I__4468 (
            .O(N__18336),
            .I(TX_ADDR_11));
    LocalMux I__4467 (
            .O(N__18333),
            .I(TX_ADDR_11));
    Odrv4 I__4466 (
            .O(N__18330),
            .I(TX_ADDR_11));
    Odrv12 I__4465 (
            .O(N__18327),
            .I(TX_ADDR_11));
    Odrv12 I__4464 (
            .O(N__18322),
            .I(TX_ADDR_11));
    Odrv4 I__4463 (
            .O(N__18317),
            .I(TX_ADDR_11));
    Odrv4 I__4462 (
            .O(N__18310),
            .I(TX_ADDR_11));
    Odrv4 I__4461 (
            .O(N__18303),
            .I(TX_ADDR_11));
    InMux I__4460 (
            .O(N__18286),
            .I(N__18283));
    LocalMux I__4459 (
            .O(N__18283),
            .I(N__18280));
    Span4Mux_v I__4458 (
            .O(N__18280),
            .I(N__18277));
    Sp12to4 I__4457 (
            .O(N__18277),
            .I(N__18274));
    Odrv12 I__4456 (
            .O(N__18274),
            .I(\line_buffer.n756 ));
    InMux I__4455 (
            .O(N__18271),
            .I(N__18268));
    LocalMux I__4454 (
            .O(N__18268),
            .I(N__18265));
    Span4Mux_v I__4453 (
            .O(N__18265),
            .I(N__18262));
    Span4Mux_v I__4452 (
            .O(N__18262),
            .I(N__18259));
    Span4Mux_v I__4451 (
            .O(N__18259),
            .I(N__18256));
    Span4Mux_h I__4450 (
            .O(N__18256),
            .I(N__18253));
    Odrv4 I__4449 (
            .O(N__18253),
            .I(\line_buffer.n748 ));
    InMux I__4448 (
            .O(N__18250),
            .I(N__18247));
    LocalMux I__4447 (
            .O(N__18247),
            .I(\line_buffer.n3025 ));
    SRMux I__4446 (
            .O(N__18244),
            .I(N__18240));
    SRMux I__4445 (
            .O(N__18243),
            .I(N__18237));
    LocalMux I__4444 (
            .O(N__18240),
            .I(N__18232));
    LocalMux I__4443 (
            .O(N__18237),
            .I(N__18229));
    SRMux I__4442 (
            .O(N__18236),
            .I(N__18226));
    SRMux I__4441 (
            .O(N__18235),
            .I(N__18223));
    Span4Mux_v I__4440 (
            .O(N__18232),
            .I(N__18220));
    Span4Mux_v I__4439 (
            .O(N__18229),
            .I(N__18213));
    LocalMux I__4438 (
            .O(N__18226),
            .I(N__18213));
    LocalMux I__4437 (
            .O(N__18223),
            .I(N__18213));
    Span4Mux_v I__4436 (
            .O(N__18220),
            .I(N__18210));
    Span4Mux_v I__4435 (
            .O(N__18213),
            .I(N__18207));
    Span4Mux_v I__4434 (
            .O(N__18210),
            .I(N__18202));
    Span4Mux_h I__4433 (
            .O(N__18207),
            .I(N__18202));
    Odrv4 I__4432 (
            .O(N__18202),
            .I(\line_buffer.n729 ));
    SRMux I__4431 (
            .O(N__18199),
            .I(N__18196));
    LocalMux I__4430 (
            .O(N__18196),
            .I(N__18193));
    Span4Mux_s3_v I__4429 (
            .O(N__18193),
            .I(N__18188));
    SRMux I__4428 (
            .O(N__18192),
            .I(N__18185));
    SRMux I__4427 (
            .O(N__18191),
            .I(N__18181));
    Span4Mux_v I__4426 (
            .O(N__18188),
            .I(N__18176));
    LocalMux I__4425 (
            .O(N__18185),
            .I(N__18176));
    SRMux I__4424 (
            .O(N__18184),
            .I(N__18173));
    LocalMux I__4423 (
            .O(N__18181),
            .I(N__18170));
    Span4Mux_h I__4422 (
            .O(N__18176),
            .I(N__18167));
    LocalMux I__4421 (
            .O(N__18173),
            .I(N__18164));
    Span4Mux_h I__4420 (
            .O(N__18170),
            .I(N__18161));
    Span4Mux_v I__4419 (
            .O(N__18167),
            .I(N__18156));
    Span4Mux_h I__4418 (
            .O(N__18164),
            .I(N__18156));
    Odrv4 I__4417 (
            .O(N__18161),
            .I(\line_buffer.n697 ));
    Odrv4 I__4416 (
            .O(N__18156),
            .I(\line_buffer.n697 ));
    InMux I__4415 (
            .O(N__18151),
            .I(N__18146));
    InMux I__4414 (
            .O(N__18150),
            .I(N__18143));
    CascadeMux I__4413 (
            .O(N__18149),
            .I(N__18140));
    LocalMux I__4412 (
            .O(N__18146),
            .I(N__18130));
    LocalMux I__4411 (
            .O(N__18143),
            .I(N__18130));
    InMux I__4410 (
            .O(N__18140),
            .I(N__18125));
    InMux I__4409 (
            .O(N__18139),
            .I(N__18125));
    InMux I__4408 (
            .O(N__18138),
            .I(N__18122));
    InMux I__4407 (
            .O(N__18137),
            .I(N__18119));
    InMux I__4406 (
            .O(N__18136),
            .I(N__18116));
    InMux I__4405 (
            .O(N__18135),
            .I(N__18113));
    Span4Mux_v I__4404 (
            .O(N__18130),
            .I(N__18108));
    LocalMux I__4403 (
            .O(N__18125),
            .I(N__18108));
    LocalMux I__4402 (
            .O(N__18122),
            .I(N__18104));
    LocalMux I__4401 (
            .O(N__18119),
            .I(N__18101));
    LocalMux I__4400 (
            .O(N__18116),
            .I(N__18098));
    LocalMux I__4399 (
            .O(N__18113),
            .I(N__18095));
    Sp12to4 I__4398 (
            .O(N__18108),
            .I(N__18092));
    InMux I__4397 (
            .O(N__18107),
            .I(N__18089));
    Span4Mux_v I__4396 (
            .O(N__18104),
            .I(N__18084));
    Span4Mux_v I__4395 (
            .O(N__18101),
            .I(N__18084));
    Span12Mux_v I__4394 (
            .O(N__18098),
            .I(N__18077));
    Span12Mux_v I__4393 (
            .O(N__18095),
            .I(N__18077));
    Span12Mux_v I__4392 (
            .O(N__18092),
            .I(N__18077));
    LocalMux I__4391 (
            .O(N__18089),
            .I(RX_ADDR_12));
    Odrv4 I__4390 (
            .O(N__18084),
            .I(RX_ADDR_12));
    Odrv12 I__4389 (
            .O(N__18077),
            .I(RX_ADDR_12));
    InMux I__4388 (
            .O(N__18070),
            .I(N__18064));
    InMux I__4387 (
            .O(N__18069),
            .I(N__18059));
    InMux I__4386 (
            .O(N__18068),
            .I(N__18059));
    InMux I__4385 (
            .O(N__18067),
            .I(N__18056));
    LocalMux I__4384 (
            .O(N__18064),
            .I(N__18051));
    LocalMux I__4383 (
            .O(N__18059),
            .I(N__18048));
    LocalMux I__4382 (
            .O(N__18056),
            .I(N__18043));
    InMux I__4381 (
            .O(N__18055),
            .I(N__18040));
    InMux I__4380 (
            .O(N__18054),
            .I(N__18037));
    Span4Mux_v I__4379 (
            .O(N__18051),
            .I(N__18032));
    Span4Mux_v I__4378 (
            .O(N__18048),
            .I(N__18032));
    InMux I__4377 (
            .O(N__18047),
            .I(N__18029));
    InMux I__4376 (
            .O(N__18046),
            .I(N__18026));
    Span4Mux_v I__4375 (
            .O(N__18043),
            .I(N__18023));
    LocalMux I__4374 (
            .O(N__18040),
            .I(N__18020));
    LocalMux I__4373 (
            .O(N__18037),
            .I(N__18017));
    Span4Mux_h I__4372 (
            .O(N__18032),
            .I(N__18014));
    LocalMux I__4371 (
            .O(N__18029),
            .I(N__18011));
    LocalMux I__4370 (
            .O(N__18026),
            .I(N__18008));
    Span4Mux_h I__4369 (
            .O(N__18023),
            .I(N__18004));
    Span4Mux_v I__4368 (
            .O(N__18020),
            .I(N__17999));
    Span4Mux_v I__4367 (
            .O(N__18017),
            .I(N__17999));
    Span4Mux_h I__4366 (
            .O(N__18014),
            .I(N__17992));
    Span4Mux_v I__4365 (
            .O(N__18011),
            .I(N__17992));
    Span4Mux_v I__4364 (
            .O(N__18008),
            .I(N__17992));
    InMux I__4363 (
            .O(N__18007),
            .I(N__17989));
    Odrv4 I__4362 (
            .O(N__18004),
            .I(RX_ADDR_11));
    Odrv4 I__4361 (
            .O(N__17999),
            .I(RX_ADDR_11));
    Odrv4 I__4360 (
            .O(N__17992),
            .I(RX_ADDR_11));
    LocalMux I__4359 (
            .O(N__17989),
            .I(RX_ADDR_11));
    CascadeMux I__4358 (
            .O(N__17980),
            .I(N__17976));
    CascadeMux I__4357 (
            .O(N__17979),
            .I(N__17968));
    InMux I__4356 (
            .O(N__17976),
            .I(N__17965));
    CascadeMux I__4355 (
            .O(N__17975),
            .I(N__17962));
    CascadeMux I__4354 (
            .O(N__17974),
            .I(N__17959));
    CascadeMux I__4353 (
            .O(N__17973),
            .I(N__17956));
    CascadeMux I__4352 (
            .O(N__17972),
            .I(N__17953));
    CascadeMux I__4351 (
            .O(N__17971),
            .I(N__17949));
    InMux I__4350 (
            .O(N__17968),
            .I(N__17946));
    LocalMux I__4349 (
            .O(N__17965),
            .I(N__17943));
    InMux I__4348 (
            .O(N__17962),
            .I(N__17940));
    InMux I__4347 (
            .O(N__17959),
            .I(N__17937));
    InMux I__4346 (
            .O(N__17956),
            .I(N__17934));
    InMux I__4345 (
            .O(N__17953),
            .I(N__17931));
    InMux I__4344 (
            .O(N__17952),
            .I(N__17926));
    InMux I__4343 (
            .O(N__17949),
            .I(N__17926));
    LocalMux I__4342 (
            .O(N__17946),
            .I(N__17922));
    Span4Mux_h I__4341 (
            .O(N__17943),
            .I(N__17919));
    LocalMux I__4340 (
            .O(N__17940),
            .I(N__17916));
    LocalMux I__4339 (
            .O(N__17937),
            .I(N__17911));
    LocalMux I__4338 (
            .O(N__17934),
            .I(N__17911));
    LocalMux I__4337 (
            .O(N__17931),
            .I(N__17908));
    LocalMux I__4336 (
            .O(N__17926),
            .I(N__17905));
    InMux I__4335 (
            .O(N__17925),
            .I(N__17902));
    Span4Mux_v I__4334 (
            .O(N__17922),
            .I(N__17897));
    Span4Mux_h I__4333 (
            .O(N__17919),
            .I(N__17897));
    Span4Mux_h I__4332 (
            .O(N__17916),
            .I(N__17892));
    Span4Mux_h I__4331 (
            .O(N__17911),
            .I(N__17892));
    Span12Mux_v I__4330 (
            .O(N__17908),
            .I(N__17887));
    Span12Mux_v I__4329 (
            .O(N__17905),
            .I(N__17887));
    LocalMux I__4328 (
            .O(N__17902),
            .I(RX_ADDR_13));
    Odrv4 I__4327 (
            .O(N__17897),
            .I(RX_ADDR_13));
    Odrv4 I__4326 (
            .O(N__17892),
            .I(RX_ADDR_13));
    Odrv12 I__4325 (
            .O(N__17887),
            .I(RX_ADDR_13));
    InMux I__4324 (
            .O(N__17878),
            .I(N__17862));
    InMux I__4323 (
            .O(N__17877),
            .I(N__17858));
    InMux I__4322 (
            .O(N__17876),
            .I(N__17854));
    InMux I__4321 (
            .O(N__17875),
            .I(N__17851));
    InMux I__4320 (
            .O(N__17874),
            .I(N__17846));
    InMux I__4319 (
            .O(N__17873),
            .I(N__17846));
    InMux I__4318 (
            .O(N__17872),
            .I(N__17839));
    InMux I__4317 (
            .O(N__17871),
            .I(N__17839));
    InMux I__4316 (
            .O(N__17870),
            .I(N__17839));
    InMux I__4315 (
            .O(N__17869),
            .I(N__17828));
    InMux I__4314 (
            .O(N__17868),
            .I(N__17828));
    InMux I__4313 (
            .O(N__17867),
            .I(N__17828));
    InMux I__4312 (
            .O(N__17866),
            .I(N__17828));
    InMux I__4311 (
            .O(N__17865),
            .I(N__17828));
    LocalMux I__4310 (
            .O(N__17862),
            .I(N__17825));
    InMux I__4309 (
            .O(N__17861),
            .I(N__17822));
    LocalMux I__4308 (
            .O(N__17858),
            .I(N__17819));
    InMux I__4307 (
            .O(N__17857),
            .I(N__17816));
    LocalMux I__4306 (
            .O(N__17854),
            .I(N__17813));
    LocalMux I__4305 (
            .O(N__17851),
            .I(N__17806));
    LocalMux I__4304 (
            .O(N__17846),
            .I(N__17806));
    LocalMux I__4303 (
            .O(N__17839),
            .I(N__17803));
    LocalMux I__4302 (
            .O(N__17828),
            .I(N__17796));
    Span4Mux_v I__4301 (
            .O(N__17825),
            .I(N__17796));
    LocalMux I__4300 (
            .O(N__17822),
            .I(N__17796));
    Span4Mux_h I__4299 (
            .O(N__17819),
            .I(N__17789));
    LocalMux I__4298 (
            .O(N__17816),
            .I(N__17789));
    Span4Mux_v I__4297 (
            .O(N__17813),
            .I(N__17789));
    InMux I__4296 (
            .O(N__17812),
            .I(N__17784));
    InMux I__4295 (
            .O(N__17811),
            .I(N__17784));
    Span4Mux_v I__4294 (
            .O(N__17806),
            .I(N__17781));
    Span4Mux_v I__4293 (
            .O(N__17803),
            .I(N__17777));
    Span4Mux_v I__4292 (
            .O(N__17796),
            .I(N__17772));
    Span4Mux_h I__4291 (
            .O(N__17789),
            .I(N__17772));
    LocalMux I__4290 (
            .O(N__17784),
            .I(N__17769));
    Span4Mux_h I__4289 (
            .O(N__17781),
            .I(N__17766));
    InMux I__4288 (
            .O(N__17780),
            .I(N__17763));
    Span4Mux_h I__4287 (
            .O(N__17777),
            .I(N__17759));
    Span4Mux_h I__4286 (
            .O(N__17772),
            .I(N__17754));
    Span4Mux_v I__4285 (
            .O(N__17769),
            .I(N__17754));
    Span4Mux_h I__4284 (
            .O(N__17766),
            .I(N__17749));
    LocalMux I__4283 (
            .O(N__17763),
            .I(N__17749));
    InMux I__4282 (
            .O(N__17762),
            .I(N__17746));
    Odrv4 I__4281 (
            .O(N__17759),
            .I(n25));
    Odrv4 I__4280 (
            .O(N__17754),
            .I(n25));
    Odrv4 I__4279 (
            .O(N__17749),
            .I(n25));
    LocalMux I__4278 (
            .O(N__17746),
            .I(n25));
    SRMux I__4277 (
            .O(N__17737),
            .I(N__17733));
    SRMux I__4276 (
            .O(N__17736),
            .I(N__17730));
    LocalMux I__4275 (
            .O(N__17733),
            .I(N__17726));
    LocalMux I__4274 (
            .O(N__17730),
            .I(N__17723));
    SRMux I__4273 (
            .O(N__17729),
            .I(N__17720));
    Span4Mux_v I__4272 (
            .O(N__17726),
            .I(N__17713));
    Span4Mux_h I__4271 (
            .O(N__17723),
            .I(N__17713));
    LocalMux I__4270 (
            .O(N__17720),
            .I(N__17713));
    Span4Mux_v I__4269 (
            .O(N__17713),
            .I(N__17709));
    SRMux I__4268 (
            .O(N__17712),
            .I(N__17706));
    Span4Mux_h I__4267 (
            .O(N__17709),
            .I(N__17701));
    LocalMux I__4266 (
            .O(N__17706),
            .I(N__17701));
    Span4Mux_h I__4265 (
            .O(N__17701),
            .I(N__17698));
    Odrv4 I__4264 (
            .O(N__17698),
            .I(\line_buffer.n633 ));
    CascadeMux I__4263 (
            .O(N__17695),
            .I(N__17690));
    InMux I__4262 (
            .O(N__17694),
            .I(N__17687));
    InMux I__4261 (
            .O(N__17693),
            .I(N__17679));
    InMux I__4260 (
            .O(N__17690),
            .I(N__17679));
    LocalMux I__4259 (
            .O(N__17687),
            .I(N__17676));
    InMux I__4258 (
            .O(N__17686),
            .I(N__17673));
    CascadeMux I__4257 (
            .O(N__17685),
            .I(N__17669));
    InMux I__4256 (
            .O(N__17684),
            .I(N__17665));
    LocalMux I__4255 (
            .O(N__17679),
            .I(N__17662));
    Span4Mux_v I__4254 (
            .O(N__17676),
            .I(N__17657));
    LocalMux I__4253 (
            .O(N__17673),
            .I(N__17657));
    InMux I__4252 (
            .O(N__17672),
            .I(N__17652));
    InMux I__4251 (
            .O(N__17669),
            .I(N__17652));
    InMux I__4250 (
            .O(N__17668),
            .I(N__17646));
    LocalMux I__4249 (
            .O(N__17665),
            .I(N__17641));
    Span4Mux_v I__4248 (
            .O(N__17662),
            .I(N__17641));
    Span4Mux_v I__4247 (
            .O(N__17657),
            .I(N__17636));
    LocalMux I__4246 (
            .O(N__17652),
            .I(N__17636));
    InMux I__4245 (
            .O(N__17651),
            .I(N__17632));
    InMux I__4244 (
            .O(N__17650),
            .I(N__17629));
    InMux I__4243 (
            .O(N__17649),
            .I(N__17626));
    LocalMux I__4242 (
            .O(N__17646),
            .I(N__17621));
    Span4Mux_h I__4241 (
            .O(N__17641),
            .I(N__17621));
    Span4Mux_h I__4240 (
            .O(N__17636),
            .I(N__17618));
    InMux I__4239 (
            .O(N__17635),
            .I(N__17615));
    LocalMux I__4238 (
            .O(N__17632),
            .I(TX_ADDR_13));
    LocalMux I__4237 (
            .O(N__17629),
            .I(TX_ADDR_13));
    LocalMux I__4236 (
            .O(N__17626),
            .I(TX_ADDR_13));
    Odrv4 I__4235 (
            .O(N__17621),
            .I(TX_ADDR_13));
    Odrv4 I__4234 (
            .O(N__17618),
            .I(TX_ADDR_13));
    LocalMux I__4233 (
            .O(N__17615),
            .I(TX_ADDR_13));
    InMux I__4232 (
            .O(N__17602),
            .I(N__17599));
    LocalMux I__4231 (
            .O(N__17599),
            .I(N__17596));
    Span4Mux_v I__4230 (
            .O(N__17596),
            .I(N__17593));
    Odrv4 I__4229 (
            .O(N__17593),
            .I(TX_DATA_4));
    ClkMux I__4228 (
            .O(N__17590),
            .I(N__17584));
    ClkMux I__4227 (
            .O(N__17589),
            .I(N__17581));
    ClkMux I__4226 (
            .O(N__17588),
            .I(N__17576));
    ClkMux I__4225 (
            .O(N__17587),
            .I(N__17573));
    LocalMux I__4224 (
            .O(N__17584),
            .I(N__17569));
    LocalMux I__4223 (
            .O(N__17581),
            .I(N__17566));
    ClkMux I__4222 (
            .O(N__17580),
            .I(N__17563));
    ClkMux I__4221 (
            .O(N__17579),
            .I(N__17560));
    LocalMux I__4220 (
            .O(N__17576),
            .I(N__17555));
    LocalMux I__4219 (
            .O(N__17573),
            .I(N__17552));
    ClkMux I__4218 (
            .O(N__17572),
            .I(N__17549));
    Span4Mux_s2_v I__4217 (
            .O(N__17569),
            .I(N__17541));
    Span4Mux_h I__4216 (
            .O(N__17566),
            .I(N__17541));
    LocalMux I__4215 (
            .O(N__17563),
            .I(N__17541));
    LocalMux I__4214 (
            .O(N__17560),
            .I(N__17538));
    ClkMux I__4213 (
            .O(N__17559),
            .I(N__17535));
    ClkMux I__4212 (
            .O(N__17558),
            .I(N__17532));
    Span4Mux_s2_v I__4211 (
            .O(N__17555),
            .I(N__17522));
    Span4Mux_h I__4210 (
            .O(N__17552),
            .I(N__17522));
    LocalMux I__4209 (
            .O(N__17549),
            .I(N__17522));
    ClkMux I__4208 (
            .O(N__17548),
            .I(N__17519));
    Span4Mux_v I__4207 (
            .O(N__17541),
            .I(N__17509));
    Span4Mux_h I__4206 (
            .O(N__17538),
            .I(N__17509));
    LocalMux I__4205 (
            .O(N__17535),
            .I(N__17509));
    LocalMux I__4204 (
            .O(N__17532),
            .I(N__17506));
    ClkMux I__4203 (
            .O(N__17531),
            .I(N__17503));
    ClkMux I__4202 (
            .O(N__17530),
            .I(N__17500));
    ClkMux I__4201 (
            .O(N__17529),
            .I(N__17492));
    Span4Mux_v I__4200 (
            .O(N__17522),
            .I(N__17485));
    LocalMux I__4199 (
            .O(N__17519),
            .I(N__17485));
    ClkMux I__4198 (
            .O(N__17518),
            .I(N__17482));
    ClkMux I__4197 (
            .O(N__17517),
            .I(N__17478));
    ClkMux I__4196 (
            .O(N__17516),
            .I(N__17475));
    Span4Mux_v I__4195 (
            .O(N__17509),
            .I(N__17467));
    Span4Mux_h I__4194 (
            .O(N__17506),
            .I(N__17467));
    LocalMux I__4193 (
            .O(N__17503),
            .I(N__17467));
    LocalMux I__4192 (
            .O(N__17500),
            .I(N__17464));
    ClkMux I__4191 (
            .O(N__17499),
            .I(N__17461));
    ClkMux I__4190 (
            .O(N__17498),
            .I(N__17458));
    ClkMux I__4189 (
            .O(N__17497),
            .I(N__17454));
    ClkMux I__4188 (
            .O(N__17496),
            .I(N__17450));
    ClkMux I__4187 (
            .O(N__17495),
            .I(N__17447));
    LocalMux I__4186 (
            .O(N__17492),
            .I(N__17443));
    ClkMux I__4185 (
            .O(N__17491),
            .I(N__17440));
    ClkMux I__4184 (
            .O(N__17490),
            .I(N__17437));
    Span4Mux_v I__4183 (
            .O(N__17485),
            .I(N__17429));
    LocalMux I__4182 (
            .O(N__17482),
            .I(N__17429));
    ClkMux I__4181 (
            .O(N__17481),
            .I(N__17426));
    LocalMux I__4180 (
            .O(N__17478),
            .I(N__17420));
    LocalMux I__4179 (
            .O(N__17475),
            .I(N__17416));
    ClkMux I__4178 (
            .O(N__17474),
            .I(N__17413));
    Span4Mux_v I__4177 (
            .O(N__17467),
            .I(N__17404));
    Span4Mux_h I__4176 (
            .O(N__17464),
            .I(N__17404));
    LocalMux I__4175 (
            .O(N__17461),
            .I(N__17404));
    LocalMux I__4174 (
            .O(N__17458),
            .I(N__17401));
    ClkMux I__4173 (
            .O(N__17457),
            .I(N__17398));
    LocalMux I__4172 (
            .O(N__17454),
            .I(N__17393));
    ClkMux I__4171 (
            .O(N__17453),
            .I(N__17390));
    LocalMux I__4170 (
            .O(N__17450),
            .I(N__17385));
    LocalMux I__4169 (
            .O(N__17447),
            .I(N__17385));
    ClkMux I__4168 (
            .O(N__17446),
            .I(N__17382));
    Span4Mux_h I__4167 (
            .O(N__17443),
            .I(N__17375));
    LocalMux I__4166 (
            .O(N__17440),
            .I(N__17375));
    LocalMux I__4165 (
            .O(N__17437),
            .I(N__17375));
    ClkMux I__4164 (
            .O(N__17436),
            .I(N__17372));
    ClkMux I__4163 (
            .O(N__17435),
            .I(N__17369));
    ClkMux I__4162 (
            .O(N__17434),
            .I(N__17366));
    Span4Mux_v I__4161 (
            .O(N__17429),
            .I(N__17361));
    LocalMux I__4160 (
            .O(N__17426),
            .I(N__17361));
    ClkMux I__4159 (
            .O(N__17425),
            .I(N__17358));
    ClkMux I__4158 (
            .O(N__17424),
            .I(N__17355));
    ClkMux I__4157 (
            .O(N__17423),
            .I(N__17352));
    Span4Mux_v I__4156 (
            .O(N__17420),
            .I(N__17349));
    ClkMux I__4155 (
            .O(N__17419),
            .I(N__17346));
    Span4Mux_v I__4154 (
            .O(N__17416),
            .I(N__17341));
    LocalMux I__4153 (
            .O(N__17413),
            .I(N__17341));
    ClkMux I__4152 (
            .O(N__17412),
            .I(N__17338));
    ClkMux I__4151 (
            .O(N__17411),
            .I(N__17334));
    Span4Mux_v I__4150 (
            .O(N__17404),
            .I(N__17320));
    Span4Mux_h I__4149 (
            .O(N__17401),
            .I(N__17320));
    LocalMux I__4148 (
            .O(N__17398),
            .I(N__17320));
    ClkMux I__4147 (
            .O(N__17397),
            .I(N__17317));
    ClkMux I__4146 (
            .O(N__17396),
            .I(N__17314));
    Span4Mux_v I__4145 (
            .O(N__17393),
            .I(N__17306));
    LocalMux I__4144 (
            .O(N__17390),
            .I(N__17306));
    Span4Mux_v I__4143 (
            .O(N__17385),
            .I(N__17301));
    LocalMux I__4142 (
            .O(N__17382),
            .I(N__17301));
    Span4Mux_h I__4141 (
            .O(N__17375),
            .I(N__17292));
    LocalMux I__4140 (
            .O(N__17372),
            .I(N__17292));
    LocalMux I__4139 (
            .O(N__17369),
            .I(N__17292));
    LocalMux I__4138 (
            .O(N__17366),
            .I(N__17292));
    Span4Mux_v I__4137 (
            .O(N__17361),
            .I(N__17287));
    LocalMux I__4136 (
            .O(N__17358),
            .I(N__17287));
    LocalMux I__4135 (
            .O(N__17355),
            .I(N__17282));
    LocalMux I__4134 (
            .O(N__17352),
            .I(N__17282));
    Span4Mux_h I__4133 (
            .O(N__17349),
            .I(N__17277));
    LocalMux I__4132 (
            .O(N__17346),
            .I(N__17277));
    Span4Mux_v I__4131 (
            .O(N__17341),
            .I(N__17272));
    LocalMux I__4130 (
            .O(N__17338),
            .I(N__17272));
    ClkMux I__4129 (
            .O(N__17337),
            .I(N__17269));
    LocalMux I__4128 (
            .O(N__17334),
            .I(N__17265));
    ClkMux I__4127 (
            .O(N__17333),
            .I(N__17262));
    ClkMux I__4126 (
            .O(N__17332),
            .I(N__17259));
    ClkMux I__4125 (
            .O(N__17331),
            .I(N__17256));
    ClkMux I__4124 (
            .O(N__17330),
            .I(N__17253));
    ClkMux I__4123 (
            .O(N__17329),
            .I(N__17250));
    ClkMux I__4122 (
            .O(N__17328),
            .I(N__17246));
    ClkMux I__4121 (
            .O(N__17327),
            .I(N__17242));
    Span4Mux_v I__4120 (
            .O(N__17320),
            .I(N__17236));
    LocalMux I__4119 (
            .O(N__17317),
            .I(N__17236));
    LocalMux I__4118 (
            .O(N__17314),
            .I(N__17233));
    ClkMux I__4117 (
            .O(N__17313),
            .I(N__17230));
    IoInMux I__4116 (
            .O(N__17312),
            .I(N__17227));
    ClkMux I__4115 (
            .O(N__17311),
            .I(N__17222));
    Span4Mux_v I__4114 (
            .O(N__17306),
            .I(N__17219));
    Span4Mux_v I__4113 (
            .O(N__17301),
            .I(N__17214));
    Span4Mux_v I__4112 (
            .O(N__17292),
            .I(N__17214));
    Span4Mux_v I__4111 (
            .O(N__17287),
            .I(N__17210));
    Span4Mux_v I__4110 (
            .O(N__17282),
            .I(N__17207));
    Span4Mux_v I__4109 (
            .O(N__17277),
            .I(N__17200));
    Span4Mux_h I__4108 (
            .O(N__17272),
            .I(N__17200));
    LocalMux I__4107 (
            .O(N__17269),
            .I(N__17200));
    ClkMux I__4106 (
            .O(N__17268),
            .I(N__17197));
    Span4Mux_v I__4105 (
            .O(N__17265),
            .I(N__17190));
    LocalMux I__4104 (
            .O(N__17262),
            .I(N__17190));
    LocalMux I__4103 (
            .O(N__17259),
            .I(N__17187));
    LocalMux I__4102 (
            .O(N__17256),
            .I(N__17180));
    LocalMux I__4101 (
            .O(N__17253),
            .I(N__17180));
    LocalMux I__4100 (
            .O(N__17250),
            .I(N__17180));
    ClkMux I__4099 (
            .O(N__17249),
            .I(N__17177));
    LocalMux I__4098 (
            .O(N__17246),
            .I(N__17174));
    ClkMux I__4097 (
            .O(N__17245),
            .I(N__17171));
    LocalMux I__4096 (
            .O(N__17242),
            .I(N__17168));
    ClkMux I__4095 (
            .O(N__17241),
            .I(N__17165));
    Span4Mux_v I__4094 (
            .O(N__17236),
            .I(N__17158));
    Span4Mux_h I__4093 (
            .O(N__17233),
            .I(N__17158));
    LocalMux I__4092 (
            .O(N__17230),
            .I(N__17158));
    LocalMux I__4091 (
            .O(N__17227),
            .I(N__17155));
    ClkMux I__4090 (
            .O(N__17226),
            .I(N__17152));
    ClkMux I__4089 (
            .O(N__17225),
            .I(N__17148));
    LocalMux I__4088 (
            .O(N__17222),
            .I(N__17145));
    Span4Mux_v I__4087 (
            .O(N__17219),
            .I(N__17140));
    Span4Mux_v I__4086 (
            .O(N__17214),
            .I(N__17140));
    ClkMux I__4085 (
            .O(N__17213),
            .I(N__17137));
    Span4Mux_h I__4084 (
            .O(N__17210),
            .I(N__17130));
    Span4Mux_v I__4083 (
            .O(N__17207),
            .I(N__17130));
    Span4Mux_v I__4082 (
            .O(N__17200),
            .I(N__17130));
    LocalMux I__4081 (
            .O(N__17197),
            .I(N__17127));
    ClkMux I__4080 (
            .O(N__17196),
            .I(N__17124));
    ClkMux I__4079 (
            .O(N__17195),
            .I(N__17121));
    Span4Mux_v I__4078 (
            .O(N__17190),
            .I(N__17112));
    Span4Mux_h I__4077 (
            .O(N__17187),
            .I(N__17112));
    Span4Mux_v I__4076 (
            .O(N__17180),
            .I(N__17112));
    LocalMux I__4075 (
            .O(N__17177),
            .I(N__17112));
    Span4Mux_h I__4074 (
            .O(N__17174),
            .I(N__17109));
    LocalMux I__4073 (
            .O(N__17171),
            .I(N__17106));
    Span12Mux_h I__4072 (
            .O(N__17168),
            .I(N__17103));
    LocalMux I__4071 (
            .O(N__17165),
            .I(N__17100));
    Span4Mux_v I__4070 (
            .O(N__17158),
            .I(N__17097));
    Span4Mux_s1_v I__4069 (
            .O(N__17155),
            .I(N__17094));
    LocalMux I__4068 (
            .O(N__17152),
            .I(N__17091));
    ClkMux I__4067 (
            .O(N__17151),
            .I(N__17088));
    LocalMux I__4066 (
            .O(N__17148),
            .I(N__17085));
    Sp12to4 I__4065 (
            .O(N__17145),
            .I(N__17080));
    Sp12to4 I__4064 (
            .O(N__17140),
            .I(N__17080));
    LocalMux I__4063 (
            .O(N__17137),
            .I(N__17075));
    Sp12to4 I__4062 (
            .O(N__17130),
            .I(N__17075));
    Span12Mux_h I__4061 (
            .O(N__17127),
            .I(N__17068));
    LocalMux I__4060 (
            .O(N__17124),
            .I(N__17068));
    LocalMux I__4059 (
            .O(N__17121),
            .I(N__17068));
    Span4Mux_v I__4058 (
            .O(N__17112),
            .I(N__17065));
    Span4Mux_v I__4057 (
            .O(N__17109),
            .I(N__17060));
    Span4Mux_h I__4056 (
            .O(N__17106),
            .I(N__17060));
    Span12Mux_v I__4055 (
            .O(N__17103),
            .I(N__17055));
    Span12Mux_h I__4054 (
            .O(N__17100),
            .I(N__17055));
    Sp12to4 I__4053 (
            .O(N__17097),
            .I(N__17048));
    Sp12to4 I__4052 (
            .O(N__17094),
            .I(N__17048));
    Sp12to4 I__4051 (
            .O(N__17091),
            .I(N__17048));
    LocalMux I__4050 (
            .O(N__17088),
            .I(N__17045));
    Span12Mux_h I__4049 (
            .O(N__17085),
            .I(N__17042));
    Span12Mux_h I__4048 (
            .O(N__17080),
            .I(N__17033));
    Span12Mux_h I__4047 (
            .O(N__17075),
            .I(N__17033));
    Span12Mux_v I__4046 (
            .O(N__17068),
            .I(N__17033));
    Sp12to4 I__4045 (
            .O(N__17065),
            .I(N__17033));
    Span4Mux_h I__4044 (
            .O(N__17060),
            .I(N__17030));
    Span12Mux_v I__4043 (
            .O(N__17055),
            .I(N__17023));
    Span12Mux_h I__4042 (
            .O(N__17048),
            .I(N__17023));
    Span12Mux_h I__4041 (
            .O(N__17045),
            .I(N__17023));
    Odrv12 I__4040 (
            .O(N__17042),
            .I(ADV_CLK_c));
    Odrv12 I__4039 (
            .O(N__17033),
            .I(ADV_CLK_c));
    Odrv4 I__4038 (
            .O(N__17030),
            .I(ADV_CLK_c));
    Odrv12 I__4037 (
            .O(N__17023),
            .I(ADV_CLK_c));
    InMux I__4036 (
            .O(N__17014),
            .I(N__17011));
    LocalMux I__4035 (
            .O(N__17011),
            .I(N__17008));
    Span4Mux_h I__4034 (
            .O(N__17008),
            .I(N__17005));
    Span4Mux_h I__4033 (
            .O(N__17005),
            .I(N__17002));
    Odrv4 I__4032 (
            .O(N__17002),
            .I(\line_buffer.n716 ));
    InMux I__4031 (
            .O(N__16999),
            .I(N__16996));
    LocalMux I__4030 (
            .O(N__16996),
            .I(N__16993));
    Span4Mux_v I__4029 (
            .O(N__16993),
            .I(N__16990));
    Span4Mux_v I__4028 (
            .O(N__16990),
            .I(N__16987));
    Sp12to4 I__4027 (
            .O(N__16987),
            .I(N__16984));
    Odrv12 I__4026 (
            .O(N__16984),
            .I(\line_buffer.n724 ));
    InMux I__4025 (
            .O(N__16981),
            .I(N__16978));
    LocalMux I__4024 (
            .O(N__16978),
            .I(\line_buffer.n3046 ));
    InMux I__4023 (
            .O(N__16975),
            .I(N__16972));
    LocalMux I__4022 (
            .O(N__16972),
            .I(N__16969));
    Odrv4 I__4021 (
            .O(N__16969),
            .I(\receive_module.n132 ));
    CascadeMux I__4020 (
            .O(N__16966),
            .I(N__16963));
    CascadeBuf I__4019 (
            .O(N__16963),
            .I(N__16959));
    CascadeMux I__4018 (
            .O(N__16962),
            .I(N__16956));
    CascadeMux I__4017 (
            .O(N__16959),
            .I(N__16953));
    CascadeBuf I__4016 (
            .O(N__16956),
            .I(N__16950));
    CascadeBuf I__4015 (
            .O(N__16953),
            .I(N__16947));
    CascadeMux I__4014 (
            .O(N__16950),
            .I(N__16944));
    CascadeMux I__4013 (
            .O(N__16947),
            .I(N__16941));
    CascadeBuf I__4012 (
            .O(N__16944),
            .I(N__16938));
    CascadeBuf I__4011 (
            .O(N__16941),
            .I(N__16935));
    CascadeMux I__4010 (
            .O(N__16938),
            .I(N__16932));
    CascadeMux I__4009 (
            .O(N__16935),
            .I(N__16929));
    CascadeBuf I__4008 (
            .O(N__16932),
            .I(N__16926));
    CascadeBuf I__4007 (
            .O(N__16929),
            .I(N__16923));
    CascadeMux I__4006 (
            .O(N__16926),
            .I(N__16920));
    CascadeMux I__4005 (
            .O(N__16923),
            .I(N__16917));
    CascadeBuf I__4004 (
            .O(N__16920),
            .I(N__16914));
    CascadeBuf I__4003 (
            .O(N__16917),
            .I(N__16911));
    CascadeMux I__4002 (
            .O(N__16914),
            .I(N__16908));
    CascadeMux I__4001 (
            .O(N__16911),
            .I(N__16905));
    CascadeBuf I__4000 (
            .O(N__16908),
            .I(N__16902));
    CascadeBuf I__3999 (
            .O(N__16905),
            .I(N__16899));
    CascadeMux I__3998 (
            .O(N__16902),
            .I(N__16896));
    CascadeMux I__3997 (
            .O(N__16899),
            .I(N__16893));
    CascadeBuf I__3996 (
            .O(N__16896),
            .I(N__16890));
    CascadeBuf I__3995 (
            .O(N__16893),
            .I(N__16887));
    CascadeMux I__3994 (
            .O(N__16890),
            .I(N__16884));
    CascadeMux I__3993 (
            .O(N__16887),
            .I(N__16881));
    CascadeBuf I__3992 (
            .O(N__16884),
            .I(N__16878));
    CascadeBuf I__3991 (
            .O(N__16881),
            .I(N__16875));
    CascadeMux I__3990 (
            .O(N__16878),
            .I(N__16872));
    CascadeMux I__3989 (
            .O(N__16875),
            .I(N__16869));
    CascadeBuf I__3988 (
            .O(N__16872),
            .I(N__16866));
    CascadeBuf I__3987 (
            .O(N__16869),
            .I(N__16863));
    CascadeMux I__3986 (
            .O(N__16866),
            .I(N__16860));
    CascadeMux I__3985 (
            .O(N__16863),
            .I(N__16857));
    CascadeBuf I__3984 (
            .O(N__16860),
            .I(N__16854));
    CascadeBuf I__3983 (
            .O(N__16857),
            .I(N__16851));
    CascadeMux I__3982 (
            .O(N__16854),
            .I(N__16848));
    CascadeMux I__3981 (
            .O(N__16851),
            .I(N__16845));
    CascadeBuf I__3980 (
            .O(N__16848),
            .I(N__16842));
    CascadeBuf I__3979 (
            .O(N__16845),
            .I(N__16839));
    CascadeMux I__3978 (
            .O(N__16842),
            .I(N__16836));
    CascadeMux I__3977 (
            .O(N__16839),
            .I(N__16833));
    CascadeBuf I__3976 (
            .O(N__16836),
            .I(N__16830));
    CascadeBuf I__3975 (
            .O(N__16833),
            .I(N__16827));
    CascadeMux I__3974 (
            .O(N__16830),
            .I(N__16824));
    CascadeMux I__3973 (
            .O(N__16827),
            .I(N__16821));
    CascadeBuf I__3972 (
            .O(N__16824),
            .I(N__16818));
    CascadeBuf I__3971 (
            .O(N__16821),
            .I(N__16815));
    CascadeMux I__3970 (
            .O(N__16818),
            .I(N__16812));
    CascadeMux I__3969 (
            .O(N__16815),
            .I(N__16809));
    CascadeBuf I__3968 (
            .O(N__16812),
            .I(N__16806));
    CascadeBuf I__3967 (
            .O(N__16809),
            .I(N__16803));
    CascadeMux I__3966 (
            .O(N__16806),
            .I(N__16800));
    CascadeMux I__3965 (
            .O(N__16803),
            .I(N__16797));
    CascadeBuf I__3964 (
            .O(N__16800),
            .I(N__16794));
    CascadeBuf I__3963 (
            .O(N__16797),
            .I(N__16791));
    CascadeMux I__3962 (
            .O(N__16794),
            .I(N__16788));
    CascadeMux I__3961 (
            .O(N__16791),
            .I(N__16785));
    CascadeBuf I__3960 (
            .O(N__16788),
            .I(N__16782));
    InMux I__3959 (
            .O(N__16785),
            .I(N__16779));
    CascadeMux I__3958 (
            .O(N__16782),
            .I(N__16776));
    LocalMux I__3957 (
            .O(N__16779),
            .I(N__16773));
    InMux I__3956 (
            .O(N__16776),
            .I(N__16770));
    Span4Mux_h I__3955 (
            .O(N__16773),
            .I(N__16767));
    LocalMux I__3954 (
            .O(N__16770),
            .I(N__16764));
    Span4Mux_h I__3953 (
            .O(N__16767),
            .I(N__16760));
    Span12Mux_s1_v I__3952 (
            .O(N__16764),
            .I(N__16757));
    InMux I__3951 (
            .O(N__16763),
            .I(N__16754));
    Sp12to4 I__3950 (
            .O(N__16760),
            .I(N__16750));
    Span12Mux_v I__3949 (
            .O(N__16757),
            .I(N__16747));
    LocalMux I__3948 (
            .O(N__16754),
            .I(N__16744));
    InMux I__3947 (
            .O(N__16753),
            .I(N__16741));
    Span12Mux_v I__3946 (
            .O(N__16750),
            .I(N__16736));
    Span12Mux_h I__3945 (
            .O(N__16747),
            .I(N__16736));
    Odrv4 I__3944 (
            .O(N__16744),
            .I(RX_ADDR_4));
    LocalMux I__3943 (
            .O(N__16741),
            .I(RX_ADDR_4));
    Odrv12 I__3942 (
            .O(N__16736),
            .I(RX_ADDR_4));
    CascadeMux I__3941 (
            .O(N__16729),
            .I(N__16726));
    InMux I__3940 (
            .O(N__16726),
            .I(N__16723));
    LocalMux I__3939 (
            .O(N__16723),
            .I(N__16720));
    Odrv4 I__3938 (
            .O(N__16720),
            .I(\receive_module.n130 ));
    CascadeMux I__3937 (
            .O(N__16717),
            .I(N__16713));
    CascadeMux I__3936 (
            .O(N__16716),
            .I(N__16710));
    CascadeBuf I__3935 (
            .O(N__16713),
            .I(N__16707));
    CascadeBuf I__3934 (
            .O(N__16710),
            .I(N__16704));
    CascadeMux I__3933 (
            .O(N__16707),
            .I(N__16701));
    CascadeMux I__3932 (
            .O(N__16704),
            .I(N__16698));
    CascadeBuf I__3931 (
            .O(N__16701),
            .I(N__16695));
    CascadeBuf I__3930 (
            .O(N__16698),
            .I(N__16692));
    CascadeMux I__3929 (
            .O(N__16695),
            .I(N__16689));
    CascadeMux I__3928 (
            .O(N__16692),
            .I(N__16686));
    CascadeBuf I__3927 (
            .O(N__16689),
            .I(N__16683));
    CascadeBuf I__3926 (
            .O(N__16686),
            .I(N__16680));
    CascadeMux I__3925 (
            .O(N__16683),
            .I(N__16677));
    CascadeMux I__3924 (
            .O(N__16680),
            .I(N__16674));
    CascadeBuf I__3923 (
            .O(N__16677),
            .I(N__16671));
    CascadeBuf I__3922 (
            .O(N__16674),
            .I(N__16668));
    CascadeMux I__3921 (
            .O(N__16671),
            .I(N__16665));
    CascadeMux I__3920 (
            .O(N__16668),
            .I(N__16662));
    CascadeBuf I__3919 (
            .O(N__16665),
            .I(N__16659));
    CascadeBuf I__3918 (
            .O(N__16662),
            .I(N__16656));
    CascadeMux I__3917 (
            .O(N__16659),
            .I(N__16653));
    CascadeMux I__3916 (
            .O(N__16656),
            .I(N__16650));
    CascadeBuf I__3915 (
            .O(N__16653),
            .I(N__16647));
    CascadeBuf I__3914 (
            .O(N__16650),
            .I(N__16644));
    CascadeMux I__3913 (
            .O(N__16647),
            .I(N__16641));
    CascadeMux I__3912 (
            .O(N__16644),
            .I(N__16638));
    CascadeBuf I__3911 (
            .O(N__16641),
            .I(N__16635));
    CascadeBuf I__3910 (
            .O(N__16638),
            .I(N__16632));
    CascadeMux I__3909 (
            .O(N__16635),
            .I(N__16629));
    CascadeMux I__3908 (
            .O(N__16632),
            .I(N__16626));
    CascadeBuf I__3907 (
            .O(N__16629),
            .I(N__16623));
    CascadeBuf I__3906 (
            .O(N__16626),
            .I(N__16620));
    CascadeMux I__3905 (
            .O(N__16623),
            .I(N__16617));
    CascadeMux I__3904 (
            .O(N__16620),
            .I(N__16614));
    CascadeBuf I__3903 (
            .O(N__16617),
            .I(N__16611));
    CascadeBuf I__3902 (
            .O(N__16614),
            .I(N__16608));
    CascadeMux I__3901 (
            .O(N__16611),
            .I(N__16605));
    CascadeMux I__3900 (
            .O(N__16608),
            .I(N__16602));
    CascadeBuf I__3899 (
            .O(N__16605),
            .I(N__16599));
    CascadeBuf I__3898 (
            .O(N__16602),
            .I(N__16596));
    CascadeMux I__3897 (
            .O(N__16599),
            .I(N__16593));
    CascadeMux I__3896 (
            .O(N__16596),
            .I(N__16590));
    CascadeBuf I__3895 (
            .O(N__16593),
            .I(N__16587));
    CascadeBuf I__3894 (
            .O(N__16590),
            .I(N__16584));
    CascadeMux I__3893 (
            .O(N__16587),
            .I(N__16581));
    CascadeMux I__3892 (
            .O(N__16584),
            .I(N__16578));
    CascadeBuf I__3891 (
            .O(N__16581),
            .I(N__16575));
    CascadeBuf I__3890 (
            .O(N__16578),
            .I(N__16572));
    CascadeMux I__3889 (
            .O(N__16575),
            .I(N__16569));
    CascadeMux I__3888 (
            .O(N__16572),
            .I(N__16566));
    CascadeBuf I__3887 (
            .O(N__16569),
            .I(N__16563));
    CascadeBuf I__3886 (
            .O(N__16566),
            .I(N__16560));
    CascadeMux I__3885 (
            .O(N__16563),
            .I(N__16557));
    CascadeMux I__3884 (
            .O(N__16560),
            .I(N__16554));
    CascadeBuf I__3883 (
            .O(N__16557),
            .I(N__16551));
    CascadeBuf I__3882 (
            .O(N__16554),
            .I(N__16548));
    CascadeMux I__3881 (
            .O(N__16551),
            .I(N__16545));
    CascadeMux I__3880 (
            .O(N__16548),
            .I(N__16542));
    CascadeBuf I__3879 (
            .O(N__16545),
            .I(N__16539));
    CascadeBuf I__3878 (
            .O(N__16542),
            .I(N__16536));
    CascadeMux I__3877 (
            .O(N__16539),
            .I(N__16533));
    CascadeMux I__3876 (
            .O(N__16536),
            .I(N__16530));
    InMux I__3875 (
            .O(N__16533),
            .I(N__16527));
    InMux I__3874 (
            .O(N__16530),
            .I(N__16524));
    LocalMux I__3873 (
            .O(N__16527),
            .I(N__16520));
    LocalMux I__3872 (
            .O(N__16524),
            .I(N__16517));
    InMux I__3871 (
            .O(N__16523),
            .I(N__16514));
    Span12Mux_h I__3870 (
            .O(N__16520),
            .I(N__16508));
    Span12Mux_h I__3869 (
            .O(N__16517),
            .I(N__16508));
    LocalMux I__3868 (
            .O(N__16514),
            .I(N__16505));
    InMux I__3867 (
            .O(N__16513),
            .I(N__16502));
    Span12Mux_v I__3866 (
            .O(N__16508),
            .I(N__16499));
    Odrv4 I__3865 (
            .O(N__16505),
            .I(RX_ADDR_6));
    LocalMux I__3864 (
            .O(N__16502),
            .I(RX_ADDR_6));
    Odrv12 I__3863 (
            .O(N__16499),
            .I(RX_ADDR_6));
    InMux I__3862 (
            .O(N__16492),
            .I(N__16489));
    LocalMux I__3861 (
            .O(N__16489),
            .I(N__16486));
    Odrv4 I__3860 (
            .O(N__16486),
            .I(\receive_module.n126 ));
    CascadeMux I__3859 (
            .O(N__16483),
            .I(N__16476));
    CascadeMux I__3858 (
            .O(N__16482),
            .I(N__16472));
    CascadeMux I__3857 (
            .O(N__16481),
            .I(N__16467));
    CascadeMux I__3856 (
            .O(N__16480),
            .I(N__16463));
    CascadeMux I__3855 (
            .O(N__16479),
            .I(N__16460));
    InMux I__3854 (
            .O(N__16476),
            .I(N__16457));
    InMux I__3853 (
            .O(N__16475),
            .I(N__16452));
    InMux I__3852 (
            .O(N__16472),
            .I(N__16452));
    InMux I__3851 (
            .O(N__16471),
            .I(N__16449));
    CascadeMux I__3850 (
            .O(N__16470),
            .I(N__16446));
    InMux I__3849 (
            .O(N__16467),
            .I(N__16440));
    InMux I__3848 (
            .O(N__16466),
            .I(N__16433));
    InMux I__3847 (
            .O(N__16463),
            .I(N__16433));
    InMux I__3846 (
            .O(N__16460),
            .I(N__16433));
    LocalMux I__3845 (
            .O(N__16457),
            .I(N__16427));
    LocalMux I__3844 (
            .O(N__16452),
            .I(N__16427));
    LocalMux I__3843 (
            .O(N__16449),
            .I(N__16424));
    InMux I__3842 (
            .O(N__16446),
            .I(N__16415));
    InMux I__3841 (
            .O(N__16445),
            .I(N__16415));
    InMux I__3840 (
            .O(N__16444),
            .I(N__16415));
    InMux I__3839 (
            .O(N__16443),
            .I(N__16415));
    LocalMux I__3838 (
            .O(N__16440),
            .I(N__16410));
    LocalMux I__3837 (
            .O(N__16433),
            .I(N__16410));
    InMux I__3836 (
            .O(N__16432),
            .I(N__16407));
    Span4Mux_v I__3835 (
            .O(N__16427),
            .I(N__16402));
    Span4Mux_v I__3834 (
            .O(N__16424),
            .I(N__16399));
    LocalMux I__3833 (
            .O(N__16415),
            .I(N__16392));
    Span4Mux_h I__3832 (
            .O(N__16410),
            .I(N__16392));
    LocalMux I__3831 (
            .O(N__16407),
            .I(N__16392));
    InMux I__3830 (
            .O(N__16406),
            .I(N__16387));
    InMux I__3829 (
            .O(N__16405),
            .I(N__16387));
    Span4Mux_h I__3828 (
            .O(N__16402),
            .I(N__16377));
    Span4Mux_h I__3827 (
            .O(N__16399),
            .I(N__16377));
    Span4Mux_v I__3826 (
            .O(N__16392),
            .I(N__16377));
    LocalMux I__3825 (
            .O(N__16387),
            .I(N__16377));
    InMux I__3824 (
            .O(N__16386),
            .I(N__16374));
    Span4Mux_v I__3823 (
            .O(N__16377),
            .I(N__16371));
    LocalMux I__3822 (
            .O(N__16374),
            .I(N__16368));
    Span4Mux_v I__3821 (
            .O(N__16371),
            .I(N__16365));
    Span12Mux_v I__3820 (
            .O(N__16368),
            .I(N__16362));
    IoSpan4Mux I__3819 (
            .O(N__16365),
            .I(N__16359));
    Odrv12 I__3818 (
            .O(N__16362),
            .I(TVP_VSYNC_c));
    Odrv4 I__3817 (
            .O(N__16359),
            .I(TVP_VSYNC_c));
    CascadeMux I__3816 (
            .O(N__16354),
            .I(N__16350));
    CascadeMux I__3815 (
            .O(N__16353),
            .I(N__16347));
    CascadeBuf I__3814 (
            .O(N__16350),
            .I(N__16344));
    CascadeBuf I__3813 (
            .O(N__16347),
            .I(N__16341));
    CascadeMux I__3812 (
            .O(N__16344),
            .I(N__16338));
    CascadeMux I__3811 (
            .O(N__16341),
            .I(N__16335));
    CascadeBuf I__3810 (
            .O(N__16338),
            .I(N__16332));
    CascadeBuf I__3809 (
            .O(N__16335),
            .I(N__16329));
    CascadeMux I__3808 (
            .O(N__16332),
            .I(N__16326));
    CascadeMux I__3807 (
            .O(N__16329),
            .I(N__16323));
    CascadeBuf I__3806 (
            .O(N__16326),
            .I(N__16320));
    CascadeBuf I__3805 (
            .O(N__16323),
            .I(N__16317));
    CascadeMux I__3804 (
            .O(N__16320),
            .I(N__16314));
    CascadeMux I__3803 (
            .O(N__16317),
            .I(N__16311));
    CascadeBuf I__3802 (
            .O(N__16314),
            .I(N__16308));
    CascadeBuf I__3801 (
            .O(N__16311),
            .I(N__16305));
    CascadeMux I__3800 (
            .O(N__16308),
            .I(N__16302));
    CascadeMux I__3799 (
            .O(N__16305),
            .I(N__16299));
    CascadeBuf I__3798 (
            .O(N__16302),
            .I(N__16296));
    CascadeBuf I__3797 (
            .O(N__16299),
            .I(N__16293));
    CascadeMux I__3796 (
            .O(N__16296),
            .I(N__16290));
    CascadeMux I__3795 (
            .O(N__16293),
            .I(N__16287));
    CascadeBuf I__3794 (
            .O(N__16290),
            .I(N__16284));
    CascadeBuf I__3793 (
            .O(N__16287),
            .I(N__16281));
    CascadeMux I__3792 (
            .O(N__16284),
            .I(N__16278));
    CascadeMux I__3791 (
            .O(N__16281),
            .I(N__16275));
    CascadeBuf I__3790 (
            .O(N__16278),
            .I(N__16272));
    CascadeBuf I__3789 (
            .O(N__16275),
            .I(N__16269));
    CascadeMux I__3788 (
            .O(N__16272),
            .I(N__16266));
    CascadeMux I__3787 (
            .O(N__16269),
            .I(N__16263));
    CascadeBuf I__3786 (
            .O(N__16266),
            .I(N__16260));
    CascadeBuf I__3785 (
            .O(N__16263),
            .I(N__16257));
    CascadeMux I__3784 (
            .O(N__16260),
            .I(N__16254));
    CascadeMux I__3783 (
            .O(N__16257),
            .I(N__16251));
    CascadeBuf I__3782 (
            .O(N__16254),
            .I(N__16248));
    CascadeBuf I__3781 (
            .O(N__16251),
            .I(N__16245));
    CascadeMux I__3780 (
            .O(N__16248),
            .I(N__16242));
    CascadeMux I__3779 (
            .O(N__16245),
            .I(N__16239));
    CascadeBuf I__3778 (
            .O(N__16242),
            .I(N__16236));
    CascadeBuf I__3777 (
            .O(N__16239),
            .I(N__16233));
    CascadeMux I__3776 (
            .O(N__16236),
            .I(N__16230));
    CascadeMux I__3775 (
            .O(N__16233),
            .I(N__16227));
    CascadeBuf I__3774 (
            .O(N__16230),
            .I(N__16224));
    CascadeBuf I__3773 (
            .O(N__16227),
            .I(N__16221));
    CascadeMux I__3772 (
            .O(N__16224),
            .I(N__16218));
    CascadeMux I__3771 (
            .O(N__16221),
            .I(N__16215));
    CascadeBuf I__3770 (
            .O(N__16218),
            .I(N__16212));
    CascadeBuf I__3769 (
            .O(N__16215),
            .I(N__16209));
    CascadeMux I__3768 (
            .O(N__16212),
            .I(N__16206));
    CascadeMux I__3767 (
            .O(N__16209),
            .I(N__16203));
    CascadeBuf I__3766 (
            .O(N__16206),
            .I(N__16200));
    CascadeBuf I__3765 (
            .O(N__16203),
            .I(N__16197));
    CascadeMux I__3764 (
            .O(N__16200),
            .I(N__16194));
    CascadeMux I__3763 (
            .O(N__16197),
            .I(N__16191));
    CascadeBuf I__3762 (
            .O(N__16194),
            .I(N__16188));
    CascadeBuf I__3761 (
            .O(N__16191),
            .I(N__16185));
    CascadeMux I__3760 (
            .O(N__16188),
            .I(N__16182));
    CascadeMux I__3759 (
            .O(N__16185),
            .I(N__16179));
    CascadeBuf I__3758 (
            .O(N__16182),
            .I(N__16176));
    CascadeBuf I__3757 (
            .O(N__16179),
            .I(N__16173));
    CascadeMux I__3756 (
            .O(N__16176),
            .I(N__16170));
    CascadeMux I__3755 (
            .O(N__16173),
            .I(N__16167));
    InMux I__3754 (
            .O(N__16170),
            .I(N__16164));
    InMux I__3753 (
            .O(N__16167),
            .I(N__16161));
    LocalMux I__3752 (
            .O(N__16164),
            .I(N__16157));
    LocalMux I__3751 (
            .O(N__16161),
            .I(N__16154));
    InMux I__3750 (
            .O(N__16160),
            .I(N__16151));
    Span12Mux_h I__3749 (
            .O(N__16157),
            .I(N__16145));
    Span12Mux_h I__3748 (
            .O(N__16154),
            .I(N__16145));
    LocalMux I__3747 (
            .O(N__16151),
            .I(N__16142));
    InMux I__3746 (
            .O(N__16150),
            .I(N__16139));
    Span12Mux_v I__3745 (
            .O(N__16145),
            .I(N__16136));
    Odrv4 I__3744 (
            .O(N__16142),
            .I(RX_ADDR_10));
    LocalMux I__3743 (
            .O(N__16139),
            .I(RX_ADDR_10));
    Odrv12 I__3742 (
            .O(N__16136),
            .I(RX_ADDR_10));
    InMux I__3741 (
            .O(N__16129),
            .I(N__16126));
    LocalMux I__3740 (
            .O(N__16126),
            .I(N__16115));
    ClkMux I__3739 (
            .O(N__16125),
            .I(N__15985));
    ClkMux I__3738 (
            .O(N__16124),
            .I(N__15985));
    ClkMux I__3737 (
            .O(N__16123),
            .I(N__15985));
    ClkMux I__3736 (
            .O(N__16122),
            .I(N__15985));
    ClkMux I__3735 (
            .O(N__16121),
            .I(N__15985));
    ClkMux I__3734 (
            .O(N__16120),
            .I(N__15985));
    ClkMux I__3733 (
            .O(N__16119),
            .I(N__15985));
    ClkMux I__3732 (
            .O(N__16118),
            .I(N__15985));
    Glb2LocalMux I__3731 (
            .O(N__16115),
            .I(N__15985));
    ClkMux I__3730 (
            .O(N__16114),
            .I(N__15985));
    ClkMux I__3729 (
            .O(N__16113),
            .I(N__15985));
    ClkMux I__3728 (
            .O(N__16112),
            .I(N__15985));
    ClkMux I__3727 (
            .O(N__16111),
            .I(N__15985));
    ClkMux I__3726 (
            .O(N__16110),
            .I(N__15985));
    ClkMux I__3725 (
            .O(N__16109),
            .I(N__15985));
    ClkMux I__3724 (
            .O(N__16108),
            .I(N__15985));
    ClkMux I__3723 (
            .O(N__16107),
            .I(N__15985));
    ClkMux I__3722 (
            .O(N__16106),
            .I(N__15985));
    ClkMux I__3721 (
            .O(N__16105),
            .I(N__15985));
    ClkMux I__3720 (
            .O(N__16104),
            .I(N__15985));
    ClkMux I__3719 (
            .O(N__16103),
            .I(N__15985));
    ClkMux I__3718 (
            .O(N__16102),
            .I(N__15985));
    ClkMux I__3717 (
            .O(N__16101),
            .I(N__15985));
    ClkMux I__3716 (
            .O(N__16100),
            .I(N__15985));
    ClkMux I__3715 (
            .O(N__16099),
            .I(N__15985));
    ClkMux I__3714 (
            .O(N__16098),
            .I(N__15985));
    ClkMux I__3713 (
            .O(N__16097),
            .I(N__15985));
    ClkMux I__3712 (
            .O(N__16096),
            .I(N__15985));
    ClkMux I__3711 (
            .O(N__16095),
            .I(N__15985));
    ClkMux I__3710 (
            .O(N__16094),
            .I(N__15985));
    ClkMux I__3709 (
            .O(N__16093),
            .I(N__15985));
    ClkMux I__3708 (
            .O(N__16092),
            .I(N__15985));
    ClkMux I__3707 (
            .O(N__16091),
            .I(N__15985));
    ClkMux I__3706 (
            .O(N__16090),
            .I(N__15985));
    ClkMux I__3705 (
            .O(N__16089),
            .I(N__15985));
    ClkMux I__3704 (
            .O(N__16088),
            .I(N__15985));
    ClkMux I__3703 (
            .O(N__16087),
            .I(N__15985));
    ClkMux I__3702 (
            .O(N__16086),
            .I(N__15985));
    ClkMux I__3701 (
            .O(N__16085),
            .I(N__15985));
    ClkMux I__3700 (
            .O(N__16084),
            .I(N__15985));
    ClkMux I__3699 (
            .O(N__16083),
            .I(N__15985));
    ClkMux I__3698 (
            .O(N__16082),
            .I(N__15985));
    ClkMux I__3697 (
            .O(N__16081),
            .I(N__15985));
    ClkMux I__3696 (
            .O(N__16080),
            .I(N__15985));
    ClkMux I__3695 (
            .O(N__16079),
            .I(N__15985));
    ClkMux I__3694 (
            .O(N__16078),
            .I(N__15985));
    GlobalMux I__3693 (
            .O(N__15985),
            .I(N__15982));
    gio2CtrlBuf I__3692 (
            .O(N__15982),
            .I(TVP_CLK_c));
    SRMux I__3691 (
            .O(N__15979),
            .I(N__15975));
    SRMux I__3690 (
            .O(N__15978),
            .I(N__15972));
    LocalMux I__3689 (
            .O(N__15975),
            .I(N__15969));
    LocalMux I__3688 (
            .O(N__15972),
            .I(N__15961));
    Span4Mux_h I__3687 (
            .O(N__15969),
            .I(N__15958));
    SRMux I__3686 (
            .O(N__15968),
            .I(N__15955));
    SRMux I__3685 (
            .O(N__15967),
            .I(N__15952));
    SRMux I__3684 (
            .O(N__15966),
            .I(N__15949));
    SRMux I__3683 (
            .O(N__15965),
            .I(N__15946));
    SRMux I__3682 (
            .O(N__15964),
            .I(N__15943));
    Span4Mux_v I__3681 (
            .O(N__15961),
            .I(N__15940));
    Span4Mux_h I__3680 (
            .O(N__15958),
            .I(N__15933));
    LocalMux I__3679 (
            .O(N__15955),
            .I(N__15933));
    LocalMux I__3678 (
            .O(N__15952),
            .I(N__15933));
    LocalMux I__3677 (
            .O(N__15949),
            .I(N__15928));
    LocalMux I__3676 (
            .O(N__15946),
            .I(N__15928));
    LocalMux I__3675 (
            .O(N__15943),
            .I(N__15925));
    Span4Mux_h I__3674 (
            .O(N__15940),
            .I(N__15920));
    Span4Mux_v I__3673 (
            .O(N__15933),
            .I(N__15920));
    Span4Mux_v I__3672 (
            .O(N__15928),
            .I(N__15917));
    Sp12to4 I__3671 (
            .O(N__15925),
            .I(N__15914));
    Span4Mux_h I__3670 (
            .O(N__15920),
            .I(N__15911));
    Odrv4 I__3669 (
            .O(N__15917),
            .I(\receive_module.n3185 ));
    Odrv12 I__3668 (
            .O(N__15914),
            .I(\receive_module.n3185 ));
    Odrv4 I__3667 (
            .O(N__15911),
            .I(\receive_module.n3185 ));
    InMux I__3666 (
            .O(N__15904),
            .I(N__15901));
    LocalMux I__3665 (
            .O(N__15901),
            .I(N__15898));
    Span12Mux_v I__3664 (
            .O(N__15898),
            .I(N__15895));
    Odrv12 I__3663 (
            .O(N__15895),
            .I(\line_buffer.n757 ));
    InMux I__3662 (
            .O(N__15892),
            .I(N__15889));
    LocalMux I__3661 (
            .O(N__15889),
            .I(N__15886));
    Span4Mux_v I__3660 (
            .O(N__15886),
            .I(N__15883));
    Span4Mux_v I__3659 (
            .O(N__15883),
            .I(N__15880));
    Span4Mux_h I__3658 (
            .O(N__15880),
            .I(N__15877));
    Odrv4 I__3657 (
            .O(N__15877),
            .I(\line_buffer.n749 ));
    InMux I__3656 (
            .O(N__15874),
            .I(N__15871));
    LocalMux I__3655 (
            .O(N__15871),
            .I(N__15868));
    Span4Mux_v I__3654 (
            .O(N__15868),
            .I(N__15865));
    Span4Mux_h I__3653 (
            .O(N__15865),
            .I(N__15862));
    Span4Mux_v I__3652 (
            .O(N__15862),
            .I(N__15859));
    Odrv4 I__3651 (
            .O(N__15859),
            .I(\line_buffer.n685 ));
    InMux I__3650 (
            .O(N__15856),
            .I(N__15853));
    LocalMux I__3649 (
            .O(N__15853),
            .I(N__15850));
    Span12Mux_v I__3648 (
            .O(N__15850),
            .I(N__15847));
    Span12Mux_h I__3647 (
            .O(N__15847),
            .I(N__15844));
    Odrv12 I__3646 (
            .O(N__15844),
            .I(\line_buffer.n693 ));
    CascadeMux I__3645 (
            .O(N__15841),
            .I(\line_buffer.n3155_cascade_ ));
    CascadeMux I__3644 (
            .O(N__15838),
            .I(N__15831));
    InMux I__3643 (
            .O(N__15837),
            .I(N__15827));
    CascadeMux I__3642 (
            .O(N__15836),
            .I(N__15822));
    InMux I__3641 (
            .O(N__15835),
            .I(N__15819));
    InMux I__3640 (
            .O(N__15834),
            .I(N__15814));
    InMux I__3639 (
            .O(N__15831),
            .I(N__15814));
    CascadeMux I__3638 (
            .O(N__15830),
            .I(N__15804));
    LocalMux I__3637 (
            .O(N__15827),
            .I(N__15801));
    InMux I__3636 (
            .O(N__15826),
            .I(N__15794));
    InMux I__3635 (
            .O(N__15825),
            .I(N__15794));
    InMux I__3634 (
            .O(N__15822),
            .I(N__15794));
    LocalMux I__3633 (
            .O(N__15819),
            .I(N__15789));
    LocalMux I__3632 (
            .O(N__15814),
            .I(N__15789));
    InMux I__3631 (
            .O(N__15813),
            .I(N__15786));
    CascadeMux I__3630 (
            .O(N__15812),
            .I(N__15782));
    CascadeMux I__3629 (
            .O(N__15811),
            .I(N__15778));
    CascadeMux I__3628 (
            .O(N__15810),
            .I(N__15773));
    CascadeMux I__3627 (
            .O(N__15809),
            .I(N__15769));
    InMux I__3626 (
            .O(N__15808),
            .I(N__15761));
    InMux I__3625 (
            .O(N__15807),
            .I(N__15761));
    InMux I__3624 (
            .O(N__15804),
            .I(N__15761));
    Span4Mux_h I__3623 (
            .O(N__15801),
            .I(N__15756));
    LocalMux I__3622 (
            .O(N__15794),
            .I(N__15756));
    Span4Mux_h I__3621 (
            .O(N__15789),
            .I(N__15751));
    LocalMux I__3620 (
            .O(N__15786),
            .I(N__15751));
    InMux I__3619 (
            .O(N__15785),
            .I(N__15746));
    InMux I__3618 (
            .O(N__15782),
            .I(N__15746));
    CascadeMux I__3617 (
            .O(N__15781),
            .I(N__15742));
    InMux I__3616 (
            .O(N__15778),
            .I(N__15739));
    InMux I__3615 (
            .O(N__15777),
            .I(N__15736));
    InMux I__3614 (
            .O(N__15776),
            .I(N__15733));
    InMux I__3613 (
            .O(N__15773),
            .I(N__15730));
    InMux I__3612 (
            .O(N__15772),
            .I(N__15727));
    InMux I__3611 (
            .O(N__15769),
            .I(N__15724));
    CascadeMux I__3610 (
            .O(N__15768),
            .I(N__15720));
    LocalMux I__3609 (
            .O(N__15761),
            .I(N__15716));
    Span4Mux_h I__3608 (
            .O(N__15756),
            .I(N__15713));
    Span4Mux_v I__3607 (
            .O(N__15751),
            .I(N__15708));
    LocalMux I__3606 (
            .O(N__15746),
            .I(N__15708));
    InMux I__3605 (
            .O(N__15745),
            .I(N__15703));
    InMux I__3604 (
            .O(N__15742),
            .I(N__15703));
    LocalMux I__3603 (
            .O(N__15739),
            .I(N__15700));
    LocalMux I__3602 (
            .O(N__15736),
            .I(N__15697));
    LocalMux I__3601 (
            .O(N__15733),
            .I(N__15694));
    LocalMux I__3600 (
            .O(N__15730),
            .I(N__15691));
    LocalMux I__3599 (
            .O(N__15727),
            .I(N__15686));
    LocalMux I__3598 (
            .O(N__15724),
            .I(N__15686));
    InMux I__3597 (
            .O(N__15723),
            .I(N__15683));
    InMux I__3596 (
            .O(N__15720),
            .I(N__15680));
    InMux I__3595 (
            .O(N__15719),
            .I(N__15677));
    Span4Mux_h I__3594 (
            .O(N__15716),
            .I(N__15670));
    Span4Mux_v I__3593 (
            .O(N__15713),
            .I(N__15670));
    Span4Mux_h I__3592 (
            .O(N__15708),
            .I(N__15670));
    LocalMux I__3591 (
            .O(N__15703),
            .I(N__15665));
    Span12Mux_v I__3590 (
            .O(N__15700),
            .I(N__15665));
    Span4Mux_h I__3589 (
            .O(N__15697),
            .I(N__15656));
    Span4Mux_h I__3588 (
            .O(N__15694),
            .I(N__15656));
    Span4Mux_v I__3587 (
            .O(N__15691),
            .I(N__15656));
    Span4Mux_h I__3586 (
            .O(N__15686),
            .I(N__15656));
    LocalMux I__3585 (
            .O(N__15683),
            .I(TX_ADDR_12));
    LocalMux I__3584 (
            .O(N__15680),
            .I(TX_ADDR_12));
    LocalMux I__3583 (
            .O(N__15677),
            .I(TX_ADDR_12));
    Odrv4 I__3582 (
            .O(N__15670),
            .I(TX_ADDR_12));
    Odrv12 I__3581 (
            .O(N__15665),
            .I(TX_ADDR_12));
    Odrv4 I__3580 (
            .O(N__15656),
            .I(TX_ADDR_12));
    InMux I__3579 (
            .O(N__15643),
            .I(N__15640));
    LocalMux I__3578 (
            .O(N__15640),
            .I(\line_buffer.n3158 ));
    InMux I__3577 (
            .O(N__15637),
            .I(N__15634));
    LocalMux I__3576 (
            .O(N__15634),
            .I(N__15631));
    Span4Mux_h I__3575 (
            .O(N__15631),
            .I(N__15628));
    Span4Mux_h I__3574 (
            .O(N__15628),
            .I(N__15625));
    Odrv4 I__3573 (
            .O(N__15625),
            .I(\line_buffer.n627 ));
    InMux I__3572 (
            .O(N__15622),
            .I(N__15619));
    LocalMux I__3571 (
            .O(N__15619),
            .I(N__15616));
    Span12Mux_v I__3570 (
            .O(N__15616),
            .I(N__15613));
    Odrv12 I__3569 (
            .O(N__15613),
            .I(\line_buffer.n619 ));
    InMux I__3568 (
            .O(N__15610),
            .I(N__15607));
    LocalMux I__3567 (
            .O(N__15607),
            .I(N__15604));
    Span4Mux_v I__3566 (
            .O(N__15604),
            .I(N__15601));
    Odrv4 I__3565 (
            .O(N__15601),
            .I(\line_buffer.n3045 ));
    InMux I__3564 (
            .O(N__15598),
            .I(N__15595));
    LocalMux I__3563 (
            .O(N__15595),
            .I(N__15592));
    Sp12to4 I__3562 (
            .O(N__15592),
            .I(N__15589));
    Span12Mux_v I__3561 (
            .O(N__15589),
            .I(N__15586));
    Odrv12 I__3560 (
            .O(N__15586),
            .I(\line_buffer.n725 ));
    InMux I__3559 (
            .O(N__15583),
            .I(N__15580));
    LocalMux I__3558 (
            .O(N__15580),
            .I(N__15577));
    Odrv12 I__3557 (
            .O(N__15577),
            .I(\line_buffer.n717 ));
    InMux I__3556 (
            .O(N__15574),
            .I(N__15571));
    LocalMux I__3555 (
            .O(N__15571),
            .I(\receive_module.n133 ));
    CascadeMux I__3554 (
            .O(N__15568),
            .I(N__15564));
    CascadeMux I__3553 (
            .O(N__15567),
            .I(N__15561));
    CascadeBuf I__3552 (
            .O(N__15564),
            .I(N__15558));
    CascadeBuf I__3551 (
            .O(N__15561),
            .I(N__15555));
    CascadeMux I__3550 (
            .O(N__15558),
            .I(N__15552));
    CascadeMux I__3549 (
            .O(N__15555),
            .I(N__15549));
    CascadeBuf I__3548 (
            .O(N__15552),
            .I(N__15546));
    CascadeBuf I__3547 (
            .O(N__15549),
            .I(N__15543));
    CascadeMux I__3546 (
            .O(N__15546),
            .I(N__15540));
    CascadeMux I__3545 (
            .O(N__15543),
            .I(N__15537));
    CascadeBuf I__3544 (
            .O(N__15540),
            .I(N__15534));
    CascadeBuf I__3543 (
            .O(N__15537),
            .I(N__15531));
    CascadeMux I__3542 (
            .O(N__15534),
            .I(N__15528));
    CascadeMux I__3541 (
            .O(N__15531),
            .I(N__15525));
    CascadeBuf I__3540 (
            .O(N__15528),
            .I(N__15522));
    CascadeBuf I__3539 (
            .O(N__15525),
            .I(N__15519));
    CascadeMux I__3538 (
            .O(N__15522),
            .I(N__15516));
    CascadeMux I__3537 (
            .O(N__15519),
            .I(N__15513));
    CascadeBuf I__3536 (
            .O(N__15516),
            .I(N__15510));
    CascadeBuf I__3535 (
            .O(N__15513),
            .I(N__15507));
    CascadeMux I__3534 (
            .O(N__15510),
            .I(N__15504));
    CascadeMux I__3533 (
            .O(N__15507),
            .I(N__15501));
    CascadeBuf I__3532 (
            .O(N__15504),
            .I(N__15498));
    CascadeBuf I__3531 (
            .O(N__15501),
            .I(N__15495));
    CascadeMux I__3530 (
            .O(N__15498),
            .I(N__15492));
    CascadeMux I__3529 (
            .O(N__15495),
            .I(N__15489));
    CascadeBuf I__3528 (
            .O(N__15492),
            .I(N__15486));
    CascadeBuf I__3527 (
            .O(N__15489),
            .I(N__15483));
    CascadeMux I__3526 (
            .O(N__15486),
            .I(N__15480));
    CascadeMux I__3525 (
            .O(N__15483),
            .I(N__15477));
    CascadeBuf I__3524 (
            .O(N__15480),
            .I(N__15474));
    CascadeBuf I__3523 (
            .O(N__15477),
            .I(N__15471));
    CascadeMux I__3522 (
            .O(N__15474),
            .I(N__15468));
    CascadeMux I__3521 (
            .O(N__15471),
            .I(N__15465));
    CascadeBuf I__3520 (
            .O(N__15468),
            .I(N__15462));
    CascadeBuf I__3519 (
            .O(N__15465),
            .I(N__15459));
    CascadeMux I__3518 (
            .O(N__15462),
            .I(N__15456));
    CascadeMux I__3517 (
            .O(N__15459),
            .I(N__15453));
    CascadeBuf I__3516 (
            .O(N__15456),
            .I(N__15450));
    CascadeBuf I__3515 (
            .O(N__15453),
            .I(N__15447));
    CascadeMux I__3514 (
            .O(N__15450),
            .I(N__15444));
    CascadeMux I__3513 (
            .O(N__15447),
            .I(N__15441));
    CascadeBuf I__3512 (
            .O(N__15444),
            .I(N__15438));
    CascadeBuf I__3511 (
            .O(N__15441),
            .I(N__15435));
    CascadeMux I__3510 (
            .O(N__15438),
            .I(N__15432));
    CascadeMux I__3509 (
            .O(N__15435),
            .I(N__15429));
    CascadeBuf I__3508 (
            .O(N__15432),
            .I(N__15426));
    CascadeBuf I__3507 (
            .O(N__15429),
            .I(N__15423));
    CascadeMux I__3506 (
            .O(N__15426),
            .I(N__15420));
    CascadeMux I__3505 (
            .O(N__15423),
            .I(N__15417));
    CascadeBuf I__3504 (
            .O(N__15420),
            .I(N__15414));
    CascadeBuf I__3503 (
            .O(N__15417),
            .I(N__15411));
    CascadeMux I__3502 (
            .O(N__15414),
            .I(N__15408));
    CascadeMux I__3501 (
            .O(N__15411),
            .I(N__15405));
    CascadeBuf I__3500 (
            .O(N__15408),
            .I(N__15402));
    CascadeBuf I__3499 (
            .O(N__15405),
            .I(N__15399));
    CascadeMux I__3498 (
            .O(N__15402),
            .I(N__15396));
    CascadeMux I__3497 (
            .O(N__15399),
            .I(N__15393));
    CascadeBuf I__3496 (
            .O(N__15396),
            .I(N__15390));
    CascadeBuf I__3495 (
            .O(N__15393),
            .I(N__15387));
    CascadeMux I__3494 (
            .O(N__15390),
            .I(N__15384));
    CascadeMux I__3493 (
            .O(N__15387),
            .I(N__15381));
    InMux I__3492 (
            .O(N__15384),
            .I(N__15378));
    InMux I__3491 (
            .O(N__15381),
            .I(N__15375));
    LocalMux I__3490 (
            .O(N__15378),
            .I(N__15372));
    LocalMux I__3489 (
            .O(N__15375),
            .I(N__15369));
    Span4Mux_v I__3488 (
            .O(N__15372),
            .I(N__15366));
    Span4Mux_v I__3487 (
            .O(N__15369),
            .I(N__15363));
    Sp12to4 I__3486 (
            .O(N__15366),
            .I(N__15360));
    Sp12to4 I__3485 (
            .O(N__15363),
            .I(N__15357));
    Span12Mux_h I__3484 (
            .O(N__15360),
            .I(N__15350));
    Span12Mux_h I__3483 (
            .O(N__15357),
            .I(N__15350));
    InMux I__3482 (
            .O(N__15356),
            .I(N__15347));
    InMux I__3481 (
            .O(N__15355),
            .I(N__15344));
    Span12Mux_v I__3480 (
            .O(N__15350),
            .I(N__15341));
    LocalMux I__3479 (
            .O(N__15347),
            .I(RX_ADDR_3));
    LocalMux I__3478 (
            .O(N__15344),
            .I(RX_ADDR_3));
    Odrv12 I__3477 (
            .O(N__15341),
            .I(RX_ADDR_3));
    CascadeMux I__3476 (
            .O(N__15334),
            .I(N__15331));
    InMux I__3475 (
            .O(N__15331),
            .I(N__15328));
    LocalMux I__3474 (
            .O(N__15328),
            .I(\receive_module.n134 ));
    CascadeMux I__3473 (
            .O(N__15325),
            .I(N__15322));
    CascadeBuf I__3472 (
            .O(N__15322),
            .I(N__15318));
    CascadeMux I__3471 (
            .O(N__15321),
            .I(N__15315));
    CascadeMux I__3470 (
            .O(N__15318),
            .I(N__15312));
    CascadeBuf I__3469 (
            .O(N__15315),
            .I(N__15309));
    CascadeBuf I__3468 (
            .O(N__15312),
            .I(N__15306));
    CascadeMux I__3467 (
            .O(N__15309),
            .I(N__15303));
    CascadeMux I__3466 (
            .O(N__15306),
            .I(N__15300));
    CascadeBuf I__3465 (
            .O(N__15303),
            .I(N__15297));
    CascadeBuf I__3464 (
            .O(N__15300),
            .I(N__15294));
    CascadeMux I__3463 (
            .O(N__15297),
            .I(N__15291));
    CascadeMux I__3462 (
            .O(N__15294),
            .I(N__15288));
    CascadeBuf I__3461 (
            .O(N__15291),
            .I(N__15285));
    CascadeBuf I__3460 (
            .O(N__15288),
            .I(N__15282));
    CascadeMux I__3459 (
            .O(N__15285),
            .I(N__15279));
    CascadeMux I__3458 (
            .O(N__15282),
            .I(N__15276));
    CascadeBuf I__3457 (
            .O(N__15279),
            .I(N__15273));
    CascadeBuf I__3456 (
            .O(N__15276),
            .I(N__15270));
    CascadeMux I__3455 (
            .O(N__15273),
            .I(N__15267));
    CascadeMux I__3454 (
            .O(N__15270),
            .I(N__15264));
    CascadeBuf I__3453 (
            .O(N__15267),
            .I(N__15261));
    CascadeBuf I__3452 (
            .O(N__15264),
            .I(N__15258));
    CascadeMux I__3451 (
            .O(N__15261),
            .I(N__15255));
    CascadeMux I__3450 (
            .O(N__15258),
            .I(N__15252));
    CascadeBuf I__3449 (
            .O(N__15255),
            .I(N__15249));
    CascadeBuf I__3448 (
            .O(N__15252),
            .I(N__15246));
    CascadeMux I__3447 (
            .O(N__15249),
            .I(N__15243));
    CascadeMux I__3446 (
            .O(N__15246),
            .I(N__15240));
    CascadeBuf I__3445 (
            .O(N__15243),
            .I(N__15237));
    CascadeBuf I__3444 (
            .O(N__15240),
            .I(N__15234));
    CascadeMux I__3443 (
            .O(N__15237),
            .I(N__15231));
    CascadeMux I__3442 (
            .O(N__15234),
            .I(N__15228));
    CascadeBuf I__3441 (
            .O(N__15231),
            .I(N__15225));
    CascadeBuf I__3440 (
            .O(N__15228),
            .I(N__15222));
    CascadeMux I__3439 (
            .O(N__15225),
            .I(N__15219));
    CascadeMux I__3438 (
            .O(N__15222),
            .I(N__15216));
    CascadeBuf I__3437 (
            .O(N__15219),
            .I(N__15213));
    CascadeBuf I__3436 (
            .O(N__15216),
            .I(N__15210));
    CascadeMux I__3435 (
            .O(N__15213),
            .I(N__15207));
    CascadeMux I__3434 (
            .O(N__15210),
            .I(N__15204));
    CascadeBuf I__3433 (
            .O(N__15207),
            .I(N__15201));
    CascadeBuf I__3432 (
            .O(N__15204),
            .I(N__15198));
    CascadeMux I__3431 (
            .O(N__15201),
            .I(N__15195));
    CascadeMux I__3430 (
            .O(N__15198),
            .I(N__15192));
    CascadeBuf I__3429 (
            .O(N__15195),
            .I(N__15189));
    CascadeBuf I__3428 (
            .O(N__15192),
            .I(N__15186));
    CascadeMux I__3427 (
            .O(N__15189),
            .I(N__15183));
    CascadeMux I__3426 (
            .O(N__15186),
            .I(N__15180));
    CascadeBuf I__3425 (
            .O(N__15183),
            .I(N__15177));
    CascadeBuf I__3424 (
            .O(N__15180),
            .I(N__15174));
    CascadeMux I__3423 (
            .O(N__15177),
            .I(N__15171));
    CascadeMux I__3422 (
            .O(N__15174),
            .I(N__15168));
    CascadeBuf I__3421 (
            .O(N__15171),
            .I(N__15165));
    CascadeBuf I__3420 (
            .O(N__15168),
            .I(N__15162));
    CascadeMux I__3419 (
            .O(N__15165),
            .I(N__15159));
    CascadeMux I__3418 (
            .O(N__15162),
            .I(N__15156));
    CascadeBuf I__3417 (
            .O(N__15159),
            .I(N__15153));
    CascadeBuf I__3416 (
            .O(N__15156),
            .I(N__15150));
    CascadeMux I__3415 (
            .O(N__15153),
            .I(N__15147));
    CascadeMux I__3414 (
            .O(N__15150),
            .I(N__15144));
    CascadeBuf I__3413 (
            .O(N__15147),
            .I(N__15141));
    InMux I__3412 (
            .O(N__15144),
            .I(N__15138));
    CascadeMux I__3411 (
            .O(N__15141),
            .I(N__15135));
    LocalMux I__3410 (
            .O(N__15138),
            .I(N__15132));
    InMux I__3409 (
            .O(N__15135),
            .I(N__15129));
    Span4Mux_s3_v I__3408 (
            .O(N__15132),
            .I(N__15126));
    LocalMux I__3407 (
            .O(N__15129),
            .I(N__15123));
    Sp12to4 I__3406 (
            .O(N__15126),
            .I(N__15120));
    Span12Mux_s5_v I__3405 (
            .O(N__15123),
            .I(N__15115));
    Span12Mux_h I__3404 (
            .O(N__15120),
            .I(N__15112));
    InMux I__3403 (
            .O(N__15119),
            .I(N__15109));
    InMux I__3402 (
            .O(N__15118),
            .I(N__15106));
    Span12Mux_v I__3401 (
            .O(N__15115),
            .I(N__15103));
    Span12Mux_v I__3400 (
            .O(N__15112),
            .I(N__15100));
    LocalMux I__3399 (
            .O(N__15109),
            .I(RX_ADDR_2));
    LocalMux I__3398 (
            .O(N__15106),
            .I(RX_ADDR_2));
    Odrv12 I__3397 (
            .O(N__15103),
            .I(RX_ADDR_2));
    Odrv12 I__3396 (
            .O(N__15100),
            .I(RX_ADDR_2));
    InMux I__3395 (
            .O(N__15091),
            .I(N__15088));
    LocalMux I__3394 (
            .O(N__15088),
            .I(\receive_module.n135 ));
    CascadeMux I__3393 (
            .O(N__15085),
            .I(N__15081));
    CascadeMux I__3392 (
            .O(N__15084),
            .I(N__15078));
    CascadeBuf I__3391 (
            .O(N__15081),
            .I(N__15075));
    CascadeBuf I__3390 (
            .O(N__15078),
            .I(N__15072));
    CascadeMux I__3389 (
            .O(N__15075),
            .I(N__15069));
    CascadeMux I__3388 (
            .O(N__15072),
            .I(N__15066));
    CascadeBuf I__3387 (
            .O(N__15069),
            .I(N__15063));
    CascadeBuf I__3386 (
            .O(N__15066),
            .I(N__15060));
    CascadeMux I__3385 (
            .O(N__15063),
            .I(N__15057));
    CascadeMux I__3384 (
            .O(N__15060),
            .I(N__15054));
    CascadeBuf I__3383 (
            .O(N__15057),
            .I(N__15051));
    CascadeBuf I__3382 (
            .O(N__15054),
            .I(N__15048));
    CascadeMux I__3381 (
            .O(N__15051),
            .I(N__15045));
    CascadeMux I__3380 (
            .O(N__15048),
            .I(N__15042));
    CascadeBuf I__3379 (
            .O(N__15045),
            .I(N__15039));
    CascadeBuf I__3378 (
            .O(N__15042),
            .I(N__15036));
    CascadeMux I__3377 (
            .O(N__15039),
            .I(N__15033));
    CascadeMux I__3376 (
            .O(N__15036),
            .I(N__15030));
    CascadeBuf I__3375 (
            .O(N__15033),
            .I(N__15027));
    CascadeBuf I__3374 (
            .O(N__15030),
            .I(N__15024));
    CascadeMux I__3373 (
            .O(N__15027),
            .I(N__15021));
    CascadeMux I__3372 (
            .O(N__15024),
            .I(N__15018));
    CascadeBuf I__3371 (
            .O(N__15021),
            .I(N__15015));
    CascadeBuf I__3370 (
            .O(N__15018),
            .I(N__15012));
    CascadeMux I__3369 (
            .O(N__15015),
            .I(N__15009));
    CascadeMux I__3368 (
            .O(N__15012),
            .I(N__15006));
    CascadeBuf I__3367 (
            .O(N__15009),
            .I(N__15003));
    CascadeBuf I__3366 (
            .O(N__15006),
            .I(N__15000));
    CascadeMux I__3365 (
            .O(N__15003),
            .I(N__14997));
    CascadeMux I__3364 (
            .O(N__15000),
            .I(N__14994));
    CascadeBuf I__3363 (
            .O(N__14997),
            .I(N__14991));
    CascadeBuf I__3362 (
            .O(N__14994),
            .I(N__14988));
    CascadeMux I__3361 (
            .O(N__14991),
            .I(N__14985));
    CascadeMux I__3360 (
            .O(N__14988),
            .I(N__14982));
    CascadeBuf I__3359 (
            .O(N__14985),
            .I(N__14979));
    CascadeBuf I__3358 (
            .O(N__14982),
            .I(N__14976));
    CascadeMux I__3357 (
            .O(N__14979),
            .I(N__14973));
    CascadeMux I__3356 (
            .O(N__14976),
            .I(N__14970));
    CascadeBuf I__3355 (
            .O(N__14973),
            .I(N__14967));
    CascadeBuf I__3354 (
            .O(N__14970),
            .I(N__14964));
    CascadeMux I__3353 (
            .O(N__14967),
            .I(N__14961));
    CascadeMux I__3352 (
            .O(N__14964),
            .I(N__14958));
    CascadeBuf I__3351 (
            .O(N__14961),
            .I(N__14955));
    CascadeBuf I__3350 (
            .O(N__14958),
            .I(N__14952));
    CascadeMux I__3349 (
            .O(N__14955),
            .I(N__14949));
    CascadeMux I__3348 (
            .O(N__14952),
            .I(N__14946));
    CascadeBuf I__3347 (
            .O(N__14949),
            .I(N__14943));
    CascadeBuf I__3346 (
            .O(N__14946),
            .I(N__14940));
    CascadeMux I__3345 (
            .O(N__14943),
            .I(N__14937));
    CascadeMux I__3344 (
            .O(N__14940),
            .I(N__14934));
    CascadeBuf I__3343 (
            .O(N__14937),
            .I(N__14931));
    CascadeBuf I__3342 (
            .O(N__14934),
            .I(N__14928));
    CascadeMux I__3341 (
            .O(N__14931),
            .I(N__14925));
    CascadeMux I__3340 (
            .O(N__14928),
            .I(N__14922));
    CascadeBuf I__3339 (
            .O(N__14925),
            .I(N__14919));
    CascadeBuf I__3338 (
            .O(N__14922),
            .I(N__14916));
    CascadeMux I__3337 (
            .O(N__14919),
            .I(N__14913));
    CascadeMux I__3336 (
            .O(N__14916),
            .I(N__14910));
    CascadeBuf I__3335 (
            .O(N__14913),
            .I(N__14907));
    CascadeBuf I__3334 (
            .O(N__14910),
            .I(N__14904));
    CascadeMux I__3333 (
            .O(N__14907),
            .I(N__14901));
    CascadeMux I__3332 (
            .O(N__14904),
            .I(N__14898));
    InMux I__3331 (
            .O(N__14901),
            .I(N__14895));
    InMux I__3330 (
            .O(N__14898),
            .I(N__14892));
    LocalMux I__3329 (
            .O(N__14895),
            .I(N__14889));
    LocalMux I__3328 (
            .O(N__14892),
            .I(N__14886));
    Span4Mux_h I__3327 (
            .O(N__14889),
            .I(N__14883));
    Span4Mux_h I__3326 (
            .O(N__14886),
            .I(N__14880));
    Sp12to4 I__3325 (
            .O(N__14883),
            .I(N__14877));
    Sp12to4 I__3324 (
            .O(N__14880),
            .I(N__14874));
    Span12Mux_s5_v I__3323 (
            .O(N__14877),
            .I(N__14869));
    Span12Mux_s5_v I__3322 (
            .O(N__14874),
            .I(N__14866));
    InMux I__3321 (
            .O(N__14873),
            .I(N__14863));
    InMux I__3320 (
            .O(N__14872),
            .I(N__14860));
    Span12Mux_v I__3319 (
            .O(N__14869),
            .I(N__14855));
    Span12Mux_v I__3318 (
            .O(N__14866),
            .I(N__14855));
    LocalMux I__3317 (
            .O(N__14863),
            .I(RX_ADDR_1));
    LocalMux I__3316 (
            .O(N__14860),
            .I(RX_ADDR_1));
    Odrv12 I__3315 (
            .O(N__14855),
            .I(RX_ADDR_1));
    InMux I__3314 (
            .O(N__14848),
            .I(N__14845));
    LocalMux I__3313 (
            .O(N__14845),
            .I(N__14842));
    Span4Mux_h I__3312 (
            .O(N__14842),
            .I(N__14839));
    Span4Mux_h I__3311 (
            .O(N__14839),
            .I(N__14836));
    Odrv4 I__3310 (
            .O(N__14836),
            .I(\line_buffer.n628 ));
    CascadeMux I__3309 (
            .O(N__14833),
            .I(N__14830));
    InMux I__3308 (
            .O(N__14830),
            .I(N__14827));
    LocalMux I__3307 (
            .O(N__14827),
            .I(N__14824));
    Span12Mux_h I__3306 (
            .O(N__14824),
            .I(N__14821));
    Span12Mux_v I__3305 (
            .O(N__14821),
            .I(N__14818));
    Odrv12 I__3304 (
            .O(N__14818),
            .I(\line_buffer.n620 ));
    InMux I__3303 (
            .O(N__14815),
            .I(N__14812));
    LocalMux I__3302 (
            .O(N__14812),
            .I(N__14809));
    Odrv12 I__3301 (
            .O(N__14809),
            .I(\line_buffer.n3149 ));
    CascadeMux I__3300 (
            .O(N__14806),
            .I(\line_buffer.n3152_cascade_ ));
    InMux I__3299 (
            .O(N__14803),
            .I(N__14800));
    LocalMux I__3298 (
            .O(N__14800),
            .I(N__14797));
    Span4Mux_h I__3297 (
            .O(N__14797),
            .I(N__14794));
    Odrv4 I__3296 (
            .O(N__14794),
            .I(TX_DATA_5));
    InMux I__3295 (
            .O(N__14791),
            .I(N__14788));
    LocalMux I__3294 (
            .O(N__14788),
            .I(N__14785));
    Span12Mux_v I__3293 (
            .O(N__14785),
            .I(N__14782));
    Odrv12 I__3292 (
            .O(N__14782),
            .I(\line_buffer.n692 ));
    InMux I__3291 (
            .O(N__14779),
            .I(N__14776));
    LocalMux I__3290 (
            .O(N__14776),
            .I(N__14773));
    Span4Mux_v I__3289 (
            .O(N__14773),
            .I(N__14770));
    Span4Mux_h I__3288 (
            .O(N__14770),
            .I(N__14767));
    Odrv4 I__3287 (
            .O(N__14767),
            .I(\line_buffer.n684 ));
    InMux I__3286 (
            .O(N__14764),
            .I(N__14761));
    LocalMux I__3285 (
            .O(N__14761),
            .I(N__14758));
    Span4Mux_v I__3284 (
            .O(N__14758),
            .I(N__14755));
    Odrv4 I__3283 (
            .O(N__14755),
            .I(\line_buffer.n3024 ));
    CascadeMux I__3282 (
            .O(N__14752),
            .I(\line_buffer.n3131_cascade_ ));
    CascadeMux I__3281 (
            .O(N__14749),
            .I(N__14745));
    CascadeMux I__3280 (
            .O(N__14748),
            .I(N__14742));
    CascadeBuf I__3279 (
            .O(N__14745),
            .I(N__14739));
    CascadeBuf I__3278 (
            .O(N__14742),
            .I(N__14736));
    CascadeMux I__3277 (
            .O(N__14739),
            .I(N__14733));
    CascadeMux I__3276 (
            .O(N__14736),
            .I(N__14730));
    CascadeBuf I__3275 (
            .O(N__14733),
            .I(N__14727));
    CascadeBuf I__3274 (
            .O(N__14730),
            .I(N__14724));
    CascadeMux I__3273 (
            .O(N__14727),
            .I(N__14721));
    CascadeMux I__3272 (
            .O(N__14724),
            .I(N__14718));
    CascadeBuf I__3271 (
            .O(N__14721),
            .I(N__14715));
    CascadeBuf I__3270 (
            .O(N__14718),
            .I(N__14712));
    CascadeMux I__3269 (
            .O(N__14715),
            .I(N__14709));
    CascadeMux I__3268 (
            .O(N__14712),
            .I(N__14706));
    CascadeBuf I__3267 (
            .O(N__14709),
            .I(N__14703));
    CascadeBuf I__3266 (
            .O(N__14706),
            .I(N__14700));
    CascadeMux I__3265 (
            .O(N__14703),
            .I(N__14697));
    CascadeMux I__3264 (
            .O(N__14700),
            .I(N__14694));
    CascadeBuf I__3263 (
            .O(N__14697),
            .I(N__14691));
    CascadeBuf I__3262 (
            .O(N__14694),
            .I(N__14688));
    CascadeMux I__3261 (
            .O(N__14691),
            .I(N__14685));
    CascadeMux I__3260 (
            .O(N__14688),
            .I(N__14682));
    CascadeBuf I__3259 (
            .O(N__14685),
            .I(N__14679));
    CascadeBuf I__3258 (
            .O(N__14682),
            .I(N__14676));
    CascadeMux I__3257 (
            .O(N__14679),
            .I(N__14673));
    CascadeMux I__3256 (
            .O(N__14676),
            .I(N__14670));
    CascadeBuf I__3255 (
            .O(N__14673),
            .I(N__14667));
    CascadeBuf I__3254 (
            .O(N__14670),
            .I(N__14664));
    CascadeMux I__3253 (
            .O(N__14667),
            .I(N__14661));
    CascadeMux I__3252 (
            .O(N__14664),
            .I(N__14658));
    CascadeBuf I__3251 (
            .O(N__14661),
            .I(N__14655));
    CascadeBuf I__3250 (
            .O(N__14658),
            .I(N__14652));
    CascadeMux I__3249 (
            .O(N__14655),
            .I(N__14649));
    CascadeMux I__3248 (
            .O(N__14652),
            .I(N__14646));
    CascadeBuf I__3247 (
            .O(N__14649),
            .I(N__14643));
    CascadeBuf I__3246 (
            .O(N__14646),
            .I(N__14640));
    CascadeMux I__3245 (
            .O(N__14643),
            .I(N__14637));
    CascadeMux I__3244 (
            .O(N__14640),
            .I(N__14634));
    CascadeBuf I__3243 (
            .O(N__14637),
            .I(N__14631));
    CascadeBuf I__3242 (
            .O(N__14634),
            .I(N__14628));
    CascadeMux I__3241 (
            .O(N__14631),
            .I(N__14625));
    CascadeMux I__3240 (
            .O(N__14628),
            .I(N__14622));
    CascadeBuf I__3239 (
            .O(N__14625),
            .I(N__14619));
    CascadeBuf I__3238 (
            .O(N__14622),
            .I(N__14616));
    CascadeMux I__3237 (
            .O(N__14619),
            .I(N__14613));
    CascadeMux I__3236 (
            .O(N__14616),
            .I(N__14610));
    CascadeBuf I__3235 (
            .O(N__14613),
            .I(N__14607));
    CascadeBuf I__3234 (
            .O(N__14610),
            .I(N__14604));
    CascadeMux I__3233 (
            .O(N__14607),
            .I(N__14601));
    CascadeMux I__3232 (
            .O(N__14604),
            .I(N__14598));
    CascadeBuf I__3231 (
            .O(N__14601),
            .I(N__14595));
    CascadeBuf I__3230 (
            .O(N__14598),
            .I(N__14592));
    CascadeMux I__3229 (
            .O(N__14595),
            .I(N__14589));
    CascadeMux I__3228 (
            .O(N__14592),
            .I(N__14586));
    CascadeBuf I__3227 (
            .O(N__14589),
            .I(N__14583));
    CascadeBuf I__3226 (
            .O(N__14586),
            .I(N__14580));
    CascadeMux I__3225 (
            .O(N__14583),
            .I(N__14577));
    CascadeMux I__3224 (
            .O(N__14580),
            .I(N__14574));
    CascadeBuf I__3223 (
            .O(N__14577),
            .I(N__14571));
    CascadeBuf I__3222 (
            .O(N__14574),
            .I(N__14568));
    CascadeMux I__3221 (
            .O(N__14571),
            .I(N__14565));
    CascadeMux I__3220 (
            .O(N__14568),
            .I(N__14562));
    InMux I__3219 (
            .O(N__14565),
            .I(N__14559));
    InMux I__3218 (
            .O(N__14562),
            .I(N__14556));
    LocalMux I__3217 (
            .O(N__14559),
            .I(N__14553));
    LocalMux I__3216 (
            .O(N__14556),
            .I(N__14550));
    Span4Mux_s1_v I__3215 (
            .O(N__14553),
            .I(N__14547));
    Span4Mux_s1_v I__3214 (
            .O(N__14550),
            .I(N__14544));
    Span4Mux_v I__3213 (
            .O(N__14547),
            .I(N__14541));
    Span4Mux_v I__3212 (
            .O(N__14544),
            .I(N__14538));
    Sp12to4 I__3211 (
            .O(N__14541),
            .I(N__14535));
    Sp12to4 I__3210 (
            .O(N__14538),
            .I(N__14532));
    Span12Mux_s9_h I__3209 (
            .O(N__14535),
            .I(N__14527));
    Span12Mux_s10_h I__3208 (
            .O(N__14532),
            .I(N__14524));
    InMux I__3207 (
            .O(N__14531),
            .I(N__14521));
    InMux I__3206 (
            .O(N__14530),
            .I(N__14518));
    Span12Mux_v I__3205 (
            .O(N__14527),
            .I(N__14513));
    Span12Mux_v I__3204 (
            .O(N__14524),
            .I(N__14513));
    LocalMux I__3203 (
            .O(N__14521),
            .I(RX_ADDR_9));
    LocalMux I__3202 (
            .O(N__14518),
            .I(RX_ADDR_9));
    Odrv12 I__3201 (
            .O(N__14513),
            .I(RX_ADDR_9));
    CascadeMux I__3200 (
            .O(N__14506),
            .I(N__14503));
    InMux I__3199 (
            .O(N__14503),
            .I(N__14500));
    LocalMux I__3198 (
            .O(N__14500),
            .I(\receive_module.n127 ));
    InMux I__3197 (
            .O(N__14497),
            .I(\receive_module.n2735 ));
    InMux I__3196 (
            .O(N__14494),
            .I(\receive_module.n2736 ));
    InMux I__3195 (
            .O(N__14491),
            .I(\receive_module.n2737 ));
    InMux I__3194 (
            .O(N__14488),
            .I(\receive_module.n2738 ));
    InMux I__3193 (
            .O(N__14485),
            .I(\receive_module.n2739 ));
    CEMux I__3192 (
            .O(N__14482),
            .I(N__14479));
    LocalMux I__3191 (
            .O(N__14479),
            .I(N__14476));
    Span4Mux_v I__3190 (
            .O(N__14476),
            .I(N__14473));
    Odrv4 I__3189 (
            .O(N__14473),
            .I(\receive_module.n3181 ));
    InMux I__3188 (
            .O(N__14470),
            .I(N__14467));
    LocalMux I__3187 (
            .O(N__14467),
            .I(N__14463));
    InMux I__3186 (
            .O(N__14466),
            .I(N__14460));
    Span4Mux_h I__3185 (
            .O(N__14463),
            .I(N__14457));
    LocalMux I__3184 (
            .O(N__14460),
            .I(\transmit_module.n388 ));
    Odrv4 I__3183 (
            .O(N__14457),
            .I(\transmit_module.n388 ));
    IoInMux I__3182 (
            .O(N__14452),
            .I(N__14449));
    LocalMux I__3181 (
            .O(N__14449),
            .I(N__14446));
    IoSpan4Mux I__3180 (
            .O(N__14446),
            .I(N__14437));
    SRMux I__3179 (
            .O(N__14445),
            .I(N__14431));
    CascadeMux I__3178 (
            .O(N__14444),
            .I(N__14428));
    CascadeMux I__3177 (
            .O(N__14443),
            .I(N__14420));
    CascadeMux I__3176 (
            .O(N__14442),
            .I(N__14417));
    CascadeMux I__3175 (
            .O(N__14441),
            .I(N__14414));
    SRMux I__3174 (
            .O(N__14440),
            .I(N__14408));
    Span4Mux_s3_h I__3173 (
            .O(N__14437),
            .I(N__14405));
    CascadeMux I__3172 (
            .O(N__14436),
            .I(N__14399));
    CascadeMux I__3171 (
            .O(N__14435),
            .I(N__14394));
    CascadeMux I__3170 (
            .O(N__14434),
            .I(N__14391));
    LocalMux I__3169 (
            .O(N__14431),
            .I(N__14388));
    InMux I__3168 (
            .O(N__14428),
            .I(N__14385));
    CascadeMux I__3167 (
            .O(N__14427),
            .I(N__14381));
    CascadeMux I__3166 (
            .O(N__14426),
            .I(N__14378));
    CascadeMux I__3165 (
            .O(N__14425),
            .I(N__14375));
    CascadeMux I__3164 (
            .O(N__14424),
            .I(N__14372));
    InMux I__3163 (
            .O(N__14423),
            .I(N__14369));
    InMux I__3162 (
            .O(N__14420),
            .I(N__14362));
    InMux I__3161 (
            .O(N__14417),
            .I(N__14362));
    InMux I__3160 (
            .O(N__14414),
            .I(N__14362));
    SRMux I__3159 (
            .O(N__14413),
            .I(N__14357));
    InMux I__3158 (
            .O(N__14412),
            .I(N__14352));
    InMux I__3157 (
            .O(N__14411),
            .I(N__14352));
    LocalMux I__3156 (
            .O(N__14408),
            .I(N__14349));
    Span4Mux_h I__3155 (
            .O(N__14405),
            .I(N__14345));
    SRMux I__3154 (
            .O(N__14404),
            .I(N__14342));
    InMux I__3153 (
            .O(N__14403),
            .I(N__14335));
    InMux I__3152 (
            .O(N__14402),
            .I(N__14335));
    InMux I__3151 (
            .O(N__14399),
            .I(N__14335));
    InMux I__3150 (
            .O(N__14398),
            .I(N__14332));
    InMux I__3149 (
            .O(N__14397),
            .I(N__14325));
    InMux I__3148 (
            .O(N__14394),
            .I(N__14325));
    InMux I__3147 (
            .O(N__14391),
            .I(N__14325));
    Span4Mux_v I__3146 (
            .O(N__14388),
            .I(N__14320));
    LocalMux I__3145 (
            .O(N__14385),
            .I(N__14320));
    InMux I__3144 (
            .O(N__14384),
            .I(N__14311));
    InMux I__3143 (
            .O(N__14381),
            .I(N__14311));
    InMux I__3142 (
            .O(N__14378),
            .I(N__14311));
    InMux I__3141 (
            .O(N__14375),
            .I(N__14311));
    InMux I__3140 (
            .O(N__14372),
            .I(N__14308));
    LocalMux I__3139 (
            .O(N__14369),
            .I(N__14303));
    LocalMux I__3138 (
            .O(N__14362),
            .I(N__14303));
    CascadeMux I__3137 (
            .O(N__14361),
            .I(N__14300));
    CascadeMux I__3136 (
            .O(N__14360),
            .I(N__14297));
    LocalMux I__3135 (
            .O(N__14357),
            .I(N__14293));
    LocalMux I__3134 (
            .O(N__14352),
            .I(N__14290));
    Span4Mux_v I__3133 (
            .O(N__14349),
            .I(N__14287));
    InMux I__3132 (
            .O(N__14348),
            .I(N__14284));
    Span4Mux_h I__3131 (
            .O(N__14345),
            .I(N__14279));
    LocalMux I__3130 (
            .O(N__14342),
            .I(N__14279));
    LocalMux I__3129 (
            .O(N__14335),
            .I(N__14264));
    LocalMux I__3128 (
            .O(N__14332),
            .I(N__14264));
    LocalMux I__3127 (
            .O(N__14325),
            .I(N__14264));
    Span4Mux_v I__3126 (
            .O(N__14320),
            .I(N__14264));
    LocalMux I__3125 (
            .O(N__14311),
            .I(N__14264));
    LocalMux I__3124 (
            .O(N__14308),
            .I(N__14264));
    Span4Mux_h I__3123 (
            .O(N__14303),
            .I(N__14264));
    InMux I__3122 (
            .O(N__14300),
            .I(N__14257));
    InMux I__3121 (
            .O(N__14297),
            .I(N__14257));
    InMux I__3120 (
            .O(N__14296),
            .I(N__14257));
    Span4Mux_h I__3119 (
            .O(N__14293),
            .I(N__14254));
    Span4Mux_v I__3118 (
            .O(N__14290),
            .I(N__14247));
    Span4Mux_h I__3117 (
            .O(N__14287),
            .I(N__14247));
    LocalMux I__3116 (
            .O(N__14284),
            .I(N__14247));
    Span4Mux_v I__3115 (
            .O(N__14279),
            .I(N__14242));
    Span4Mux_v I__3114 (
            .O(N__14264),
            .I(N__14242));
    LocalMux I__3113 (
            .O(N__14257),
            .I(ADV_VSYNC_c));
    Odrv4 I__3112 (
            .O(N__14254),
            .I(ADV_VSYNC_c));
    Odrv4 I__3111 (
            .O(N__14247),
            .I(ADV_VSYNC_c));
    Odrv4 I__3110 (
            .O(N__14242),
            .I(ADV_VSYNC_c));
    IoInMux I__3109 (
            .O(N__14233),
            .I(N__14230));
    LocalMux I__3108 (
            .O(N__14230),
            .I(N__14226));
    CascadeMux I__3107 (
            .O(N__14229),
            .I(N__14223));
    Span12Mux_s3_h I__3106 (
            .O(N__14226),
            .I(N__14220));
    InMux I__3105 (
            .O(N__14223),
            .I(N__14216));
    Span12Mux_h I__3104 (
            .O(N__14220),
            .I(N__14213));
    CascadeMux I__3103 (
            .O(N__14219),
            .I(N__14210));
    LocalMux I__3102 (
            .O(N__14216),
            .I(N__14207));
    Span12Mux_v I__3101 (
            .O(N__14213),
            .I(N__14203));
    InMux I__3100 (
            .O(N__14210),
            .I(N__14200));
    Span4Mux_v I__3099 (
            .O(N__14207),
            .I(N__14197));
    InMux I__3098 (
            .O(N__14206),
            .I(N__14194));
    Odrv12 I__3097 (
            .O(N__14203),
            .I(DEBUG_c_0));
    LocalMux I__3096 (
            .O(N__14200),
            .I(DEBUG_c_0));
    Odrv4 I__3095 (
            .O(N__14197),
            .I(DEBUG_c_0));
    LocalMux I__3094 (
            .O(N__14194),
            .I(DEBUG_c_0));
    InMux I__3093 (
            .O(N__14185),
            .I(N__14168));
    SRMux I__3092 (
            .O(N__14184),
            .I(N__14161));
    InMux I__3091 (
            .O(N__14183),
            .I(N__14158));
    InMux I__3090 (
            .O(N__14182),
            .I(N__14149));
    InMux I__3089 (
            .O(N__14181),
            .I(N__14149));
    InMux I__3088 (
            .O(N__14180),
            .I(N__14149));
    InMux I__3087 (
            .O(N__14179),
            .I(N__14149));
    InMux I__3086 (
            .O(N__14178),
            .I(N__14142));
    InMux I__3085 (
            .O(N__14177),
            .I(N__14142));
    InMux I__3084 (
            .O(N__14176),
            .I(N__14142));
    InMux I__3083 (
            .O(N__14175),
            .I(N__14132));
    InMux I__3082 (
            .O(N__14174),
            .I(N__14132));
    InMux I__3081 (
            .O(N__14173),
            .I(N__14132));
    InMux I__3080 (
            .O(N__14172),
            .I(N__14125));
    InMux I__3079 (
            .O(N__14171),
            .I(N__14125));
    LocalMux I__3078 (
            .O(N__14168),
            .I(N__14122));
    InMux I__3077 (
            .O(N__14167),
            .I(N__14113));
    InMux I__3076 (
            .O(N__14166),
            .I(N__14113));
    InMux I__3075 (
            .O(N__14165),
            .I(N__14113));
    InMux I__3074 (
            .O(N__14164),
            .I(N__14113));
    LocalMux I__3073 (
            .O(N__14161),
            .I(N__14110));
    LocalMux I__3072 (
            .O(N__14158),
            .I(N__14103));
    LocalMux I__3071 (
            .O(N__14149),
            .I(N__14103));
    LocalMux I__3070 (
            .O(N__14142),
            .I(N__14103));
    InMux I__3069 (
            .O(N__14141),
            .I(N__14096));
    InMux I__3068 (
            .O(N__14140),
            .I(N__14096));
    InMux I__3067 (
            .O(N__14139),
            .I(N__14093));
    LocalMux I__3066 (
            .O(N__14132),
            .I(N__14090));
    InMux I__3065 (
            .O(N__14131),
            .I(N__14087));
    SRMux I__3064 (
            .O(N__14130),
            .I(N__14084));
    LocalMux I__3063 (
            .O(N__14125),
            .I(N__14073));
    Span4Mux_v I__3062 (
            .O(N__14122),
            .I(N__14073));
    LocalMux I__3061 (
            .O(N__14113),
            .I(N__14073));
    Span4Mux_v I__3060 (
            .O(N__14110),
            .I(N__14073));
    Span4Mux_h I__3059 (
            .O(N__14103),
            .I(N__14073));
    SRMux I__3058 (
            .O(N__14102),
            .I(N__14070));
    SRMux I__3057 (
            .O(N__14101),
            .I(N__14067));
    LocalMux I__3056 (
            .O(N__14096),
            .I(VGA_VISIBLE));
    LocalMux I__3055 (
            .O(N__14093),
            .I(VGA_VISIBLE));
    Odrv4 I__3054 (
            .O(N__14090),
            .I(VGA_VISIBLE));
    LocalMux I__3053 (
            .O(N__14087),
            .I(VGA_VISIBLE));
    LocalMux I__3052 (
            .O(N__14084),
            .I(VGA_VISIBLE));
    Odrv4 I__3051 (
            .O(N__14073),
            .I(VGA_VISIBLE));
    LocalMux I__3050 (
            .O(N__14070),
            .I(VGA_VISIBLE));
    LocalMux I__3049 (
            .O(N__14067),
            .I(VGA_VISIBLE));
    CascadeMux I__3048 (
            .O(N__14050),
            .I(N__14046));
    CascadeMux I__3047 (
            .O(N__14049),
            .I(N__14043));
    CascadeBuf I__3046 (
            .O(N__14046),
            .I(N__14040));
    CascadeBuf I__3045 (
            .O(N__14043),
            .I(N__14037));
    CascadeMux I__3044 (
            .O(N__14040),
            .I(N__14034));
    CascadeMux I__3043 (
            .O(N__14037),
            .I(N__14031));
    CascadeBuf I__3042 (
            .O(N__14034),
            .I(N__14028));
    CascadeBuf I__3041 (
            .O(N__14031),
            .I(N__14025));
    CascadeMux I__3040 (
            .O(N__14028),
            .I(N__14022));
    CascadeMux I__3039 (
            .O(N__14025),
            .I(N__14019));
    CascadeBuf I__3038 (
            .O(N__14022),
            .I(N__14016));
    CascadeBuf I__3037 (
            .O(N__14019),
            .I(N__14013));
    CascadeMux I__3036 (
            .O(N__14016),
            .I(N__14010));
    CascadeMux I__3035 (
            .O(N__14013),
            .I(N__14007));
    CascadeBuf I__3034 (
            .O(N__14010),
            .I(N__14004));
    CascadeBuf I__3033 (
            .O(N__14007),
            .I(N__14001));
    CascadeMux I__3032 (
            .O(N__14004),
            .I(N__13998));
    CascadeMux I__3031 (
            .O(N__14001),
            .I(N__13995));
    CascadeBuf I__3030 (
            .O(N__13998),
            .I(N__13992));
    CascadeBuf I__3029 (
            .O(N__13995),
            .I(N__13989));
    CascadeMux I__3028 (
            .O(N__13992),
            .I(N__13986));
    CascadeMux I__3027 (
            .O(N__13989),
            .I(N__13983));
    CascadeBuf I__3026 (
            .O(N__13986),
            .I(N__13980));
    CascadeBuf I__3025 (
            .O(N__13983),
            .I(N__13977));
    CascadeMux I__3024 (
            .O(N__13980),
            .I(N__13974));
    CascadeMux I__3023 (
            .O(N__13977),
            .I(N__13971));
    CascadeBuf I__3022 (
            .O(N__13974),
            .I(N__13968));
    CascadeBuf I__3021 (
            .O(N__13971),
            .I(N__13965));
    CascadeMux I__3020 (
            .O(N__13968),
            .I(N__13962));
    CascadeMux I__3019 (
            .O(N__13965),
            .I(N__13959));
    CascadeBuf I__3018 (
            .O(N__13962),
            .I(N__13956));
    CascadeBuf I__3017 (
            .O(N__13959),
            .I(N__13953));
    CascadeMux I__3016 (
            .O(N__13956),
            .I(N__13950));
    CascadeMux I__3015 (
            .O(N__13953),
            .I(N__13947));
    CascadeBuf I__3014 (
            .O(N__13950),
            .I(N__13944));
    CascadeBuf I__3013 (
            .O(N__13947),
            .I(N__13941));
    CascadeMux I__3012 (
            .O(N__13944),
            .I(N__13938));
    CascadeMux I__3011 (
            .O(N__13941),
            .I(N__13935));
    CascadeBuf I__3010 (
            .O(N__13938),
            .I(N__13932));
    CascadeBuf I__3009 (
            .O(N__13935),
            .I(N__13929));
    CascadeMux I__3008 (
            .O(N__13932),
            .I(N__13926));
    CascadeMux I__3007 (
            .O(N__13929),
            .I(N__13923));
    CascadeBuf I__3006 (
            .O(N__13926),
            .I(N__13920));
    CascadeBuf I__3005 (
            .O(N__13923),
            .I(N__13917));
    CascadeMux I__3004 (
            .O(N__13920),
            .I(N__13914));
    CascadeMux I__3003 (
            .O(N__13917),
            .I(N__13911));
    CascadeBuf I__3002 (
            .O(N__13914),
            .I(N__13908));
    CascadeBuf I__3001 (
            .O(N__13911),
            .I(N__13905));
    CascadeMux I__3000 (
            .O(N__13908),
            .I(N__13902));
    CascadeMux I__2999 (
            .O(N__13905),
            .I(N__13899));
    CascadeBuf I__2998 (
            .O(N__13902),
            .I(N__13896));
    CascadeBuf I__2997 (
            .O(N__13899),
            .I(N__13893));
    CascadeMux I__2996 (
            .O(N__13896),
            .I(N__13890));
    CascadeMux I__2995 (
            .O(N__13893),
            .I(N__13887));
    CascadeBuf I__2994 (
            .O(N__13890),
            .I(N__13884));
    CascadeBuf I__2993 (
            .O(N__13887),
            .I(N__13881));
    CascadeMux I__2992 (
            .O(N__13884),
            .I(N__13878));
    CascadeMux I__2991 (
            .O(N__13881),
            .I(N__13875));
    CascadeBuf I__2990 (
            .O(N__13878),
            .I(N__13872));
    CascadeBuf I__2989 (
            .O(N__13875),
            .I(N__13869));
    CascadeMux I__2988 (
            .O(N__13872),
            .I(N__13866));
    CascadeMux I__2987 (
            .O(N__13869),
            .I(N__13863));
    InMux I__2986 (
            .O(N__13866),
            .I(N__13860));
    InMux I__2985 (
            .O(N__13863),
            .I(N__13857));
    LocalMux I__2984 (
            .O(N__13860),
            .I(N__13854));
    LocalMux I__2983 (
            .O(N__13857),
            .I(N__13851));
    Span12Mux_h I__2982 (
            .O(N__13854),
            .I(N__13848));
    Span12Mux_s11_h I__2981 (
            .O(N__13851),
            .I(N__13845));
    Span12Mux_v I__2980 (
            .O(N__13848),
            .I(N__13842));
    Span12Mux_v I__2979 (
            .O(N__13845),
            .I(N__13839));
    Odrv12 I__2978 (
            .O(N__13842),
            .I(n28));
    Odrv12 I__2977 (
            .O(N__13839),
            .I(n28));
    CascadeMux I__2976 (
            .O(N__13834),
            .I(N__13831));
    InMux I__2975 (
            .O(N__13831),
            .I(N__13828));
    LocalMux I__2974 (
            .O(N__13828),
            .I(N__13825));
    Span4Mux_v I__2973 (
            .O(N__13825),
            .I(N__13822));
    Sp12to4 I__2972 (
            .O(N__13822),
            .I(N__13819));
    Span12Mux_h I__2971 (
            .O(N__13819),
            .I(N__13816));
    Span12Mux_v I__2970 (
            .O(N__13816),
            .I(N__13813));
    Odrv12 I__2969 (
            .O(N__13813),
            .I(\line_buffer.n744 ));
    InMux I__2968 (
            .O(N__13810),
            .I(N__13807));
    LocalMux I__2967 (
            .O(N__13807),
            .I(N__13804));
    Span4Mux_v I__2966 (
            .O(N__13804),
            .I(N__13801));
    Sp12to4 I__2965 (
            .O(N__13801),
            .I(N__13798));
    Odrv12 I__2964 (
            .O(N__13798),
            .I(\line_buffer.n752 ));
    InMux I__2963 (
            .O(N__13795),
            .I(N__13792));
    LocalMux I__2962 (
            .O(N__13792),
            .I(N__13789));
    Span4Mux_v I__2961 (
            .O(N__13789),
            .I(N__13786));
    Odrv4 I__2960 (
            .O(N__13786),
            .I(\line_buffer.n3119 ));
    InMux I__2959 (
            .O(N__13783),
            .I(N__13780));
    LocalMux I__2958 (
            .O(N__13780),
            .I(N__13777));
    Odrv12 I__2957 (
            .O(N__13777),
            .I(\line_buffer.n695 ));
    InMux I__2956 (
            .O(N__13774),
            .I(N__13771));
    LocalMux I__2955 (
            .O(N__13771),
            .I(N__13768));
    Span4Mux_h I__2954 (
            .O(N__13768),
            .I(N__13765));
    Sp12to4 I__2953 (
            .O(N__13765),
            .I(N__13762));
    Span12Mux_v I__2952 (
            .O(N__13762),
            .I(N__13759));
    Span12Mux_v I__2951 (
            .O(N__13759),
            .I(N__13756));
    Odrv12 I__2950 (
            .O(N__13756),
            .I(\line_buffer.n687 ));
    InMux I__2949 (
            .O(N__13753),
            .I(N__13750));
    LocalMux I__2948 (
            .O(N__13750),
            .I(\line_buffer.n3027 ));
    CascadeMux I__2947 (
            .O(N__13747),
            .I(N__13743));
    CascadeMux I__2946 (
            .O(N__13746),
            .I(N__13740));
    CascadeBuf I__2945 (
            .O(N__13743),
            .I(N__13737));
    CascadeBuf I__2944 (
            .O(N__13740),
            .I(N__13734));
    CascadeMux I__2943 (
            .O(N__13737),
            .I(N__13731));
    CascadeMux I__2942 (
            .O(N__13734),
            .I(N__13728));
    CascadeBuf I__2941 (
            .O(N__13731),
            .I(N__13725));
    CascadeBuf I__2940 (
            .O(N__13728),
            .I(N__13722));
    CascadeMux I__2939 (
            .O(N__13725),
            .I(N__13719));
    CascadeMux I__2938 (
            .O(N__13722),
            .I(N__13716));
    CascadeBuf I__2937 (
            .O(N__13719),
            .I(N__13713));
    CascadeBuf I__2936 (
            .O(N__13716),
            .I(N__13710));
    CascadeMux I__2935 (
            .O(N__13713),
            .I(N__13707));
    CascadeMux I__2934 (
            .O(N__13710),
            .I(N__13704));
    CascadeBuf I__2933 (
            .O(N__13707),
            .I(N__13701));
    CascadeBuf I__2932 (
            .O(N__13704),
            .I(N__13698));
    CascadeMux I__2931 (
            .O(N__13701),
            .I(N__13695));
    CascadeMux I__2930 (
            .O(N__13698),
            .I(N__13692));
    CascadeBuf I__2929 (
            .O(N__13695),
            .I(N__13689));
    CascadeBuf I__2928 (
            .O(N__13692),
            .I(N__13686));
    CascadeMux I__2927 (
            .O(N__13689),
            .I(N__13683));
    CascadeMux I__2926 (
            .O(N__13686),
            .I(N__13680));
    CascadeBuf I__2925 (
            .O(N__13683),
            .I(N__13677));
    CascadeBuf I__2924 (
            .O(N__13680),
            .I(N__13674));
    CascadeMux I__2923 (
            .O(N__13677),
            .I(N__13671));
    CascadeMux I__2922 (
            .O(N__13674),
            .I(N__13668));
    CascadeBuf I__2921 (
            .O(N__13671),
            .I(N__13665));
    CascadeBuf I__2920 (
            .O(N__13668),
            .I(N__13662));
    CascadeMux I__2919 (
            .O(N__13665),
            .I(N__13659));
    CascadeMux I__2918 (
            .O(N__13662),
            .I(N__13656));
    CascadeBuf I__2917 (
            .O(N__13659),
            .I(N__13653));
    CascadeBuf I__2916 (
            .O(N__13656),
            .I(N__13650));
    CascadeMux I__2915 (
            .O(N__13653),
            .I(N__13647));
    CascadeMux I__2914 (
            .O(N__13650),
            .I(N__13644));
    CascadeBuf I__2913 (
            .O(N__13647),
            .I(N__13641));
    CascadeBuf I__2912 (
            .O(N__13644),
            .I(N__13638));
    CascadeMux I__2911 (
            .O(N__13641),
            .I(N__13635));
    CascadeMux I__2910 (
            .O(N__13638),
            .I(N__13632));
    CascadeBuf I__2909 (
            .O(N__13635),
            .I(N__13629));
    CascadeBuf I__2908 (
            .O(N__13632),
            .I(N__13626));
    CascadeMux I__2907 (
            .O(N__13629),
            .I(N__13623));
    CascadeMux I__2906 (
            .O(N__13626),
            .I(N__13620));
    CascadeBuf I__2905 (
            .O(N__13623),
            .I(N__13617));
    CascadeBuf I__2904 (
            .O(N__13620),
            .I(N__13614));
    CascadeMux I__2903 (
            .O(N__13617),
            .I(N__13611));
    CascadeMux I__2902 (
            .O(N__13614),
            .I(N__13608));
    CascadeBuf I__2901 (
            .O(N__13611),
            .I(N__13605));
    CascadeBuf I__2900 (
            .O(N__13608),
            .I(N__13602));
    CascadeMux I__2899 (
            .O(N__13605),
            .I(N__13599));
    CascadeMux I__2898 (
            .O(N__13602),
            .I(N__13596));
    CascadeBuf I__2897 (
            .O(N__13599),
            .I(N__13593));
    CascadeBuf I__2896 (
            .O(N__13596),
            .I(N__13590));
    CascadeMux I__2895 (
            .O(N__13593),
            .I(N__13587));
    CascadeMux I__2894 (
            .O(N__13590),
            .I(N__13584));
    CascadeBuf I__2893 (
            .O(N__13587),
            .I(N__13581));
    CascadeBuf I__2892 (
            .O(N__13584),
            .I(N__13578));
    CascadeMux I__2891 (
            .O(N__13581),
            .I(N__13575));
    CascadeMux I__2890 (
            .O(N__13578),
            .I(N__13572));
    CascadeBuf I__2889 (
            .O(N__13575),
            .I(N__13569));
    CascadeBuf I__2888 (
            .O(N__13572),
            .I(N__13566));
    CascadeMux I__2887 (
            .O(N__13569),
            .I(N__13563));
    CascadeMux I__2886 (
            .O(N__13566),
            .I(N__13560));
    InMux I__2885 (
            .O(N__13563),
            .I(N__13557));
    InMux I__2884 (
            .O(N__13560),
            .I(N__13554));
    LocalMux I__2883 (
            .O(N__13557),
            .I(N__13551));
    LocalMux I__2882 (
            .O(N__13554),
            .I(N__13548));
    Span4Mux_h I__2881 (
            .O(N__13551),
            .I(N__13545));
    Sp12to4 I__2880 (
            .O(N__13548),
            .I(N__13541));
    Sp12to4 I__2879 (
            .O(N__13545),
            .I(N__13538));
    CascadeMux I__2878 (
            .O(N__13544),
            .I(N__13535));
    Span12Mux_s5_v I__2877 (
            .O(N__13541),
            .I(N__13531));
    Span12Mux_s5_v I__2876 (
            .O(N__13538),
            .I(N__13528));
    InMux I__2875 (
            .O(N__13535),
            .I(N__13525));
    InMux I__2874 (
            .O(N__13534),
            .I(N__13522));
    Span12Mux_v I__2873 (
            .O(N__13531),
            .I(N__13519));
    Span12Mux_v I__2872 (
            .O(N__13528),
            .I(N__13516));
    LocalMux I__2871 (
            .O(N__13525),
            .I(RX_ADDR_0));
    LocalMux I__2870 (
            .O(N__13522),
            .I(RX_ADDR_0));
    Odrv12 I__2869 (
            .O(N__13519),
            .I(RX_ADDR_0));
    Odrv12 I__2868 (
            .O(N__13516),
            .I(RX_ADDR_0));
    InMux I__2867 (
            .O(N__13507),
            .I(N__13504));
    LocalMux I__2866 (
            .O(N__13504),
            .I(\receive_module.n136 ));
    InMux I__2865 (
            .O(N__13501),
            .I(bfn_18_14_0_));
    InMux I__2864 (
            .O(N__13498),
            .I(\receive_module.n2727 ));
    InMux I__2863 (
            .O(N__13495),
            .I(\receive_module.n2728 ));
    InMux I__2862 (
            .O(N__13492),
            .I(\receive_module.n2729 ));
    InMux I__2861 (
            .O(N__13489),
            .I(\receive_module.n2730 ));
    CascadeMux I__2860 (
            .O(N__13486),
            .I(N__13482));
    CascadeMux I__2859 (
            .O(N__13485),
            .I(N__13479));
    CascadeBuf I__2858 (
            .O(N__13482),
            .I(N__13476));
    CascadeBuf I__2857 (
            .O(N__13479),
            .I(N__13473));
    CascadeMux I__2856 (
            .O(N__13476),
            .I(N__13470));
    CascadeMux I__2855 (
            .O(N__13473),
            .I(N__13467));
    CascadeBuf I__2854 (
            .O(N__13470),
            .I(N__13464));
    CascadeBuf I__2853 (
            .O(N__13467),
            .I(N__13461));
    CascadeMux I__2852 (
            .O(N__13464),
            .I(N__13458));
    CascadeMux I__2851 (
            .O(N__13461),
            .I(N__13455));
    CascadeBuf I__2850 (
            .O(N__13458),
            .I(N__13452));
    CascadeBuf I__2849 (
            .O(N__13455),
            .I(N__13449));
    CascadeMux I__2848 (
            .O(N__13452),
            .I(N__13446));
    CascadeMux I__2847 (
            .O(N__13449),
            .I(N__13443));
    CascadeBuf I__2846 (
            .O(N__13446),
            .I(N__13440));
    CascadeBuf I__2845 (
            .O(N__13443),
            .I(N__13437));
    CascadeMux I__2844 (
            .O(N__13440),
            .I(N__13434));
    CascadeMux I__2843 (
            .O(N__13437),
            .I(N__13431));
    CascadeBuf I__2842 (
            .O(N__13434),
            .I(N__13428));
    CascadeBuf I__2841 (
            .O(N__13431),
            .I(N__13425));
    CascadeMux I__2840 (
            .O(N__13428),
            .I(N__13422));
    CascadeMux I__2839 (
            .O(N__13425),
            .I(N__13419));
    CascadeBuf I__2838 (
            .O(N__13422),
            .I(N__13416));
    CascadeBuf I__2837 (
            .O(N__13419),
            .I(N__13413));
    CascadeMux I__2836 (
            .O(N__13416),
            .I(N__13410));
    CascadeMux I__2835 (
            .O(N__13413),
            .I(N__13407));
    CascadeBuf I__2834 (
            .O(N__13410),
            .I(N__13404));
    CascadeBuf I__2833 (
            .O(N__13407),
            .I(N__13401));
    CascadeMux I__2832 (
            .O(N__13404),
            .I(N__13398));
    CascadeMux I__2831 (
            .O(N__13401),
            .I(N__13395));
    CascadeBuf I__2830 (
            .O(N__13398),
            .I(N__13392));
    CascadeBuf I__2829 (
            .O(N__13395),
            .I(N__13389));
    CascadeMux I__2828 (
            .O(N__13392),
            .I(N__13386));
    CascadeMux I__2827 (
            .O(N__13389),
            .I(N__13383));
    CascadeBuf I__2826 (
            .O(N__13386),
            .I(N__13380));
    CascadeBuf I__2825 (
            .O(N__13383),
            .I(N__13377));
    CascadeMux I__2824 (
            .O(N__13380),
            .I(N__13374));
    CascadeMux I__2823 (
            .O(N__13377),
            .I(N__13371));
    CascadeBuf I__2822 (
            .O(N__13374),
            .I(N__13368));
    CascadeBuf I__2821 (
            .O(N__13371),
            .I(N__13365));
    CascadeMux I__2820 (
            .O(N__13368),
            .I(N__13362));
    CascadeMux I__2819 (
            .O(N__13365),
            .I(N__13359));
    CascadeBuf I__2818 (
            .O(N__13362),
            .I(N__13356));
    CascadeBuf I__2817 (
            .O(N__13359),
            .I(N__13353));
    CascadeMux I__2816 (
            .O(N__13356),
            .I(N__13350));
    CascadeMux I__2815 (
            .O(N__13353),
            .I(N__13347));
    CascadeBuf I__2814 (
            .O(N__13350),
            .I(N__13344));
    CascadeBuf I__2813 (
            .O(N__13347),
            .I(N__13341));
    CascadeMux I__2812 (
            .O(N__13344),
            .I(N__13338));
    CascadeMux I__2811 (
            .O(N__13341),
            .I(N__13335));
    CascadeBuf I__2810 (
            .O(N__13338),
            .I(N__13332));
    CascadeBuf I__2809 (
            .O(N__13335),
            .I(N__13329));
    CascadeMux I__2808 (
            .O(N__13332),
            .I(N__13326));
    CascadeMux I__2807 (
            .O(N__13329),
            .I(N__13323));
    CascadeBuf I__2806 (
            .O(N__13326),
            .I(N__13320));
    CascadeBuf I__2805 (
            .O(N__13323),
            .I(N__13317));
    CascadeMux I__2804 (
            .O(N__13320),
            .I(N__13314));
    CascadeMux I__2803 (
            .O(N__13317),
            .I(N__13311));
    CascadeBuf I__2802 (
            .O(N__13314),
            .I(N__13308));
    CascadeBuf I__2801 (
            .O(N__13311),
            .I(N__13305));
    CascadeMux I__2800 (
            .O(N__13308),
            .I(N__13302));
    CascadeMux I__2799 (
            .O(N__13305),
            .I(N__13299));
    InMux I__2798 (
            .O(N__13302),
            .I(N__13296));
    InMux I__2797 (
            .O(N__13299),
            .I(N__13293));
    LocalMux I__2796 (
            .O(N__13296),
            .I(N__13290));
    LocalMux I__2795 (
            .O(N__13293),
            .I(N__13287));
    Span4Mux_s1_v I__2794 (
            .O(N__13290),
            .I(N__13284));
    Span4Mux_s1_v I__2793 (
            .O(N__13287),
            .I(N__13281));
    Span4Mux_h I__2792 (
            .O(N__13284),
            .I(N__13278));
    Span4Mux_h I__2791 (
            .O(N__13281),
            .I(N__13275));
    Span4Mux_h I__2790 (
            .O(N__13278),
            .I(N__13269));
    Span4Mux_h I__2789 (
            .O(N__13275),
            .I(N__13269));
    CascadeMux I__2788 (
            .O(N__13274),
            .I(N__13266));
    Sp12to4 I__2787 (
            .O(N__13269),
            .I(N__13262));
    InMux I__2786 (
            .O(N__13266),
            .I(N__13259));
    InMux I__2785 (
            .O(N__13265),
            .I(N__13256));
    Span12Mux_s11_v I__2784 (
            .O(N__13262),
            .I(N__13253));
    LocalMux I__2783 (
            .O(N__13259),
            .I(RX_ADDR_5));
    LocalMux I__2782 (
            .O(N__13256),
            .I(RX_ADDR_5));
    Odrv12 I__2781 (
            .O(N__13253),
            .I(RX_ADDR_5));
    InMux I__2780 (
            .O(N__13246),
            .I(N__13243));
    LocalMux I__2779 (
            .O(N__13243),
            .I(\receive_module.n131 ));
    InMux I__2778 (
            .O(N__13240),
            .I(\receive_module.n2731 ));
    InMux I__2777 (
            .O(N__13237),
            .I(\receive_module.n2732 ));
    CascadeMux I__2776 (
            .O(N__13234),
            .I(N__13231));
    CascadeBuf I__2775 (
            .O(N__13231),
            .I(N__13228));
    CascadeMux I__2774 (
            .O(N__13228),
            .I(N__13224));
    CascadeMux I__2773 (
            .O(N__13227),
            .I(N__13221));
    CascadeBuf I__2772 (
            .O(N__13224),
            .I(N__13218));
    CascadeBuf I__2771 (
            .O(N__13221),
            .I(N__13215));
    CascadeMux I__2770 (
            .O(N__13218),
            .I(N__13212));
    CascadeMux I__2769 (
            .O(N__13215),
            .I(N__13209));
    CascadeBuf I__2768 (
            .O(N__13212),
            .I(N__13206));
    CascadeBuf I__2767 (
            .O(N__13209),
            .I(N__13203));
    CascadeMux I__2766 (
            .O(N__13206),
            .I(N__13200));
    CascadeMux I__2765 (
            .O(N__13203),
            .I(N__13197));
    CascadeBuf I__2764 (
            .O(N__13200),
            .I(N__13194));
    CascadeBuf I__2763 (
            .O(N__13197),
            .I(N__13191));
    CascadeMux I__2762 (
            .O(N__13194),
            .I(N__13188));
    CascadeMux I__2761 (
            .O(N__13191),
            .I(N__13185));
    CascadeBuf I__2760 (
            .O(N__13188),
            .I(N__13182));
    CascadeBuf I__2759 (
            .O(N__13185),
            .I(N__13179));
    CascadeMux I__2758 (
            .O(N__13182),
            .I(N__13176));
    CascadeMux I__2757 (
            .O(N__13179),
            .I(N__13173));
    CascadeBuf I__2756 (
            .O(N__13176),
            .I(N__13170));
    CascadeBuf I__2755 (
            .O(N__13173),
            .I(N__13167));
    CascadeMux I__2754 (
            .O(N__13170),
            .I(N__13164));
    CascadeMux I__2753 (
            .O(N__13167),
            .I(N__13161));
    CascadeBuf I__2752 (
            .O(N__13164),
            .I(N__13158));
    CascadeBuf I__2751 (
            .O(N__13161),
            .I(N__13155));
    CascadeMux I__2750 (
            .O(N__13158),
            .I(N__13152));
    CascadeMux I__2749 (
            .O(N__13155),
            .I(N__13149));
    CascadeBuf I__2748 (
            .O(N__13152),
            .I(N__13146));
    CascadeBuf I__2747 (
            .O(N__13149),
            .I(N__13143));
    CascadeMux I__2746 (
            .O(N__13146),
            .I(N__13140));
    CascadeMux I__2745 (
            .O(N__13143),
            .I(N__13137));
    CascadeBuf I__2744 (
            .O(N__13140),
            .I(N__13134));
    CascadeBuf I__2743 (
            .O(N__13137),
            .I(N__13131));
    CascadeMux I__2742 (
            .O(N__13134),
            .I(N__13128));
    CascadeMux I__2741 (
            .O(N__13131),
            .I(N__13125));
    CascadeBuf I__2740 (
            .O(N__13128),
            .I(N__13122));
    CascadeBuf I__2739 (
            .O(N__13125),
            .I(N__13119));
    CascadeMux I__2738 (
            .O(N__13122),
            .I(N__13116));
    CascadeMux I__2737 (
            .O(N__13119),
            .I(N__13113));
    CascadeBuf I__2736 (
            .O(N__13116),
            .I(N__13110));
    CascadeBuf I__2735 (
            .O(N__13113),
            .I(N__13107));
    CascadeMux I__2734 (
            .O(N__13110),
            .I(N__13104));
    CascadeMux I__2733 (
            .O(N__13107),
            .I(N__13101));
    CascadeBuf I__2732 (
            .O(N__13104),
            .I(N__13098));
    CascadeBuf I__2731 (
            .O(N__13101),
            .I(N__13095));
    CascadeMux I__2730 (
            .O(N__13098),
            .I(N__13092));
    CascadeMux I__2729 (
            .O(N__13095),
            .I(N__13089));
    CascadeBuf I__2728 (
            .O(N__13092),
            .I(N__13086));
    CascadeBuf I__2727 (
            .O(N__13089),
            .I(N__13083));
    CascadeMux I__2726 (
            .O(N__13086),
            .I(N__13080));
    CascadeMux I__2725 (
            .O(N__13083),
            .I(N__13077));
    CascadeBuf I__2724 (
            .O(N__13080),
            .I(N__13074));
    CascadeBuf I__2723 (
            .O(N__13077),
            .I(N__13071));
    CascadeMux I__2722 (
            .O(N__13074),
            .I(N__13068));
    CascadeMux I__2721 (
            .O(N__13071),
            .I(N__13065));
    CascadeBuf I__2720 (
            .O(N__13068),
            .I(N__13062));
    CascadeBuf I__2719 (
            .O(N__13065),
            .I(N__13059));
    CascadeMux I__2718 (
            .O(N__13062),
            .I(N__13056));
    CascadeMux I__2717 (
            .O(N__13059),
            .I(N__13053));
    InMux I__2716 (
            .O(N__13056),
            .I(N__13050));
    CascadeBuf I__2715 (
            .O(N__13053),
            .I(N__13047));
    LocalMux I__2714 (
            .O(N__13050),
            .I(N__13044));
    CascadeMux I__2713 (
            .O(N__13047),
            .I(N__13041));
    Span4Mux_s1_v I__2712 (
            .O(N__13044),
            .I(N__13038));
    InMux I__2711 (
            .O(N__13041),
            .I(N__13035));
    Span4Mux_h I__2710 (
            .O(N__13038),
            .I(N__13032));
    LocalMux I__2709 (
            .O(N__13035),
            .I(N__13029));
    Sp12to4 I__2708 (
            .O(N__13032),
            .I(N__13026));
    Sp12to4 I__2707 (
            .O(N__13029),
            .I(N__13023));
    Span12Mux_s5_v I__2706 (
            .O(N__13026),
            .I(N__13018));
    Span12Mux_s5_v I__2705 (
            .O(N__13023),
            .I(N__13015));
    InMux I__2704 (
            .O(N__13022),
            .I(N__13012));
    InMux I__2703 (
            .O(N__13021),
            .I(N__13009));
    Span12Mux_v I__2702 (
            .O(N__13018),
            .I(N__13004));
    Span12Mux_v I__2701 (
            .O(N__13015),
            .I(N__13004));
    LocalMux I__2700 (
            .O(N__13012),
            .I(RX_ADDR_7));
    LocalMux I__2699 (
            .O(N__13009),
            .I(RX_ADDR_7));
    Odrv12 I__2698 (
            .O(N__13004),
            .I(RX_ADDR_7));
    InMux I__2697 (
            .O(N__12997),
            .I(N__12994));
    LocalMux I__2696 (
            .O(N__12994),
            .I(\receive_module.n129 ));
    InMux I__2695 (
            .O(N__12991),
            .I(\receive_module.n2733 ));
    CascadeMux I__2694 (
            .O(N__12988),
            .I(N__12984));
    CascadeMux I__2693 (
            .O(N__12987),
            .I(N__12981));
    CascadeBuf I__2692 (
            .O(N__12984),
            .I(N__12978));
    CascadeBuf I__2691 (
            .O(N__12981),
            .I(N__12975));
    CascadeMux I__2690 (
            .O(N__12978),
            .I(N__12972));
    CascadeMux I__2689 (
            .O(N__12975),
            .I(N__12969));
    CascadeBuf I__2688 (
            .O(N__12972),
            .I(N__12966));
    CascadeBuf I__2687 (
            .O(N__12969),
            .I(N__12963));
    CascadeMux I__2686 (
            .O(N__12966),
            .I(N__12960));
    CascadeMux I__2685 (
            .O(N__12963),
            .I(N__12957));
    CascadeBuf I__2684 (
            .O(N__12960),
            .I(N__12954));
    CascadeBuf I__2683 (
            .O(N__12957),
            .I(N__12951));
    CascadeMux I__2682 (
            .O(N__12954),
            .I(N__12948));
    CascadeMux I__2681 (
            .O(N__12951),
            .I(N__12945));
    CascadeBuf I__2680 (
            .O(N__12948),
            .I(N__12942));
    CascadeBuf I__2679 (
            .O(N__12945),
            .I(N__12939));
    CascadeMux I__2678 (
            .O(N__12942),
            .I(N__12936));
    CascadeMux I__2677 (
            .O(N__12939),
            .I(N__12933));
    CascadeBuf I__2676 (
            .O(N__12936),
            .I(N__12930));
    CascadeBuf I__2675 (
            .O(N__12933),
            .I(N__12927));
    CascadeMux I__2674 (
            .O(N__12930),
            .I(N__12924));
    CascadeMux I__2673 (
            .O(N__12927),
            .I(N__12921));
    CascadeBuf I__2672 (
            .O(N__12924),
            .I(N__12918));
    CascadeBuf I__2671 (
            .O(N__12921),
            .I(N__12915));
    CascadeMux I__2670 (
            .O(N__12918),
            .I(N__12912));
    CascadeMux I__2669 (
            .O(N__12915),
            .I(N__12909));
    CascadeBuf I__2668 (
            .O(N__12912),
            .I(N__12906));
    CascadeBuf I__2667 (
            .O(N__12909),
            .I(N__12903));
    CascadeMux I__2666 (
            .O(N__12906),
            .I(N__12900));
    CascadeMux I__2665 (
            .O(N__12903),
            .I(N__12897));
    CascadeBuf I__2664 (
            .O(N__12900),
            .I(N__12894));
    CascadeBuf I__2663 (
            .O(N__12897),
            .I(N__12891));
    CascadeMux I__2662 (
            .O(N__12894),
            .I(N__12888));
    CascadeMux I__2661 (
            .O(N__12891),
            .I(N__12885));
    CascadeBuf I__2660 (
            .O(N__12888),
            .I(N__12882));
    CascadeBuf I__2659 (
            .O(N__12885),
            .I(N__12879));
    CascadeMux I__2658 (
            .O(N__12882),
            .I(N__12876));
    CascadeMux I__2657 (
            .O(N__12879),
            .I(N__12873));
    CascadeBuf I__2656 (
            .O(N__12876),
            .I(N__12870));
    CascadeBuf I__2655 (
            .O(N__12873),
            .I(N__12867));
    CascadeMux I__2654 (
            .O(N__12870),
            .I(N__12864));
    CascadeMux I__2653 (
            .O(N__12867),
            .I(N__12861));
    CascadeBuf I__2652 (
            .O(N__12864),
            .I(N__12858));
    CascadeBuf I__2651 (
            .O(N__12861),
            .I(N__12855));
    CascadeMux I__2650 (
            .O(N__12858),
            .I(N__12852));
    CascadeMux I__2649 (
            .O(N__12855),
            .I(N__12849));
    CascadeBuf I__2648 (
            .O(N__12852),
            .I(N__12846));
    CascadeBuf I__2647 (
            .O(N__12849),
            .I(N__12843));
    CascadeMux I__2646 (
            .O(N__12846),
            .I(N__12840));
    CascadeMux I__2645 (
            .O(N__12843),
            .I(N__12837));
    CascadeBuf I__2644 (
            .O(N__12840),
            .I(N__12834));
    CascadeBuf I__2643 (
            .O(N__12837),
            .I(N__12831));
    CascadeMux I__2642 (
            .O(N__12834),
            .I(N__12828));
    CascadeMux I__2641 (
            .O(N__12831),
            .I(N__12825));
    CascadeBuf I__2640 (
            .O(N__12828),
            .I(N__12822));
    CascadeBuf I__2639 (
            .O(N__12825),
            .I(N__12819));
    CascadeMux I__2638 (
            .O(N__12822),
            .I(N__12816));
    CascadeMux I__2637 (
            .O(N__12819),
            .I(N__12813));
    CascadeBuf I__2636 (
            .O(N__12816),
            .I(N__12810));
    CascadeBuf I__2635 (
            .O(N__12813),
            .I(N__12807));
    CascadeMux I__2634 (
            .O(N__12810),
            .I(N__12804));
    CascadeMux I__2633 (
            .O(N__12807),
            .I(N__12801));
    InMux I__2632 (
            .O(N__12804),
            .I(N__12798));
    InMux I__2631 (
            .O(N__12801),
            .I(N__12795));
    LocalMux I__2630 (
            .O(N__12798),
            .I(N__12792));
    LocalMux I__2629 (
            .O(N__12795),
            .I(N__12789));
    Span4Mux_h I__2628 (
            .O(N__12792),
            .I(N__12786));
    Span4Mux_h I__2627 (
            .O(N__12789),
            .I(N__12783));
    Sp12to4 I__2626 (
            .O(N__12786),
            .I(N__12780));
    Sp12to4 I__2625 (
            .O(N__12783),
            .I(N__12777));
    Span12Mux_s5_v I__2624 (
            .O(N__12780),
            .I(N__12772));
    Span12Mux_s5_v I__2623 (
            .O(N__12777),
            .I(N__12769));
    InMux I__2622 (
            .O(N__12776),
            .I(N__12766));
    InMux I__2621 (
            .O(N__12775),
            .I(N__12763));
    Span12Mux_v I__2620 (
            .O(N__12772),
            .I(N__12758));
    Span12Mux_v I__2619 (
            .O(N__12769),
            .I(N__12758));
    LocalMux I__2618 (
            .O(N__12766),
            .I(RX_ADDR_8));
    LocalMux I__2617 (
            .O(N__12763),
            .I(RX_ADDR_8));
    Odrv12 I__2616 (
            .O(N__12758),
            .I(RX_ADDR_8));
    InMux I__2615 (
            .O(N__12751),
            .I(N__12748));
    LocalMux I__2614 (
            .O(N__12748),
            .I(\receive_module.n128 ));
    InMux I__2613 (
            .O(N__12745),
            .I(bfn_18_15_0_));
    InMux I__2612 (
            .O(N__12742),
            .I(N__12739));
    LocalMux I__2611 (
            .O(N__12739),
            .I(N__12736));
    Span4Mux_v I__2610 (
            .O(N__12736),
            .I(N__12733));
    Sp12to4 I__2609 (
            .O(N__12733),
            .I(N__12730));
    Odrv12 I__2608 (
            .O(N__12730),
            .I(\line_buffer.n726 ));
    InMux I__2607 (
            .O(N__12727),
            .I(N__12724));
    LocalMux I__2606 (
            .O(N__12724),
            .I(N__12721));
    Span12Mux_v I__2605 (
            .O(N__12721),
            .I(N__12718));
    Span12Mux_v I__2604 (
            .O(N__12718),
            .I(N__12715));
    Odrv12 I__2603 (
            .O(N__12715),
            .I(\line_buffer.n718 ));
    InMux I__2602 (
            .O(N__12712),
            .I(N__12709));
    LocalMux I__2601 (
            .O(N__12709),
            .I(N__12706));
    Span12Mux_v I__2600 (
            .O(N__12706),
            .I(N__12703));
    Odrv12 I__2599 (
            .O(N__12703),
            .I(\line_buffer.n629 ));
    InMux I__2598 (
            .O(N__12700),
            .I(N__12697));
    LocalMux I__2597 (
            .O(N__12697),
            .I(N__12694));
    Span4Mux_v I__2596 (
            .O(N__12694),
            .I(N__12691));
    Span4Mux_h I__2595 (
            .O(N__12691),
            .I(N__12688));
    Span4Mux_h I__2594 (
            .O(N__12688),
            .I(N__12685));
    Odrv4 I__2593 (
            .O(N__12685),
            .I(\line_buffer.n621 ));
    CascadeMux I__2592 (
            .O(N__12682),
            .I(\line_buffer.n3161_cascade_ ));
    InMux I__2591 (
            .O(N__12679),
            .I(N__12676));
    LocalMux I__2590 (
            .O(N__12676),
            .I(\line_buffer.n3164 ));
    InMux I__2589 (
            .O(N__12673),
            .I(N__12670));
    LocalMux I__2588 (
            .O(N__12670),
            .I(N__12667));
    Span4Mux_h I__2587 (
            .O(N__12667),
            .I(N__12664));
    Span4Mux_h I__2586 (
            .O(N__12664),
            .I(N__12661));
    Odrv4 I__2585 (
            .O(N__12661),
            .I(\line_buffer.n630 ));
    InMux I__2584 (
            .O(N__12658),
            .I(N__12655));
    LocalMux I__2583 (
            .O(N__12655),
            .I(N__12652));
    Span4Mux_h I__2582 (
            .O(N__12652),
            .I(N__12649));
    Span4Mux_h I__2581 (
            .O(N__12649),
            .I(N__12646));
    Span4Mux_h I__2580 (
            .O(N__12646),
            .I(N__12643));
    Odrv4 I__2579 (
            .O(N__12643),
            .I(\line_buffer.n622 ));
    InMux I__2578 (
            .O(N__12640),
            .I(N__12637));
    LocalMux I__2577 (
            .O(N__12637),
            .I(N__12634));
    Odrv4 I__2576 (
            .O(N__12634),
            .I(\line_buffer.n3042 ));
    SRMux I__2575 (
            .O(N__12631),
            .I(N__12628));
    LocalMux I__2574 (
            .O(N__12628),
            .I(N__12623));
    SRMux I__2573 (
            .O(N__12627),
            .I(N__12620));
    SRMux I__2572 (
            .O(N__12626),
            .I(N__12617));
    Span4Mux_s2_v I__2571 (
            .O(N__12623),
            .I(N__12607));
    LocalMux I__2570 (
            .O(N__12620),
            .I(N__12607));
    LocalMux I__2569 (
            .O(N__12617),
            .I(N__12607));
    SRMux I__2568 (
            .O(N__12616),
            .I(N__12604));
    SRMux I__2567 (
            .O(N__12615),
            .I(N__12601));
    SRMux I__2566 (
            .O(N__12614),
            .I(N__12596));
    Span4Mux_v I__2565 (
            .O(N__12607),
            .I(N__12587));
    LocalMux I__2564 (
            .O(N__12604),
            .I(N__12587));
    LocalMux I__2563 (
            .O(N__12601),
            .I(N__12587));
    SRMux I__2562 (
            .O(N__12600),
            .I(N__12584));
    SRMux I__2561 (
            .O(N__12599),
            .I(N__12581));
    LocalMux I__2560 (
            .O(N__12596),
            .I(N__12576));
    SRMux I__2559 (
            .O(N__12595),
            .I(N__12573));
    SRMux I__2558 (
            .O(N__12594),
            .I(N__12570));
    Span4Mux_v I__2557 (
            .O(N__12587),
            .I(N__12561));
    LocalMux I__2556 (
            .O(N__12584),
            .I(N__12561));
    LocalMux I__2555 (
            .O(N__12581),
            .I(N__12561));
    SRMux I__2554 (
            .O(N__12580),
            .I(N__12558));
    SRMux I__2553 (
            .O(N__12579),
            .I(N__12555));
    Span4Mux_s2_v I__2552 (
            .O(N__12576),
            .I(N__12546));
    LocalMux I__2551 (
            .O(N__12573),
            .I(N__12546));
    LocalMux I__2550 (
            .O(N__12570),
            .I(N__12546));
    SRMux I__2549 (
            .O(N__12569),
            .I(N__12543));
    SRMux I__2548 (
            .O(N__12568),
            .I(N__12540));
    Span4Mux_v I__2547 (
            .O(N__12561),
            .I(N__12529));
    LocalMux I__2546 (
            .O(N__12558),
            .I(N__12529));
    LocalMux I__2545 (
            .O(N__12555),
            .I(N__12529));
    SRMux I__2544 (
            .O(N__12554),
            .I(N__12526));
    SRMux I__2543 (
            .O(N__12553),
            .I(N__12523));
    Span4Mux_v I__2542 (
            .O(N__12546),
            .I(N__12514));
    LocalMux I__2541 (
            .O(N__12543),
            .I(N__12514));
    LocalMux I__2540 (
            .O(N__12540),
            .I(N__12514));
    SRMux I__2539 (
            .O(N__12539),
            .I(N__12511));
    SRMux I__2538 (
            .O(N__12538),
            .I(N__12508));
    IoInMux I__2537 (
            .O(N__12537),
            .I(N__12503));
    IoInMux I__2536 (
            .O(N__12536),
            .I(N__12500));
    Span4Mux_v I__2535 (
            .O(N__12529),
            .I(N__12493));
    LocalMux I__2534 (
            .O(N__12526),
            .I(N__12493));
    LocalMux I__2533 (
            .O(N__12523),
            .I(N__12493));
    SRMux I__2532 (
            .O(N__12522),
            .I(N__12490));
    SRMux I__2531 (
            .O(N__12521),
            .I(N__12487));
    Span4Mux_v I__2530 (
            .O(N__12514),
            .I(N__12478));
    LocalMux I__2529 (
            .O(N__12511),
            .I(N__12478));
    LocalMux I__2528 (
            .O(N__12508),
            .I(N__12478));
    SRMux I__2527 (
            .O(N__12507),
            .I(N__12475));
    SRMux I__2526 (
            .O(N__12506),
            .I(N__12472));
    LocalMux I__2525 (
            .O(N__12503),
            .I(N__12465));
    LocalMux I__2524 (
            .O(N__12500),
            .I(N__12465));
    Span4Mux_v I__2523 (
            .O(N__12493),
            .I(N__12458));
    LocalMux I__2522 (
            .O(N__12490),
            .I(N__12458));
    LocalMux I__2521 (
            .O(N__12487),
            .I(N__12458));
    SRMux I__2520 (
            .O(N__12486),
            .I(N__12455));
    SRMux I__2519 (
            .O(N__12485),
            .I(N__12452));
    Span4Mux_v I__2518 (
            .O(N__12478),
            .I(N__12444));
    LocalMux I__2517 (
            .O(N__12475),
            .I(N__12444));
    LocalMux I__2516 (
            .O(N__12472),
            .I(N__12444));
    SRMux I__2515 (
            .O(N__12471),
            .I(N__12441));
    SRMux I__2514 (
            .O(N__12470),
            .I(N__12438));
    IoSpan4Mux I__2513 (
            .O(N__12465),
            .I(N__12433));
    Span4Mux_v I__2512 (
            .O(N__12458),
            .I(N__12426));
    LocalMux I__2511 (
            .O(N__12455),
            .I(N__12426));
    LocalMux I__2510 (
            .O(N__12452),
            .I(N__12426));
    SRMux I__2509 (
            .O(N__12451),
            .I(N__12423));
    Span4Mux_v I__2508 (
            .O(N__12444),
            .I(N__12416));
    LocalMux I__2507 (
            .O(N__12441),
            .I(N__12416));
    LocalMux I__2506 (
            .O(N__12438),
            .I(N__12416));
    SRMux I__2505 (
            .O(N__12437),
            .I(N__12413));
    SRMux I__2504 (
            .O(N__12436),
            .I(N__12410));
    Span4Mux_s0_v I__2503 (
            .O(N__12433),
            .I(N__12404));
    Span4Mux_v I__2502 (
            .O(N__12426),
            .I(N__12399));
    LocalMux I__2501 (
            .O(N__12423),
            .I(N__12399));
    Span4Mux_v I__2500 (
            .O(N__12416),
            .I(N__12392));
    LocalMux I__2499 (
            .O(N__12413),
            .I(N__12392));
    LocalMux I__2498 (
            .O(N__12410),
            .I(N__12392));
    SRMux I__2497 (
            .O(N__12409),
            .I(N__12389));
    SRMux I__2496 (
            .O(N__12408),
            .I(N__12386));
    SRMux I__2495 (
            .O(N__12407),
            .I(N__12383));
    Sp12to4 I__2494 (
            .O(N__12404),
            .I(N__12380));
    Span4Mux_s1_v I__2493 (
            .O(N__12399),
            .I(N__12377));
    Span4Mux_v I__2492 (
            .O(N__12392),
            .I(N__12370));
    LocalMux I__2491 (
            .O(N__12389),
            .I(N__12370));
    LocalMux I__2490 (
            .O(N__12386),
            .I(N__12370));
    LocalMux I__2489 (
            .O(N__12383),
            .I(N__12367));
    Span12Mux_s11_v I__2488 (
            .O(N__12380),
            .I(N__12364));
    Span4Mux_h I__2487 (
            .O(N__12377),
            .I(N__12361));
    Span4Mux_v I__2486 (
            .O(N__12370),
            .I(N__12356));
    Span4Mux_s1_v I__2485 (
            .O(N__12367),
            .I(N__12356));
    Span12Mux_v I__2484 (
            .O(N__12364),
            .I(N__12353));
    Span4Mux_h I__2483 (
            .O(N__12361),
            .I(N__12348));
    Span4Mux_h I__2482 (
            .O(N__12356),
            .I(N__12348));
    Odrv12 I__2481 (
            .O(N__12353),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2480 (
            .O(N__12348),
            .I(CONSTANT_ONE_NET));
    InMux I__2479 (
            .O(N__12343),
            .I(N__12340));
    LocalMux I__2478 (
            .O(N__12340),
            .I(N__12337));
    Span4Mux_v I__2477 (
            .O(N__12337),
            .I(N__12334));
    Sp12to4 I__2476 (
            .O(N__12334),
            .I(N__12331));
    Span12Mux_h I__2475 (
            .O(N__12331),
            .I(N__12328));
    Odrv12 I__2474 (
            .O(N__12328),
            .I(\line_buffer.n623 ));
    CascadeMux I__2473 (
            .O(N__12325),
            .I(N__12322));
    InMux I__2472 (
            .O(N__12322),
            .I(N__12319));
    LocalMux I__2471 (
            .O(N__12319),
            .I(N__12316));
    Span4Mux_h I__2470 (
            .O(N__12316),
            .I(N__12313));
    Span4Mux_h I__2469 (
            .O(N__12313),
            .I(N__12310));
    Span4Mux_v I__2468 (
            .O(N__12310),
            .I(N__12307));
    Odrv4 I__2467 (
            .O(N__12307),
            .I(\line_buffer.n615 ));
    InMux I__2466 (
            .O(N__12304),
            .I(N__12301));
    LocalMux I__2465 (
            .O(N__12301),
            .I(N__12298));
    Span4Mux_v I__2464 (
            .O(N__12298),
            .I(N__12295));
    Sp12to4 I__2463 (
            .O(N__12295),
            .I(N__12292));
    Odrv12 I__2462 (
            .O(N__12292),
            .I(\line_buffer.n720 ));
    InMux I__2461 (
            .O(N__12289),
            .I(N__12286));
    LocalMux I__2460 (
            .O(N__12286),
            .I(N__12283));
    Span4Mux_h I__2459 (
            .O(N__12283),
            .I(N__12280));
    Span4Mux_v I__2458 (
            .O(N__12280),
            .I(N__12277));
    Span4Mux_h I__2457 (
            .O(N__12277),
            .I(N__12274));
    Odrv4 I__2456 (
            .O(N__12274),
            .I(\line_buffer.n712 ));
    InMux I__2455 (
            .O(N__12271),
            .I(N__12268));
    LocalMux I__2454 (
            .O(N__12268),
            .I(\line_buffer.n3113 ));
    InMux I__2453 (
            .O(N__12265),
            .I(N__12262));
    LocalMux I__2452 (
            .O(N__12262),
            .I(N__12259));
    Span4Mux_v I__2451 (
            .O(N__12259),
            .I(N__12256));
    Span4Mux_v I__2450 (
            .O(N__12256),
            .I(N__12253));
    Sp12to4 I__2449 (
            .O(N__12253),
            .I(N__12250));
    Odrv12 I__2448 (
            .O(N__12250),
            .I(\line_buffer.n688 ));
    CascadeMux I__2447 (
            .O(N__12247),
            .I(N__12244));
    InMux I__2446 (
            .O(N__12244),
            .I(N__12241));
    LocalMux I__2445 (
            .O(N__12241),
            .I(N__12238));
    Span4Mux_v I__2444 (
            .O(N__12238),
            .I(N__12235));
    Span4Mux_h I__2443 (
            .O(N__12235),
            .I(N__12232));
    Odrv4 I__2442 (
            .O(N__12232),
            .I(\line_buffer.n680 ));
    CascadeMux I__2441 (
            .O(N__12229),
            .I(\line_buffer.n3122_cascade_ ));
    InMux I__2440 (
            .O(N__12226),
            .I(N__12223));
    LocalMux I__2439 (
            .O(N__12223),
            .I(\line_buffer.n3116 ));
    InMux I__2438 (
            .O(N__12220),
            .I(N__12217));
    LocalMux I__2437 (
            .O(N__12217),
            .I(N__12214));
    Span4Mux_h I__2436 (
            .O(N__12214),
            .I(N__12211));
    Odrv4 I__2435 (
            .O(N__12211),
            .I(TX_DATA_0));
    InMux I__2434 (
            .O(N__12208),
            .I(N__12205));
    LocalMux I__2433 (
            .O(N__12205),
            .I(N__12202));
    Span12Mux_v I__2432 (
            .O(N__12202),
            .I(N__12199));
    Span12Mux_v I__2431 (
            .O(N__12199),
            .I(N__12196));
    Odrv12 I__2430 (
            .O(N__12196),
            .I(\line_buffer.n745 ));
    CascadeMux I__2429 (
            .O(N__12193),
            .I(N__12190));
    InMux I__2428 (
            .O(N__12190),
            .I(N__12187));
    LocalMux I__2427 (
            .O(N__12187),
            .I(N__12184));
    Span4Mux_h I__2426 (
            .O(N__12184),
            .I(N__12181));
    Span4Mux_h I__2425 (
            .O(N__12181),
            .I(N__12178));
    Span4Mux_h I__2424 (
            .O(N__12178),
            .I(N__12175));
    Odrv4 I__2423 (
            .O(N__12175),
            .I(\line_buffer.n753 ));
    InMux I__2422 (
            .O(N__12172),
            .I(N__12169));
    LocalMux I__2421 (
            .O(N__12169),
            .I(\line_buffer.n3137 ));
    SRMux I__2420 (
            .O(N__12166),
            .I(N__12162));
    SRMux I__2419 (
            .O(N__12165),
            .I(N__12157));
    LocalMux I__2418 (
            .O(N__12162),
            .I(N__12154));
    SRMux I__2417 (
            .O(N__12161),
            .I(N__12151));
    SRMux I__2416 (
            .O(N__12160),
            .I(N__12148));
    LocalMux I__2415 (
            .O(N__12157),
            .I(N__12145));
    Span4Mux_s1_v I__2414 (
            .O(N__12154),
            .I(N__12138));
    LocalMux I__2413 (
            .O(N__12151),
            .I(N__12138));
    LocalMux I__2412 (
            .O(N__12148),
            .I(N__12138));
    Span4Mux_h I__2411 (
            .O(N__12145),
            .I(N__12135));
    Sp12to4 I__2410 (
            .O(N__12138),
            .I(N__12132));
    Span4Mux_h I__2409 (
            .O(N__12135),
            .I(N__12129));
    Span12Mux_v I__2408 (
            .O(N__12132),
            .I(N__12126));
    Span4Mux_h I__2407 (
            .O(N__12129),
            .I(N__12123));
    Odrv12 I__2406 (
            .O(N__12126),
            .I(\line_buffer.n761 ));
    Odrv4 I__2405 (
            .O(N__12123),
            .I(\line_buffer.n761 ));
    InMux I__2404 (
            .O(N__12118),
            .I(N__12115));
    LocalMux I__2403 (
            .O(N__12115),
            .I(N__12111));
    InMux I__2402 (
            .O(N__12114),
            .I(N__12108));
    Span4Mux_h I__2401 (
            .O(N__12111),
            .I(N__12105));
    LocalMux I__2400 (
            .O(N__12108),
            .I(\transmit_module.n387 ));
    Odrv4 I__2399 (
            .O(N__12105),
            .I(\transmit_module.n387 ));
    IoInMux I__2398 (
            .O(N__12100),
            .I(N__12097));
    LocalMux I__2397 (
            .O(N__12097),
            .I(N__12094));
    Span12Mux_s10_h I__2396 (
            .O(N__12094),
            .I(N__12090));
    InMux I__2395 (
            .O(N__12093),
            .I(N__12087));
    Span12Mux_v I__2394 (
            .O(N__12090),
            .I(N__12082));
    LocalMux I__2393 (
            .O(N__12087),
            .I(N__12079));
    InMux I__2392 (
            .O(N__12086),
            .I(N__12076));
    InMux I__2391 (
            .O(N__12085),
            .I(N__12073));
    Odrv12 I__2390 (
            .O(N__12082),
            .I(DEBUG_c_1));
    Odrv4 I__2389 (
            .O(N__12079),
            .I(DEBUG_c_1));
    LocalMux I__2388 (
            .O(N__12076),
            .I(DEBUG_c_1));
    LocalMux I__2387 (
            .O(N__12073),
            .I(DEBUG_c_1));
    CascadeMux I__2386 (
            .O(N__12064),
            .I(N__12060));
    CascadeMux I__2385 (
            .O(N__12063),
            .I(N__12057));
    CascadeBuf I__2384 (
            .O(N__12060),
            .I(N__12054));
    CascadeBuf I__2383 (
            .O(N__12057),
            .I(N__12051));
    CascadeMux I__2382 (
            .O(N__12054),
            .I(N__12048));
    CascadeMux I__2381 (
            .O(N__12051),
            .I(N__12045));
    CascadeBuf I__2380 (
            .O(N__12048),
            .I(N__12042));
    CascadeBuf I__2379 (
            .O(N__12045),
            .I(N__12039));
    CascadeMux I__2378 (
            .O(N__12042),
            .I(N__12036));
    CascadeMux I__2377 (
            .O(N__12039),
            .I(N__12033));
    CascadeBuf I__2376 (
            .O(N__12036),
            .I(N__12030));
    CascadeBuf I__2375 (
            .O(N__12033),
            .I(N__12027));
    CascadeMux I__2374 (
            .O(N__12030),
            .I(N__12024));
    CascadeMux I__2373 (
            .O(N__12027),
            .I(N__12021));
    CascadeBuf I__2372 (
            .O(N__12024),
            .I(N__12018));
    CascadeBuf I__2371 (
            .O(N__12021),
            .I(N__12015));
    CascadeMux I__2370 (
            .O(N__12018),
            .I(N__12012));
    CascadeMux I__2369 (
            .O(N__12015),
            .I(N__12009));
    CascadeBuf I__2368 (
            .O(N__12012),
            .I(N__12006));
    CascadeBuf I__2367 (
            .O(N__12009),
            .I(N__12003));
    CascadeMux I__2366 (
            .O(N__12006),
            .I(N__12000));
    CascadeMux I__2365 (
            .O(N__12003),
            .I(N__11997));
    CascadeBuf I__2364 (
            .O(N__12000),
            .I(N__11994));
    CascadeBuf I__2363 (
            .O(N__11997),
            .I(N__11991));
    CascadeMux I__2362 (
            .O(N__11994),
            .I(N__11988));
    CascadeMux I__2361 (
            .O(N__11991),
            .I(N__11985));
    CascadeBuf I__2360 (
            .O(N__11988),
            .I(N__11982));
    CascadeBuf I__2359 (
            .O(N__11985),
            .I(N__11979));
    CascadeMux I__2358 (
            .O(N__11982),
            .I(N__11976));
    CascadeMux I__2357 (
            .O(N__11979),
            .I(N__11973));
    CascadeBuf I__2356 (
            .O(N__11976),
            .I(N__11970));
    CascadeBuf I__2355 (
            .O(N__11973),
            .I(N__11967));
    CascadeMux I__2354 (
            .O(N__11970),
            .I(N__11964));
    CascadeMux I__2353 (
            .O(N__11967),
            .I(N__11961));
    CascadeBuf I__2352 (
            .O(N__11964),
            .I(N__11958));
    CascadeBuf I__2351 (
            .O(N__11961),
            .I(N__11955));
    CascadeMux I__2350 (
            .O(N__11958),
            .I(N__11952));
    CascadeMux I__2349 (
            .O(N__11955),
            .I(N__11949));
    CascadeBuf I__2348 (
            .O(N__11952),
            .I(N__11946));
    CascadeBuf I__2347 (
            .O(N__11949),
            .I(N__11943));
    CascadeMux I__2346 (
            .O(N__11946),
            .I(N__11940));
    CascadeMux I__2345 (
            .O(N__11943),
            .I(N__11937));
    CascadeBuf I__2344 (
            .O(N__11940),
            .I(N__11934));
    CascadeBuf I__2343 (
            .O(N__11937),
            .I(N__11931));
    CascadeMux I__2342 (
            .O(N__11934),
            .I(N__11928));
    CascadeMux I__2341 (
            .O(N__11931),
            .I(N__11925));
    CascadeBuf I__2340 (
            .O(N__11928),
            .I(N__11922));
    CascadeBuf I__2339 (
            .O(N__11925),
            .I(N__11919));
    CascadeMux I__2338 (
            .O(N__11922),
            .I(N__11916));
    CascadeMux I__2337 (
            .O(N__11919),
            .I(N__11913));
    CascadeBuf I__2336 (
            .O(N__11916),
            .I(N__11910));
    CascadeBuf I__2335 (
            .O(N__11913),
            .I(N__11907));
    CascadeMux I__2334 (
            .O(N__11910),
            .I(N__11904));
    CascadeMux I__2333 (
            .O(N__11907),
            .I(N__11901));
    CascadeBuf I__2332 (
            .O(N__11904),
            .I(N__11898));
    CascadeBuf I__2331 (
            .O(N__11901),
            .I(N__11895));
    CascadeMux I__2330 (
            .O(N__11898),
            .I(N__11892));
    CascadeMux I__2329 (
            .O(N__11895),
            .I(N__11889));
    CascadeBuf I__2328 (
            .O(N__11892),
            .I(N__11886));
    CascadeBuf I__2327 (
            .O(N__11889),
            .I(N__11883));
    CascadeMux I__2326 (
            .O(N__11886),
            .I(N__11880));
    CascadeMux I__2325 (
            .O(N__11883),
            .I(N__11877));
    InMux I__2324 (
            .O(N__11880),
            .I(N__11874));
    InMux I__2323 (
            .O(N__11877),
            .I(N__11871));
    LocalMux I__2322 (
            .O(N__11874),
            .I(N__11868));
    LocalMux I__2321 (
            .O(N__11871),
            .I(N__11865));
    Span12Mux_s11_h I__2320 (
            .O(N__11868),
            .I(N__11862));
    Span12Mux_s8_h I__2319 (
            .O(N__11865),
            .I(N__11859));
    Span12Mux_v I__2318 (
            .O(N__11862),
            .I(N__11854));
    Span12Mux_v I__2317 (
            .O(N__11859),
            .I(N__11854));
    Odrv12 I__2316 (
            .O(N__11854),
            .I(n27));
    IoInMux I__2315 (
            .O(N__11851),
            .I(N__11848));
    LocalMux I__2314 (
            .O(N__11848),
            .I(N__11845));
    Span4Mux_s3_h I__2313 (
            .O(N__11845),
            .I(N__11842));
    Span4Mux_h I__2312 (
            .O(N__11842),
            .I(N__11839));
    Span4Mux_h I__2311 (
            .O(N__11839),
            .I(N__11836));
    Span4Mux_h I__2310 (
            .O(N__11836),
            .I(N__11830));
    InMux I__2309 (
            .O(N__11835),
            .I(N__11827));
    InMux I__2308 (
            .O(N__11834),
            .I(N__11824));
    InMux I__2307 (
            .O(N__11833),
            .I(N__11821));
    Odrv4 I__2306 (
            .O(N__11830),
            .I(DEBUG_c_7));
    LocalMux I__2305 (
            .O(N__11827),
            .I(DEBUG_c_7));
    LocalMux I__2304 (
            .O(N__11824),
            .I(DEBUG_c_7));
    LocalMux I__2303 (
            .O(N__11821),
            .I(DEBUG_c_7));
    InMux I__2302 (
            .O(N__11812),
            .I(N__11808));
    CascadeMux I__2301 (
            .O(N__11811),
            .I(N__11805));
    LocalMux I__2300 (
            .O(N__11808),
            .I(N__11802));
    InMux I__2299 (
            .O(N__11805),
            .I(N__11799));
    Span4Mux_h I__2298 (
            .O(N__11802),
            .I(N__11796));
    LocalMux I__2297 (
            .O(N__11799),
            .I(\transmit_module.n381 ));
    Odrv4 I__2296 (
            .O(N__11796),
            .I(\transmit_module.n381 ));
    CascadeMux I__2295 (
            .O(N__11791),
            .I(N__11788));
    CascadeBuf I__2294 (
            .O(N__11788),
            .I(N__11785));
    CascadeMux I__2293 (
            .O(N__11785),
            .I(N__11781));
    CascadeMux I__2292 (
            .O(N__11784),
            .I(N__11778));
    CascadeBuf I__2291 (
            .O(N__11781),
            .I(N__11775));
    CascadeBuf I__2290 (
            .O(N__11778),
            .I(N__11772));
    CascadeMux I__2289 (
            .O(N__11775),
            .I(N__11769));
    CascadeMux I__2288 (
            .O(N__11772),
            .I(N__11766));
    CascadeBuf I__2287 (
            .O(N__11769),
            .I(N__11763));
    CascadeBuf I__2286 (
            .O(N__11766),
            .I(N__11760));
    CascadeMux I__2285 (
            .O(N__11763),
            .I(N__11757));
    CascadeMux I__2284 (
            .O(N__11760),
            .I(N__11754));
    CascadeBuf I__2283 (
            .O(N__11757),
            .I(N__11751));
    CascadeBuf I__2282 (
            .O(N__11754),
            .I(N__11748));
    CascadeMux I__2281 (
            .O(N__11751),
            .I(N__11745));
    CascadeMux I__2280 (
            .O(N__11748),
            .I(N__11742));
    CascadeBuf I__2279 (
            .O(N__11745),
            .I(N__11739));
    CascadeBuf I__2278 (
            .O(N__11742),
            .I(N__11736));
    CascadeMux I__2277 (
            .O(N__11739),
            .I(N__11733));
    CascadeMux I__2276 (
            .O(N__11736),
            .I(N__11730));
    CascadeBuf I__2275 (
            .O(N__11733),
            .I(N__11727));
    CascadeBuf I__2274 (
            .O(N__11730),
            .I(N__11724));
    CascadeMux I__2273 (
            .O(N__11727),
            .I(N__11721));
    CascadeMux I__2272 (
            .O(N__11724),
            .I(N__11718));
    CascadeBuf I__2271 (
            .O(N__11721),
            .I(N__11715));
    CascadeBuf I__2270 (
            .O(N__11718),
            .I(N__11712));
    CascadeMux I__2269 (
            .O(N__11715),
            .I(N__11709));
    CascadeMux I__2268 (
            .O(N__11712),
            .I(N__11706));
    CascadeBuf I__2267 (
            .O(N__11709),
            .I(N__11703));
    CascadeBuf I__2266 (
            .O(N__11706),
            .I(N__11700));
    CascadeMux I__2265 (
            .O(N__11703),
            .I(N__11697));
    CascadeMux I__2264 (
            .O(N__11700),
            .I(N__11694));
    CascadeBuf I__2263 (
            .O(N__11697),
            .I(N__11691));
    CascadeBuf I__2262 (
            .O(N__11694),
            .I(N__11688));
    CascadeMux I__2261 (
            .O(N__11691),
            .I(N__11685));
    CascadeMux I__2260 (
            .O(N__11688),
            .I(N__11682));
    CascadeBuf I__2259 (
            .O(N__11685),
            .I(N__11679));
    CascadeBuf I__2258 (
            .O(N__11682),
            .I(N__11676));
    CascadeMux I__2257 (
            .O(N__11679),
            .I(N__11673));
    CascadeMux I__2256 (
            .O(N__11676),
            .I(N__11670));
    CascadeBuf I__2255 (
            .O(N__11673),
            .I(N__11667));
    CascadeBuf I__2254 (
            .O(N__11670),
            .I(N__11664));
    CascadeMux I__2253 (
            .O(N__11667),
            .I(N__11661));
    CascadeMux I__2252 (
            .O(N__11664),
            .I(N__11658));
    CascadeBuf I__2251 (
            .O(N__11661),
            .I(N__11655));
    CascadeBuf I__2250 (
            .O(N__11658),
            .I(N__11652));
    CascadeMux I__2249 (
            .O(N__11655),
            .I(N__11649));
    CascadeMux I__2248 (
            .O(N__11652),
            .I(N__11646));
    CascadeBuf I__2247 (
            .O(N__11649),
            .I(N__11643));
    CascadeBuf I__2246 (
            .O(N__11646),
            .I(N__11640));
    CascadeMux I__2245 (
            .O(N__11643),
            .I(N__11637));
    CascadeMux I__2244 (
            .O(N__11640),
            .I(N__11634));
    CascadeBuf I__2243 (
            .O(N__11637),
            .I(N__11631));
    CascadeBuf I__2242 (
            .O(N__11634),
            .I(N__11628));
    CascadeMux I__2241 (
            .O(N__11631),
            .I(N__11625));
    CascadeMux I__2240 (
            .O(N__11628),
            .I(N__11622));
    CascadeBuf I__2239 (
            .O(N__11625),
            .I(N__11619));
    CascadeBuf I__2238 (
            .O(N__11622),
            .I(N__11616));
    CascadeMux I__2237 (
            .O(N__11619),
            .I(N__11613));
    CascadeMux I__2236 (
            .O(N__11616),
            .I(N__11610));
    InMux I__2235 (
            .O(N__11613),
            .I(N__11607));
    CascadeBuf I__2234 (
            .O(N__11610),
            .I(N__11604));
    LocalMux I__2233 (
            .O(N__11607),
            .I(N__11601));
    CascadeMux I__2232 (
            .O(N__11604),
            .I(N__11598));
    Span4Mux_h I__2231 (
            .O(N__11601),
            .I(N__11595));
    InMux I__2230 (
            .O(N__11598),
            .I(N__11592));
    Sp12to4 I__2229 (
            .O(N__11595),
            .I(N__11589));
    LocalMux I__2228 (
            .O(N__11592),
            .I(N__11586));
    Span12Mux_h I__2227 (
            .O(N__11589),
            .I(N__11581));
    Span12Mux_s10_h I__2226 (
            .O(N__11586),
            .I(N__11581));
    Span12Mux_v I__2225 (
            .O(N__11581),
            .I(N__11578));
    Odrv12 I__2224 (
            .O(N__11578),
            .I(n21));
    InMux I__2223 (
            .O(N__11575),
            .I(N__11572));
    LocalMux I__2222 (
            .O(N__11572),
            .I(N__11568));
    InMux I__2221 (
            .O(N__11571),
            .I(N__11565));
    Span4Mux_v I__2220 (
            .O(N__11568),
            .I(N__11562));
    LocalMux I__2219 (
            .O(N__11565),
            .I(\transmit_module.n385 ));
    Odrv4 I__2218 (
            .O(N__11562),
            .I(\transmit_module.n385 ));
    IoInMux I__2217 (
            .O(N__11557),
            .I(N__11554));
    LocalMux I__2216 (
            .O(N__11554),
            .I(N__11551));
    Span4Mux_s3_h I__2215 (
            .O(N__11551),
            .I(N__11548));
    Span4Mux_v I__2214 (
            .O(N__11548),
            .I(N__11545));
    Span4Mux_h I__2213 (
            .O(N__11545),
            .I(N__11542));
    Span4Mux_h I__2212 (
            .O(N__11542),
            .I(N__11537));
    CascadeMux I__2211 (
            .O(N__11541),
            .I(N__11534));
    InMux I__2210 (
            .O(N__11540),
            .I(N__11531));
    Span4Mux_h I__2209 (
            .O(N__11537),
            .I(N__11527));
    InMux I__2208 (
            .O(N__11534),
            .I(N__11524));
    LocalMux I__2207 (
            .O(N__11531),
            .I(N__11521));
    InMux I__2206 (
            .O(N__11530),
            .I(N__11518));
    Odrv4 I__2205 (
            .O(N__11527),
            .I(DEBUG_c_3));
    LocalMux I__2204 (
            .O(N__11524),
            .I(DEBUG_c_3));
    Odrv4 I__2203 (
            .O(N__11521),
            .I(DEBUG_c_3));
    LocalMux I__2202 (
            .O(N__11518),
            .I(DEBUG_c_3));
    CascadeMux I__2201 (
            .O(N__11509),
            .I(N__11505));
    CascadeMux I__2200 (
            .O(N__11508),
            .I(N__11502));
    CascadeBuf I__2199 (
            .O(N__11505),
            .I(N__11499));
    CascadeBuf I__2198 (
            .O(N__11502),
            .I(N__11496));
    CascadeMux I__2197 (
            .O(N__11499),
            .I(N__11493));
    CascadeMux I__2196 (
            .O(N__11496),
            .I(N__11490));
    CascadeBuf I__2195 (
            .O(N__11493),
            .I(N__11487));
    CascadeBuf I__2194 (
            .O(N__11490),
            .I(N__11484));
    CascadeMux I__2193 (
            .O(N__11487),
            .I(N__11481));
    CascadeMux I__2192 (
            .O(N__11484),
            .I(N__11478));
    CascadeBuf I__2191 (
            .O(N__11481),
            .I(N__11475));
    CascadeBuf I__2190 (
            .O(N__11478),
            .I(N__11472));
    CascadeMux I__2189 (
            .O(N__11475),
            .I(N__11469));
    CascadeMux I__2188 (
            .O(N__11472),
            .I(N__11466));
    CascadeBuf I__2187 (
            .O(N__11469),
            .I(N__11463));
    CascadeBuf I__2186 (
            .O(N__11466),
            .I(N__11460));
    CascadeMux I__2185 (
            .O(N__11463),
            .I(N__11457));
    CascadeMux I__2184 (
            .O(N__11460),
            .I(N__11454));
    CascadeBuf I__2183 (
            .O(N__11457),
            .I(N__11451));
    CascadeBuf I__2182 (
            .O(N__11454),
            .I(N__11448));
    CascadeMux I__2181 (
            .O(N__11451),
            .I(N__11445));
    CascadeMux I__2180 (
            .O(N__11448),
            .I(N__11442));
    CascadeBuf I__2179 (
            .O(N__11445),
            .I(N__11439));
    CascadeBuf I__2178 (
            .O(N__11442),
            .I(N__11436));
    CascadeMux I__2177 (
            .O(N__11439),
            .I(N__11433));
    CascadeMux I__2176 (
            .O(N__11436),
            .I(N__11430));
    CascadeBuf I__2175 (
            .O(N__11433),
            .I(N__11427));
    CascadeBuf I__2174 (
            .O(N__11430),
            .I(N__11424));
    CascadeMux I__2173 (
            .O(N__11427),
            .I(N__11421));
    CascadeMux I__2172 (
            .O(N__11424),
            .I(N__11418));
    CascadeBuf I__2171 (
            .O(N__11421),
            .I(N__11415));
    CascadeBuf I__2170 (
            .O(N__11418),
            .I(N__11412));
    CascadeMux I__2169 (
            .O(N__11415),
            .I(N__11409));
    CascadeMux I__2168 (
            .O(N__11412),
            .I(N__11406));
    CascadeBuf I__2167 (
            .O(N__11409),
            .I(N__11403));
    CascadeBuf I__2166 (
            .O(N__11406),
            .I(N__11400));
    CascadeMux I__2165 (
            .O(N__11403),
            .I(N__11397));
    CascadeMux I__2164 (
            .O(N__11400),
            .I(N__11394));
    CascadeBuf I__2163 (
            .O(N__11397),
            .I(N__11391));
    CascadeBuf I__2162 (
            .O(N__11394),
            .I(N__11388));
    CascadeMux I__2161 (
            .O(N__11391),
            .I(N__11385));
    CascadeMux I__2160 (
            .O(N__11388),
            .I(N__11382));
    CascadeBuf I__2159 (
            .O(N__11385),
            .I(N__11379));
    CascadeBuf I__2158 (
            .O(N__11382),
            .I(N__11376));
    CascadeMux I__2157 (
            .O(N__11379),
            .I(N__11373));
    CascadeMux I__2156 (
            .O(N__11376),
            .I(N__11370));
    CascadeBuf I__2155 (
            .O(N__11373),
            .I(N__11367));
    CascadeBuf I__2154 (
            .O(N__11370),
            .I(N__11364));
    CascadeMux I__2153 (
            .O(N__11367),
            .I(N__11361));
    CascadeMux I__2152 (
            .O(N__11364),
            .I(N__11358));
    CascadeBuf I__2151 (
            .O(N__11361),
            .I(N__11355));
    CascadeBuf I__2150 (
            .O(N__11358),
            .I(N__11352));
    CascadeMux I__2149 (
            .O(N__11355),
            .I(N__11349));
    CascadeMux I__2148 (
            .O(N__11352),
            .I(N__11346));
    CascadeBuf I__2147 (
            .O(N__11349),
            .I(N__11343));
    CascadeBuf I__2146 (
            .O(N__11346),
            .I(N__11340));
    CascadeMux I__2145 (
            .O(N__11343),
            .I(N__11337));
    CascadeMux I__2144 (
            .O(N__11340),
            .I(N__11334));
    CascadeBuf I__2143 (
            .O(N__11337),
            .I(N__11331));
    CascadeBuf I__2142 (
            .O(N__11334),
            .I(N__11328));
    CascadeMux I__2141 (
            .O(N__11331),
            .I(N__11325));
    CascadeMux I__2140 (
            .O(N__11328),
            .I(N__11322));
    InMux I__2139 (
            .O(N__11325),
            .I(N__11319));
    InMux I__2138 (
            .O(N__11322),
            .I(N__11316));
    LocalMux I__2137 (
            .O(N__11319),
            .I(N__11313));
    LocalMux I__2136 (
            .O(N__11316),
            .I(N__11310));
    Span12Mux_h I__2135 (
            .O(N__11313),
            .I(N__11307));
    Sp12to4 I__2134 (
            .O(N__11310),
            .I(N__11304));
    Span12Mux_v I__2133 (
            .O(N__11307),
            .I(N__11299));
    Span12Mux_v I__2132 (
            .O(N__11304),
            .I(N__11299));
    Odrv12 I__2131 (
            .O(N__11299),
            .I(n25_adj_573));
    InMux I__2130 (
            .O(N__11296),
            .I(N__11293));
    LocalMux I__2129 (
            .O(N__11293),
            .I(N__11290));
    Odrv12 I__2128 (
            .O(N__11290),
            .I(\line_buffer.n3028 ));
    CascadeMux I__2127 (
            .O(N__11287),
            .I(\line_buffer.n3125_cascade_ ));
    InMux I__2126 (
            .O(N__11284),
            .I(N__11281));
    LocalMux I__2125 (
            .O(N__11281),
            .I(N__11278));
    Odrv4 I__2124 (
            .O(N__11278),
            .I(TX_DATA_7));
    InMux I__2123 (
            .O(N__11275),
            .I(N__11272));
    LocalMux I__2122 (
            .O(N__11272),
            .I(N__11269));
    Span4Mux_v I__2121 (
            .O(N__11269),
            .I(N__11266));
    Sp12to4 I__2120 (
            .O(N__11266),
            .I(N__11263));
    Odrv12 I__2119 (
            .O(N__11263),
            .I(\line_buffer.n727 ));
    InMux I__2118 (
            .O(N__11260),
            .I(N__11257));
    LocalMux I__2117 (
            .O(N__11257),
            .I(N__11254));
    Span12Mux_v I__2116 (
            .O(N__11254),
            .I(N__11251));
    Span12Mux_v I__2115 (
            .O(N__11251),
            .I(N__11248));
    Odrv12 I__2114 (
            .O(N__11248),
            .I(\line_buffer.n719 ));
    InMux I__2113 (
            .O(N__11245),
            .I(N__11242));
    LocalMux I__2112 (
            .O(N__11242),
            .I(\line_buffer.n3043 ));
    InMux I__2111 (
            .O(N__11239),
            .I(N__11236));
    LocalMux I__2110 (
            .O(N__11236),
            .I(N__11233));
    Span4Mux_v I__2109 (
            .O(N__11233),
            .I(N__11230));
    Span4Mux_h I__2108 (
            .O(N__11230),
            .I(N__11227));
    Span4Mux_h I__2107 (
            .O(N__11227),
            .I(N__11224));
    Span4Mux_v I__2106 (
            .O(N__11224),
            .I(N__11221));
    Odrv4 I__2105 (
            .O(N__11221),
            .I(\line_buffer.n689 ));
    CascadeMux I__2104 (
            .O(N__11218),
            .I(N__11215));
    InMux I__2103 (
            .O(N__11215),
            .I(N__11212));
    LocalMux I__2102 (
            .O(N__11212),
            .I(N__11209));
    Span4Mux_v I__2101 (
            .O(N__11209),
            .I(N__11206));
    Span4Mux_h I__2100 (
            .O(N__11206),
            .I(N__11203));
    Span4Mux_h I__2099 (
            .O(N__11203),
            .I(N__11200));
    Odrv4 I__2098 (
            .O(N__11200),
            .I(\line_buffer.n681 ));
    CascadeMux I__2097 (
            .O(N__11197),
            .I(\line_buffer.n3140_cascade_ ));
    InMux I__2096 (
            .O(N__11194),
            .I(N__11191));
    LocalMux I__2095 (
            .O(N__11191),
            .I(TX_DATA_1));
    InMux I__2094 (
            .O(N__11188),
            .I(N__11185));
    LocalMux I__2093 (
            .O(N__11185),
            .I(N__11182));
    Odrv12 I__2092 (
            .O(N__11182),
            .I(\line_buffer.n713 ));
    InMux I__2091 (
            .O(N__11179),
            .I(N__11176));
    LocalMux I__2090 (
            .O(N__11176),
            .I(N__11173));
    Span4Mux_v I__2089 (
            .O(N__11173),
            .I(N__11170));
    Span4Mux_h I__2088 (
            .O(N__11170),
            .I(N__11167));
    Span4Mux_h I__2087 (
            .O(N__11167),
            .I(N__11164));
    Odrv4 I__2086 (
            .O(N__11164),
            .I(\line_buffer.n721 ));
    InMux I__2085 (
            .O(N__11161),
            .I(N__11158));
    LocalMux I__2084 (
            .O(N__11158),
            .I(N__11155));
    Span12Mux_v I__2083 (
            .O(N__11155),
            .I(N__11152));
    Odrv12 I__2082 (
            .O(N__11152),
            .I(\line_buffer.n624 ));
    InMux I__2081 (
            .O(N__11149),
            .I(N__11146));
    LocalMux I__2080 (
            .O(N__11146),
            .I(N__11143));
    Span12Mux_v I__2079 (
            .O(N__11143),
            .I(N__11140));
    Odrv12 I__2078 (
            .O(N__11140),
            .I(\line_buffer.n616 ));
    CascadeMux I__2077 (
            .O(N__11137),
            .I(\line_buffer.n3107_cascade_ ));
    InMux I__2076 (
            .O(N__11134),
            .I(N__11131));
    LocalMux I__2075 (
            .O(N__11131),
            .I(\line_buffer.n3110 ));
    CascadeMux I__2074 (
            .O(N__11128),
            .I(N__11124));
    CascadeMux I__2073 (
            .O(N__11127),
            .I(N__11121));
    CascadeBuf I__2072 (
            .O(N__11124),
            .I(N__11118));
    CascadeBuf I__2071 (
            .O(N__11121),
            .I(N__11115));
    CascadeMux I__2070 (
            .O(N__11118),
            .I(N__11112));
    CascadeMux I__2069 (
            .O(N__11115),
            .I(N__11109));
    CascadeBuf I__2068 (
            .O(N__11112),
            .I(N__11106));
    CascadeBuf I__2067 (
            .O(N__11109),
            .I(N__11103));
    CascadeMux I__2066 (
            .O(N__11106),
            .I(N__11100));
    CascadeMux I__2065 (
            .O(N__11103),
            .I(N__11097));
    CascadeBuf I__2064 (
            .O(N__11100),
            .I(N__11094));
    CascadeBuf I__2063 (
            .O(N__11097),
            .I(N__11091));
    CascadeMux I__2062 (
            .O(N__11094),
            .I(N__11088));
    CascadeMux I__2061 (
            .O(N__11091),
            .I(N__11085));
    CascadeBuf I__2060 (
            .O(N__11088),
            .I(N__11082));
    CascadeBuf I__2059 (
            .O(N__11085),
            .I(N__11079));
    CascadeMux I__2058 (
            .O(N__11082),
            .I(N__11076));
    CascadeMux I__2057 (
            .O(N__11079),
            .I(N__11073));
    CascadeBuf I__2056 (
            .O(N__11076),
            .I(N__11070));
    CascadeBuf I__2055 (
            .O(N__11073),
            .I(N__11067));
    CascadeMux I__2054 (
            .O(N__11070),
            .I(N__11064));
    CascadeMux I__2053 (
            .O(N__11067),
            .I(N__11061));
    CascadeBuf I__2052 (
            .O(N__11064),
            .I(N__11058));
    CascadeBuf I__2051 (
            .O(N__11061),
            .I(N__11055));
    CascadeMux I__2050 (
            .O(N__11058),
            .I(N__11052));
    CascadeMux I__2049 (
            .O(N__11055),
            .I(N__11049));
    CascadeBuf I__2048 (
            .O(N__11052),
            .I(N__11046));
    CascadeBuf I__2047 (
            .O(N__11049),
            .I(N__11043));
    CascadeMux I__2046 (
            .O(N__11046),
            .I(N__11040));
    CascadeMux I__2045 (
            .O(N__11043),
            .I(N__11037));
    CascadeBuf I__2044 (
            .O(N__11040),
            .I(N__11034));
    CascadeBuf I__2043 (
            .O(N__11037),
            .I(N__11031));
    CascadeMux I__2042 (
            .O(N__11034),
            .I(N__11028));
    CascadeMux I__2041 (
            .O(N__11031),
            .I(N__11025));
    CascadeBuf I__2040 (
            .O(N__11028),
            .I(N__11022));
    CascadeBuf I__2039 (
            .O(N__11025),
            .I(N__11019));
    CascadeMux I__2038 (
            .O(N__11022),
            .I(N__11016));
    CascadeMux I__2037 (
            .O(N__11019),
            .I(N__11013));
    CascadeBuf I__2036 (
            .O(N__11016),
            .I(N__11010));
    CascadeBuf I__2035 (
            .O(N__11013),
            .I(N__11007));
    CascadeMux I__2034 (
            .O(N__11010),
            .I(N__11004));
    CascadeMux I__2033 (
            .O(N__11007),
            .I(N__11001));
    CascadeBuf I__2032 (
            .O(N__11004),
            .I(N__10998));
    CascadeBuf I__2031 (
            .O(N__11001),
            .I(N__10995));
    CascadeMux I__2030 (
            .O(N__10998),
            .I(N__10992));
    CascadeMux I__2029 (
            .O(N__10995),
            .I(N__10989));
    CascadeBuf I__2028 (
            .O(N__10992),
            .I(N__10986));
    CascadeBuf I__2027 (
            .O(N__10989),
            .I(N__10983));
    CascadeMux I__2026 (
            .O(N__10986),
            .I(N__10980));
    CascadeMux I__2025 (
            .O(N__10983),
            .I(N__10977));
    CascadeBuf I__2024 (
            .O(N__10980),
            .I(N__10974));
    CascadeBuf I__2023 (
            .O(N__10977),
            .I(N__10971));
    CascadeMux I__2022 (
            .O(N__10974),
            .I(N__10968));
    CascadeMux I__2021 (
            .O(N__10971),
            .I(N__10965));
    CascadeBuf I__2020 (
            .O(N__10968),
            .I(N__10962));
    CascadeBuf I__2019 (
            .O(N__10965),
            .I(N__10959));
    CascadeMux I__2018 (
            .O(N__10962),
            .I(N__10956));
    CascadeMux I__2017 (
            .O(N__10959),
            .I(N__10953));
    CascadeBuf I__2016 (
            .O(N__10956),
            .I(N__10950));
    CascadeBuf I__2015 (
            .O(N__10953),
            .I(N__10947));
    CascadeMux I__2014 (
            .O(N__10950),
            .I(N__10944));
    CascadeMux I__2013 (
            .O(N__10947),
            .I(N__10941));
    InMux I__2012 (
            .O(N__10944),
            .I(N__10938));
    InMux I__2011 (
            .O(N__10941),
            .I(N__10935));
    LocalMux I__2010 (
            .O(N__10938),
            .I(N__10932));
    LocalMux I__2009 (
            .O(N__10935),
            .I(N__10929));
    Sp12to4 I__2008 (
            .O(N__10932),
            .I(N__10926));
    Span12Mux_s8_h I__2007 (
            .O(N__10929),
            .I(N__10923));
    Span12Mux_s11_h I__2006 (
            .O(N__10926),
            .I(N__10920));
    Span12Mux_v I__2005 (
            .O(N__10923),
            .I(N__10915));
    Span12Mux_v I__2004 (
            .O(N__10920),
            .I(N__10915));
    Odrv12 I__2003 (
            .O(N__10915),
            .I(n19));
    InMux I__2002 (
            .O(N__10912),
            .I(N__10906));
    InMux I__2001 (
            .O(N__10911),
            .I(N__10906));
    LocalMux I__2000 (
            .O(N__10906),
            .I(\transmit_module.n379 ));
    CascadeMux I__1999 (
            .O(N__10903),
            .I(N__10899));
    CascadeMux I__1998 (
            .O(N__10902),
            .I(N__10895));
    InMux I__1997 (
            .O(N__10899),
            .I(N__10890));
    InMux I__1996 (
            .O(N__10898),
            .I(N__10890));
    InMux I__1995 (
            .O(N__10895),
            .I(N__10887));
    LocalMux I__1994 (
            .O(N__10890),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__1993 (
            .O(N__10887),
            .I(\transmit_module.TX_ADDR_9 ));
    InMux I__1992 (
            .O(N__10882),
            .I(N__10877));
    InMux I__1991 (
            .O(N__10881),
            .I(N__10874));
    InMux I__1990 (
            .O(N__10880),
            .I(N__10871));
    LocalMux I__1989 (
            .O(N__10877),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__1988 (
            .O(N__10874),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__1987 (
            .O(N__10871),
            .I(\transmit_module.TX_ADDR_8 ));
    CascadeMux I__1986 (
            .O(N__10864),
            .I(N__10861));
    InMux I__1985 (
            .O(N__10861),
            .I(N__10857));
    InMux I__1984 (
            .O(N__10860),
            .I(N__10854));
    LocalMux I__1983 (
            .O(N__10857),
            .I(\transmit_module.n380 ));
    LocalMux I__1982 (
            .O(N__10854),
            .I(\transmit_module.n380 ));
    CascadeMux I__1981 (
            .O(N__10849),
            .I(N__10846));
    CascadeBuf I__1980 (
            .O(N__10846),
            .I(N__10842));
    CascadeMux I__1979 (
            .O(N__10845),
            .I(N__10839));
    CascadeMux I__1978 (
            .O(N__10842),
            .I(N__10836));
    CascadeBuf I__1977 (
            .O(N__10839),
            .I(N__10833));
    CascadeBuf I__1976 (
            .O(N__10836),
            .I(N__10830));
    CascadeMux I__1975 (
            .O(N__10833),
            .I(N__10827));
    CascadeMux I__1974 (
            .O(N__10830),
            .I(N__10824));
    CascadeBuf I__1973 (
            .O(N__10827),
            .I(N__10821));
    CascadeBuf I__1972 (
            .O(N__10824),
            .I(N__10818));
    CascadeMux I__1971 (
            .O(N__10821),
            .I(N__10815));
    CascadeMux I__1970 (
            .O(N__10818),
            .I(N__10812));
    CascadeBuf I__1969 (
            .O(N__10815),
            .I(N__10809));
    CascadeBuf I__1968 (
            .O(N__10812),
            .I(N__10806));
    CascadeMux I__1967 (
            .O(N__10809),
            .I(N__10803));
    CascadeMux I__1966 (
            .O(N__10806),
            .I(N__10800));
    CascadeBuf I__1965 (
            .O(N__10803),
            .I(N__10797));
    CascadeBuf I__1964 (
            .O(N__10800),
            .I(N__10794));
    CascadeMux I__1963 (
            .O(N__10797),
            .I(N__10791));
    CascadeMux I__1962 (
            .O(N__10794),
            .I(N__10788));
    CascadeBuf I__1961 (
            .O(N__10791),
            .I(N__10785));
    CascadeBuf I__1960 (
            .O(N__10788),
            .I(N__10782));
    CascadeMux I__1959 (
            .O(N__10785),
            .I(N__10779));
    CascadeMux I__1958 (
            .O(N__10782),
            .I(N__10776));
    CascadeBuf I__1957 (
            .O(N__10779),
            .I(N__10773));
    CascadeBuf I__1956 (
            .O(N__10776),
            .I(N__10770));
    CascadeMux I__1955 (
            .O(N__10773),
            .I(N__10767));
    CascadeMux I__1954 (
            .O(N__10770),
            .I(N__10764));
    CascadeBuf I__1953 (
            .O(N__10767),
            .I(N__10761));
    CascadeBuf I__1952 (
            .O(N__10764),
            .I(N__10758));
    CascadeMux I__1951 (
            .O(N__10761),
            .I(N__10755));
    CascadeMux I__1950 (
            .O(N__10758),
            .I(N__10752));
    CascadeBuf I__1949 (
            .O(N__10755),
            .I(N__10749));
    CascadeBuf I__1948 (
            .O(N__10752),
            .I(N__10746));
    CascadeMux I__1947 (
            .O(N__10749),
            .I(N__10743));
    CascadeMux I__1946 (
            .O(N__10746),
            .I(N__10740));
    CascadeBuf I__1945 (
            .O(N__10743),
            .I(N__10737));
    CascadeBuf I__1944 (
            .O(N__10740),
            .I(N__10734));
    CascadeMux I__1943 (
            .O(N__10737),
            .I(N__10731));
    CascadeMux I__1942 (
            .O(N__10734),
            .I(N__10728));
    CascadeBuf I__1941 (
            .O(N__10731),
            .I(N__10725));
    CascadeBuf I__1940 (
            .O(N__10728),
            .I(N__10722));
    CascadeMux I__1939 (
            .O(N__10725),
            .I(N__10719));
    CascadeMux I__1938 (
            .O(N__10722),
            .I(N__10716));
    CascadeBuf I__1937 (
            .O(N__10719),
            .I(N__10713));
    CascadeBuf I__1936 (
            .O(N__10716),
            .I(N__10710));
    CascadeMux I__1935 (
            .O(N__10713),
            .I(N__10707));
    CascadeMux I__1934 (
            .O(N__10710),
            .I(N__10704));
    CascadeBuf I__1933 (
            .O(N__10707),
            .I(N__10701));
    CascadeBuf I__1932 (
            .O(N__10704),
            .I(N__10698));
    CascadeMux I__1931 (
            .O(N__10701),
            .I(N__10695));
    CascadeMux I__1930 (
            .O(N__10698),
            .I(N__10692));
    CascadeBuf I__1929 (
            .O(N__10695),
            .I(N__10689));
    CascadeBuf I__1928 (
            .O(N__10692),
            .I(N__10686));
    CascadeMux I__1927 (
            .O(N__10689),
            .I(N__10683));
    CascadeMux I__1926 (
            .O(N__10686),
            .I(N__10680));
    CascadeBuf I__1925 (
            .O(N__10683),
            .I(N__10677));
    CascadeBuf I__1924 (
            .O(N__10680),
            .I(N__10674));
    CascadeMux I__1923 (
            .O(N__10677),
            .I(N__10671));
    CascadeMux I__1922 (
            .O(N__10674),
            .I(N__10668));
    CascadeBuf I__1921 (
            .O(N__10671),
            .I(N__10665));
    InMux I__1920 (
            .O(N__10668),
            .I(N__10662));
    CascadeMux I__1919 (
            .O(N__10665),
            .I(N__10659));
    LocalMux I__1918 (
            .O(N__10662),
            .I(N__10656));
    InMux I__1917 (
            .O(N__10659),
            .I(N__10653));
    Span12Mux_h I__1916 (
            .O(N__10656),
            .I(N__10650));
    LocalMux I__1915 (
            .O(N__10653),
            .I(N__10647));
    Span12Mux_v I__1914 (
            .O(N__10650),
            .I(N__10642));
    Span12Mux_v I__1913 (
            .O(N__10647),
            .I(N__10642));
    Odrv12 I__1912 (
            .O(N__10642),
            .I(n20));
    InMux I__1911 (
            .O(N__10639),
            .I(N__10636));
    LocalMux I__1910 (
            .O(N__10636),
            .I(N__10631));
    CascadeMux I__1909 (
            .O(N__10635),
            .I(N__10628));
    InMux I__1908 (
            .O(N__10634),
            .I(N__10625));
    Span4Mux_v I__1907 (
            .O(N__10631),
            .I(N__10622));
    InMux I__1906 (
            .O(N__10628),
            .I(N__10619));
    LocalMux I__1905 (
            .O(N__10625),
            .I(\transmit_module.TX_ADDR_10 ));
    Odrv4 I__1904 (
            .O(N__10622),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__1903 (
            .O(N__10619),
            .I(\transmit_module.TX_ADDR_10 ));
    CascadeMux I__1902 (
            .O(N__10612),
            .I(N__10609));
    InMux I__1901 (
            .O(N__10609),
            .I(N__10605));
    InMux I__1900 (
            .O(N__10608),
            .I(N__10602));
    LocalMux I__1899 (
            .O(N__10605),
            .I(\transmit_module.n378 ));
    LocalMux I__1898 (
            .O(N__10602),
            .I(\transmit_module.n378 ));
    CascadeMux I__1897 (
            .O(N__10597),
            .I(N__10594));
    CascadeBuf I__1896 (
            .O(N__10594),
            .I(N__10590));
    CascadeMux I__1895 (
            .O(N__10593),
            .I(N__10587));
    CascadeMux I__1894 (
            .O(N__10590),
            .I(N__10584));
    CascadeBuf I__1893 (
            .O(N__10587),
            .I(N__10581));
    CascadeBuf I__1892 (
            .O(N__10584),
            .I(N__10578));
    CascadeMux I__1891 (
            .O(N__10581),
            .I(N__10575));
    CascadeMux I__1890 (
            .O(N__10578),
            .I(N__10572));
    CascadeBuf I__1889 (
            .O(N__10575),
            .I(N__10569));
    CascadeBuf I__1888 (
            .O(N__10572),
            .I(N__10566));
    CascadeMux I__1887 (
            .O(N__10569),
            .I(N__10563));
    CascadeMux I__1886 (
            .O(N__10566),
            .I(N__10560));
    CascadeBuf I__1885 (
            .O(N__10563),
            .I(N__10557));
    CascadeBuf I__1884 (
            .O(N__10560),
            .I(N__10554));
    CascadeMux I__1883 (
            .O(N__10557),
            .I(N__10551));
    CascadeMux I__1882 (
            .O(N__10554),
            .I(N__10548));
    CascadeBuf I__1881 (
            .O(N__10551),
            .I(N__10545));
    CascadeBuf I__1880 (
            .O(N__10548),
            .I(N__10542));
    CascadeMux I__1879 (
            .O(N__10545),
            .I(N__10539));
    CascadeMux I__1878 (
            .O(N__10542),
            .I(N__10536));
    CascadeBuf I__1877 (
            .O(N__10539),
            .I(N__10533));
    CascadeBuf I__1876 (
            .O(N__10536),
            .I(N__10530));
    CascadeMux I__1875 (
            .O(N__10533),
            .I(N__10527));
    CascadeMux I__1874 (
            .O(N__10530),
            .I(N__10524));
    CascadeBuf I__1873 (
            .O(N__10527),
            .I(N__10521));
    CascadeBuf I__1872 (
            .O(N__10524),
            .I(N__10518));
    CascadeMux I__1871 (
            .O(N__10521),
            .I(N__10515));
    CascadeMux I__1870 (
            .O(N__10518),
            .I(N__10512));
    CascadeBuf I__1869 (
            .O(N__10515),
            .I(N__10509));
    CascadeBuf I__1868 (
            .O(N__10512),
            .I(N__10506));
    CascadeMux I__1867 (
            .O(N__10509),
            .I(N__10503));
    CascadeMux I__1866 (
            .O(N__10506),
            .I(N__10500));
    CascadeBuf I__1865 (
            .O(N__10503),
            .I(N__10497));
    CascadeBuf I__1864 (
            .O(N__10500),
            .I(N__10494));
    CascadeMux I__1863 (
            .O(N__10497),
            .I(N__10491));
    CascadeMux I__1862 (
            .O(N__10494),
            .I(N__10488));
    CascadeBuf I__1861 (
            .O(N__10491),
            .I(N__10485));
    CascadeBuf I__1860 (
            .O(N__10488),
            .I(N__10482));
    CascadeMux I__1859 (
            .O(N__10485),
            .I(N__10479));
    CascadeMux I__1858 (
            .O(N__10482),
            .I(N__10476));
    CascadeBuf I__1857 (
            .O(N__10479),
            .I(N__10473));
    CascadeBuf I__1856 (
            .O(N__10476),
            .I(N__10470));
    CascadeMux I__1855 (
            .O(N__10473),
            .I(N__10467));
    CascadeMux I__1854 (
            .O(N__10470),
            .I(N__10464));
    CascadeBuf I__1853 (
            .O(N__10467),
            .I(N__10461));
    CascadeBuf I__1852 (
            .O(N__10464),
            .I(N__10458));
    CascadeMux I__1851 (
            .O(N__10461),
            .I(N__10455));
    CascadeMux I__1850 (
            .O(N__10458),
            .I(N__10452));
    CascadeBuf I__1849 (
            .O(N__10455),
            .I(N__10449));
    CascadeBuf I__1848 (
            .O(N__10452),
            .I(N__10446));
    CascadeMux I__1847 (
            .O(N__10449),
            .I(N__10443));
    CascadeMux I__1846 (
            .O(N__10446),
            .I(N__10440));
    CascadeBuf I__1845 (
            .O(N__10443),
            .I(N__10437));
    CascadeBuf I__1844 (
            .O(N__10440),
            .I(N__10434));
    CascadeMux I__1843 (
            .O(N__10437),
            .I(N__10431));
    CascadeMux I__1842 (
            .O(N__10434),
            .I(N__10428));
    CascadeBuf I__1841 (
            .O(N__10431),
            .I(N__10425));
    CascadeBuf I__1840 (
            .O(N__10428),
            .I(N__10422));
    CascadeMux I__1839 (
            .O(N__10425),
            .I(N__10419));
    CascadeMux I__1838 (
            .O(N__10422),
            .I(N__10416));
    CascadeBuf I__1837 (
            .O(N__10419),
            .I(N__10413));
    InMux I__1836 (
            .O(N__10416),
            .I(N__10410));
    CascadeMux I__1835 (
            .O(N__10413),
            .I(N__10407));
    LocalMux I__1834 (
            .O(N__10410),
            .I(N__10404));
    InMux I__1833 (
            .O(N__10407),
            .I(N__10401));
    Sp12to4 I__1832 (
            .O(N__10404),
            .I(N__10398));
    LocalMux I__1831 (
            .O(N__10401),
            .I(N__10395));
    Span12Mux_h I__1830 (
            .O(N__10398),
            .I(N__10392));
    Span12Mux_v I__1829 (
            .O(N__10395),
            .I(N__10387));
    Span12Mux_v I__1828 (
            .O(N__10392),
            .I(N__10387));
    Odrv12 I__1827 (
            .O(N__10387),
            .I(n18));
    InMux I__1826 (
            .O(N__10384),
            .I(N__10381));
    LocalMux I__1825 (
            .O(N__10381),
            .I(N__10378));
    Odrv4 I__1824 (
            .O(N__10378),
            .I(\line_buffer.n3104 ));
    InMux I__1823 (
            .O(N__10375),
            .I(N__10372));
    LocalMux I__1822 (
            .O(N__10372),
            .I(N__10369));
    Odrv12 I__1821 (
            .O(N__10369),
            .I(TX_DATA_6));
    IoInMux I__1820 (
            .O(N__10366),
            .I(N__10363));
    LocalMux I__1819 (
            .O(N__10363),
            .I(N__10360));
    IoSpan4Mux I__1818 (
            .O(N__10360),
            .I(N__10357));
    Span4Mux_s0_v I__1817 (
            .O(N__10357),
            .I(N__10354));
    Odrv4 I__1816 (
            .O(N__10354),
            .I(GB_BUFFER_TVP_CLK_c_THRU_CO));
    InMux I__1815 (
            .O(N__10351),
            .I(N__10348));
    LocalMux I__1814 (
            .O(N__10348),
            .I(\receive_module.old_VS ));
    CEMux I__1813 (
            .O(N__10345),
            .I(N__10342));
    LocalMux I__1812 (
            .O(N__10342),
            .I(N__10338));
    CEMux I__1811 (
            .O(N__10341),
            .I(N__10335));
    Span4Mux_h I__1810 (
            .O(N__10338),
            .I(N__10331));
    LocalMux I__1809 (
            .O(N__10335),
            .I(N__10328));
    InMux I__1808 (
            .O(N__10334),
            .I(N__10325));
    Odrv4 I__1807 (
            .O(N__10331),
            .I(\receive_module.n252 ));
    Odrv12 I__1806 (
            .O(N__10328),
            .I(\receive_module.n252 ));
    LocalMux I__1805 (
            .O(N__10325),
            .I(\receive_module.n252 ));
    IoInMux I__1804 (
            .O(N__10318),
            .I(N__10315));
    LocalMux I__1803 (
            .O(N__10315),
            .I(N__10312));
    Span4Mux_s3_h I__1802 (
            .O(N__10312),
            .I(N__10307));
    IoInMux I__1801 (
            .O(N__10311),
            .I(N__10304));
    IoInMux I__1800 (
            .O(N__10310),
            .I(N__10301));
    Span4Mux_h I__1799 (
            .O(N__10307),
            .I(N__10298));
    LocalMux I__1798 (
            .O(N__10304),
            .I(N__10295));
    LocalMux I__1797 (
            .O(N__10301),
            .I(N__10292));
    Span4Mux_h I__1796 (
            .O(N__10298),
            .I(N__10289));
    Span4Mux_s3_v I__1795 (
            .O(N__10295),
            .I(N__10286));
    Span12Mux_s3_v I__1794 (
            .O(N__10292),
            .I(N__10283));
    Span4Mux_h I__1793 (
            .O(N__10289),
            .I(N__10280));
    Sp12to4 I__1792 (
            .O(N__10286),
            .I(N__10277));
    Span12Mux_h I__1791 (
            .O(N__10283),
            .I(N__10270));
    Sp12to4 I__1790 (
            .O(N__10280),
            .I(N__10270));
    Span12Mux_h I__1789 (
            .O(N__10277),
            .I(N__10270));
    Span12Mux_v I__1788 (
            .O(N__10270),
            .I(N__10267));
    Odrv12 I__1787 (
            .O(N__10267),
            .I(n1950));
    IoInMux I__1786 (
            .O(N__10264),
            .I(N__10261));
    LocalMux I__1785 (
            .O(N__10261),
            .I(N__10258));
    IoSpan4Mux I__1784 (
            .O(N__10258),
            .I(N__10253));
    IoInMux I__1783 (
            .O(N__10257),
            .I(N__10250));
    IoInMux I__1782 (
            .O(N__10256),
            .I(N__10247));
    Span4Mux_s1_v I__1781 (
            .O(N__10253),
            .I(N__10244));
    LocalMux I__1780 (
            .O(N__10250),
            .I(N__10241));
    LocalMux I__1779 (
            .O(N__10247),
            .I(N__10238));
    Span4Mux_v I__1778 (
            .O(N__10244),
            .I(N__10233));
    Span4Mux_s3_h I__1777 (
            .O(N__10241),
            .I(N__10233));
    Span4Mux_s3_v I__1776 (
            .O(N__10238),
            .I(N__10230));
    Sp12to4 I__1775 (
            .O(N__10233),
            .I(N__10227));
    Span4Mux_v I__1774 (
            .O(N__10230),
            .I(N__10224));
    Span12Mux_s7_v I__1773 (
            .O(N__10227),
            .I(N__10221));
    Span4Mux_v I__1772 (
            .O(N__10224),
            .I(N__10218));
    Span12Mux_h I__1771 (
            .O(N__10221),
            .I(N__10215));
    Span4Mux_v I__1770 (
            .O(N__10218),
            .I(N__10212));
    Odrv12 I__1769 (
            .O(N__10215),
            .I(n1954));
    Odrv4 I__1768 (
            .O(N__10212),
            .I(n1954));
    InMux I__1767 (
            .O(N__10207),
            .I(N__10204));
    LocalMux I__1766 (
            .O(N__10204),
            .I(N__10201));
    Odrv4 I__1765 (
            .O(N__10201),
            .I(TX_DATA_3));
    IoInMux I__1764 (
            .O(N__10198),
            .I(N__10193));
    IoInMux I__1763 (
            .O(N__10197),
            .I(N__10190));
    IoInMux I__1762 (
            .O(N__10196),
            .I(N__10187));
    LocalMux I__1761 (
            .O(N__10193),
            .I(N__10184));
    LocalMux I__1760 (
            .O(N__10190),
            .I(N__10181));
    LocalMux I__1759 (
            .O(N__10187),
            .I(N__10178));
    Span4Mux_s3_v I__1758 (
            .O(N__10184),
            .I(N__10175));
    Span4Mux_s3_v I__1757 (
            .O(N__10181),
            .I(N__10172));
    Span4Mux_s3_h I__1756 (
            .O(N__10178),
            .I(N__10169));
    Sp12to4 I__1755 (
            .O(N__10175),
            .I(N__10166));
    Sp12to4 I__1754 (
            .O(N__10172),
            .I(N__10163));
    Sp12to4 I__1753 (
            .O(N__10169),
            .I(N__10160));
    Span12Mux_s8_h I__1752 (
            .O(N__10166),
            .I(N__10157));
    Span12Mux_s11_h I__1751 (
            .O(N__10163),
            .I(N__10154));
    Span12Mux_v I__1750 (
            .O(N__10160),
            .I(N__10151));
    Span12Mux_v I__1749 (
            .O(N__10157),
            .I(N__10146));
    Span12Mux_v I__1748 (
            .O(N__10154),
            .I(N__10146));
    Span12Mux_h I__1747 (
            .O(N__10151),
            .I(N__10143));
    Odrv12 I__1746 (
            .O(N__10146),
            .I(n1952));
    Odrv12 I__1745 (
            .O(N__10143),
            .I(n1952));
    IoInMux I__1744 (
            .O(N__10138),
            .I(N__10134));
    IoInMux I__1743 (
            .O(N__10137),
            .I(N__10131));
    LocalMux I__1742 (
            .O(N__10134),
            .I(N__10128));
    LocalMux I__1741 (
            .O(N__10131),
            .I(N__10124));
    IoSpan4Mux I__1740 (
            .O(N__10128),
            .I(N__10121));
    IoInMux I__1739 (
            .O(N__10127),
            .I(N__10118));
    IoSpan4Mux I__1738 (
            .O(N__10124),
            .I(N__10115));
    Span4Mux_s3_v I__1737 (
            .O(N__10121),
            .I(N__10112));
    LocalMux I__1736 (
            .O(N__10118),
            .I(N__10109));
    Span4Mux_s3_v I__1735 (
            .O(N__10115),
            .I(N__10106));
    Span4Mux_v I__1734 (
            .O(N__10112),
            .I(N__10101));
    Span4Mux_s3_h I__1733 (
            .O(N__10109),
            .I(N__10101));
    Span4Mux_v I__1732 (
            .O(N__10106),
            .I(N__10098));
    Sp12to4 I__1731 (
            .O(N__10101),
            .I(N__10095));
    Sp12to4 I__1730 (
            .O(N__10098),
            .I(N__10092));
    Span12Mux_v I__1729 (
            .O(N__10095),
            .I(N__10089));
    Span12Mux_v I__1728 (
            .O(N__10092),
            .I(N__10084));
    Span12Mux_h I__1727 (
            .O(N__10089),
            .I(N__10084));
    Odrv12 I__1726 (
            .O(N__10084),
            .I(n1951));
    IoInMux I__1725 (
            .O(N__10081),
            .I(N__10078));
    LocalMux I__1724 (
            .O(N__10078),
            .I(N__10073));
    IoInMux I__1723 (
            .O(N__10077),
            .I(N__10070));
    IoInMux I__1722 (
            .O(N__10076),
            .I(N__10067));
    IoSpan4Mux I__1721 (
            .O(N__10073),
            .I(N__10064));
    LocalMux I__1720 (
            .O(N__10070),
            .I(N__10061));
    LocalMux I__1719 (
            .O(N__10067),
            .I(N__10058));
    Span4Mux_s1_h I__1718 (
            .O(N__10064),
            .I(N__10055));
    Span4Mux_s3_v I__1717 (
            .O(N__10061),
            .I(N__10052));
    Span12Mux_s3_v I__1716 (
            .O(N__10058),
            .I(N__10049));
    Sp12to4 I__1715 (
            .O(N__10055),
            .I(N__10046));
    Span4Mux_h I__1714 (
            .O(N__10052),
            .I(N__10043));
    Span12Mux_v I__1713 (
            .O(N__10049),
            .I(N__10040));
    Span12Mux_v I__1712 (
            .O(N__10046),
            .I(N__10037));
    Sp12to4 I__1711 (
            .O(N__10043),
            .I(N__10034));
    Span12Mux_h I__1710 (
            .O(N__10040),
            .I(N__10031));
    Span12Mux_h I__1709 (
            .O(N__10037),
            .I(N__10026));
    Span12Mux_v I__1708 (
            .O(N__10034),
            .I(N__10026));
    Odrv12 I__1707 (
            .O(N__10031),
            .I(n1949));
    Odrv12 I__1706 (
            .O(N__10026),
            .I(n1949));
    IoInMux I__1705 (
            .O(N__10021),
            .I(N__10016));
    IoInMux I__1704 (
            .O(N__10020),
            .I(N__10013));
    IoInMux I__1703 (
            .O(N__10019),
            .I(N__10010));
    LocalMux I__1702 (
            .O(N__10016),
            .I(N__10007));
    LocalMux I__1701 (
            .O(N__10013),
            .I(N__10004));
    LocalMux I__1700 (
            .O(N__10010),
            .I(N__10001));
    Span4Mux_s3_v I__1699 (
            .O(N__10007),
            .I(N__9998));
    Span4Mux_s0_h I__1698 (
            .O(N__10004),
            .I(N__9995));
    Span4Mux_s3_v I__1697 (
            .O(N__10001),
            .I(N__9992));
    Sp12to4 I__1696 (
            .O(N__9998),
            .I(N__9989));
    Sp12to4 I__1695 (
            .O(N__9995),
            .I(N__9986));
    Sp12to4 I__1694 (
            .O(N__9992),
            .I(N__9983));
    Span12Mux_s7_h I__1693 (
            .O(N__9989),
            .I(N__9980));
    Span12Mux_v I__1692 (
            .O(N__9986),
            .I(N__9977));
    Span12Mux_h I__1691 (
            .O(N__9983),
            .I(N__9974));
    Span12Mux_v I__1690 (
            .O(N__9980),
            .I(N__9967));
    Span12Mux_h I__1689 (
            .O(N__9977),
            .I(N__9967));
    Span12Mux_v I__1688 (
            .O(N__9974),
            .I(N__9967));
    Odrv12 I__1687 (
            .O(N__9967),
            .I(ADV_B_c));
    InMux I__1686 (
            .O(N__9964),
            .I(\transmit_module.n2752 ));
    CEMux I__1685 (
            .O(N__9961),
            .I(N__9957));
    CEMux I__1684 (
            .O(N__9960),
            .I(N__9952));
    LocalMux I__1683 (
            .O(N__9957),
            .I(N__9949));
    CEMux I__1682 (
            .O(N__9956),
            .I(N__9946));
    CEMux I__1681 (
            .O(N__9955),
            .I(N__9943));
    LocalMux I__1680 (
            .O(N__9952),
            .I(\transmit_module.n2200 ));
    Odrv12 I__1679 (
            .O(N__9949),
            .I(\transmit_module.n2200 ));
    LocalMux I__1678 (
            .O(N__9946),
            .I(\transmit_module.n2200 ));
    LocalMux I__1677 (
            .O(N__9943),
            .I(\transmit_module.n2200 ));
    IoInMux I__1676 (
            .O(N__9934),
            .I(N__9931));
    LocalMux I__1675 (
            .O(N__9931),
            .I(N__9926));
    CascadeMux I__1674 (
            .O(N__9930),
            .I(N__9923));
    CascadeMux I__1673 (
            .O(N__9929),
            .I(N__9919));
    Span12Mux_s5_h I__1672 (
            .O(N__9926),
            .I(N__9916));
    InMux I__1671 (
            .O(N__9923),
            .I(N__9913));
    InMux I__1670 (
            .O(N__9922),
            .I(N__9910));
    InMux I__1669 (
            .O(N__9919),
            .I(N__9907));
    Odrv12 I__1668 (
            .O(N__9916),
            .I(DEBUG_c_6));
    LocalMux I__1667 (
            .O(N__9913),
            .I(DEBUG_c_6));
    LocalMux I__1666 (
            .O(N__9910),
            .I(DEBUG_c_6));
    LocalMux I__1665 (
            .O(N__9907),
            .I(DEBUG_c_6));
    InMux I__1664 (
            .O(N__9898),
            .I(N__9894));
    InMux I__1663 (
            .O(N__9897),
            .I(N__9891));
    LocalMux I__1662 (
            .O(N__9894),
            .I(N__9888));
    LocalMux I__1661 (
            .O(N__9891),
            .I(\transmit_module.n382 ));
    Odrv4 I__1660 (
            .O(N__9888),
            .I(\transmit_module.n382 ));
    CascadeMux I__1659 (
            .O(N__9883),
            .I(N__9879));
    CascadeMux I__1658 (
            .O(N__9882),
            .I(N__9876));
    CascadeBuf I__1657 (
            .O(N__9879),
            .I(N__9873));
    CascadeBuf I__1656 (
            .O(N__9876),
            .I(N__9870));
    CascadeMux I__1655 (
            .O(N__9873),
            .I(N__9867));
    CascadeMux I__1654 (
            .O(N__9870),
            .I(N__9864));
    CascadeBuf I__1653 (
            .O(N__9867),
            .I(N__9861));
    CascadeBuf I__1652 (
            .O(N__9864),
            .I(N__9858));
    CascadeMux I__1651 (
            .O(N__9861),
            .I(N__9855));
    CascadeMux I__1650 (
            .O(N__9858),
            .I(N__9852));
    CascadeBuf I__1649 (
            .O(N__9855),
            .I(N__9849));
    CascadeBuf I__1648 (
            .O(N__9852),
            .I(N__9846));
    CascadeMux I__1647 (
            .O(N__9849),
            .I(N__9843));
    CascadeMux I__1646 (
            .O(N__9846),
            .I(N__9840));
    CascadeBuf I__1645 (
            .O(N__9843),
            .I(N__9837));
    CascadeBuf I__1644 (
            .O(N__9840),
            .I(N__9834));
    CascadeMux I__1643 (
            .O(N__9837),
            .I(N__9831));
    CascadeMux I__1642 (
            .O(N__9834),
            .I(N__9828));
    CascadeBuf I__1641 (
            .O(N__9831),
            .I(N__9825));
    CascadeBuf I__1640 (
            .O(N__9828),
            .I(N__9822));
    CascadeMux I__1639 (
            .O(N__9825),
            .I(N__9819));
    CascadeMux I__1638 (
            .O(N__9822),
            .I(N__9816));
    CascadeBuf I__1637 (
            .O(N__9819),
            .I(N__9813));
    CascadeBuf I__1636 (
            .O(N__9816),
            .I(N__9810));
    CascadeMux I__1635 (
            .O(N__9813),
            .I(N__9807));
    CascadeMux I__1634 (
            .O(N__9810),
            .I(N__9804));
    CascadeBuf I__1633 (
            .O(N__9807),
            .I(N__9801));
    CascadeBuf I__1632 (
            .O(N__9804),
            .I(N__9798));
    CascadeMux I__1631 (
            .O(N__9801),
            .I(N__9795));
    CascadeMux I__1630 (
            .O(N__9798),
            .I(N__9792));
    CascadeBuf I__1629 (
            .O(N__9795),
            .I(N__9789));
    CascadeBuf I__1628 (
            .O(N__9792),
            .I(N__9786));
    CascadeMux I__1627 (
            .O(N__9789),
            .I(N__9783));
    CascadeMux I__1626 (
            .O(N__9786),
            .I(N__9780));
    CascadeBuf I__1625 (
            .O(N__9783),
            .I(N__9777));
    CascadeBuf I__1624 (
            .O(N__9780),
            .I(N__9774));
    CascadeMux I__1623 (
            .O(N__9777),
            .I(N__9771));
    CascadeMux I__1622 (
            .O(N__9774),
            .I(N__9768));
    CascadeBuf I__1621 (
            .O(N__9771),
            .I(N__9765));
    CascadeBuf I__1620 (
            .O(N__9768),
            .I(N__9762));
    CascadeMux I__1619 (
            .O(N__9765),
            .I(N__9759));
    CascadeMux I__1618 (
            .O(N__9762),
            .I(N__9756));
    CascadeBuf I__1617 (
            .O(N__9759),
            .I(N__9753));
    CascadeBuf I__1616 (
            .O(N__9756),
            .I(N__9750));
    CascadeMux I__1615 (
            .O(N__9753),
            .I(N__9747));
    CascadeMux I__1614 (
            .O(N__9750),
            .I(N__9744));
    CascadeBuf I__1613 (
            .O(N__9747),
            .I(N__9741));
    CascadeBuf I__1612 (
            .O(N__9744),
            .I(N__9738));
    CascadeMux I__1611 (
            .O(N__9741),
            .I(N__9735));
    CascadeMux I__1610 (
            .O(N__9738),
            .I(N__9732));
    CascadeBuf I__1609 (
            .O(N__9735),
            .I(N__9729));
    CascadeBuf I__1608 (
            .O(N__9732),
            .I(N__9726));
    CascadeMux I__1607 (
            .O(N__9729),
            .I(N__9723));
    CascadeMux I__1606 (
            .O(N__9726),
            .I(N__9720));
    CascadeBuf I__1605 (
            .O(N__9723),
            .I(N__9717));
    CascadeBuf I__1604 (
            .O(N__9720),
            .I(N__9714));
    CascadeMux I__1603 (
            .O(N__9717),
            .I(N__9711));
    CascadeMux I__1602 (
            .O(N__9714),
            .I(N__9708));
    CascadeBuf I__1601 (
            .O(N__9711),
            .I(N__9705));
    CascadeBuf I__1600 (
            .O(N__9708),
            .I(N__9702));
    CascadeMux I__1599 (
            .O(N__9705),
            .I(N__9699));
    CascadeMux I__1598 (
            .O(N__9702),
            .I(N__9696));
    InMux I__1597 (
            .O(N__9699),
            .I(N__9693));
    InMux I__1596 (
            .O(N__9696),
            .I(N__9690));
    LocalMux I__1595 (
            .O(N__9693),
            .I(N__9687));
    LocalMux I__1594 (
            .O(N__9690),
            .I(N__9684));
    Span4Mux_v I__1593 (
            .O(N__9687),
            .I(N__9681));
    Span4Mux_h I__1592 (
            .O(N__9684),
            .I(N__9678));
    Span4Mux_h I__1591 (
            .O(N__9681),
            .I(N__9675));
    Sp12to4 I__1590 (
            .O(N__9678),
            .I(N__9672));
    Span4Mux_v I__1589 (
            .O(N__9675),
            .I(N__9669));
    Span12Mux_v I__1588 (
            .O(N__9672),
            .I(N__9666));
    Span4Mux_v I__1587 (
            .O(N__9669),
            .I(N__9663));
    Odrv12 I__1586 (
            .O(N__9666),
            .I(n22));
    Odrv4 I__1585 (
            .O(N__9663),
            .I(n22));
    InMux I__1584 (
            .O(N__9658),
            .I(N__9654));
    InMux I__1583 (
            .O(N__9657),
            .I(N__9651));
    LocalMux I__1582 (
            .O(N__9654),
            .I(N__9648));
    LocalMux I__1581 (
            .O(N__9651),
            .I(\transmit_module.n383 ));
    Odrv4 I__1580 (
            .O(N__9648),
            .I(\transmit_module.n383 ));
    IoInMux I__1579 (
            .O(N__9643),
            .I(N__9640));
    LocalMux I__1578 (
            .O(N__9640),
            .I(N__9637));
    Span4Mux_s2_h I__1577 (
            .O(N__9637),
            .I(N__9634));
    Span4Mux_h I__1576 (
            .O(N__9634),
            .I(N__9631));
    Span4Mux_h I__1575 (
            .O(N__9631),
            .I(N__9627));
    InMux I__1574 (
            .O(N__9630),
            .I(N__9623));
    Span4Mux_h I__1573 (
            .O(N__9627),
            .I(N__9619));
    InMux I__1572 (
            .O(N__9626),
            .I(N__9616));
    LocalMux I__1571 (
            .O(N__9623),
            .I(N__9613));
    InMux I__1570 (
            .O(N__9622),
            .I(N__9610));
    Odrv4 I__1569 (
            .O(N__9619),
            .I(DEBUG_c_5));
    LocalMux I__1568 (
            .O(N__9616),
            .I(DEBUG_c_5));
    Odrv4 I__1567 (
            .O(N__9613),
            .I(DEBUG_c_5));
    LocalMux I__1566 (
            .O(N__9610),
            .I(DEBUG_c_5));
    CascadeMux I__1565 (
            .O(N__9601),
            .I(N__9597));
    CascadeMux I__1564 (
            .O(N__9600),
            .I(N__9594));
    CascadeBuf I__1563 (
            .O(N__9597),
            .I(N__9591));
    CascadeBuf I__1562 (
            .O(N__9594),
            .I(N__9588));
    CascadeMux I__1561 (
            .O(N__9591),
            .I(N__9585));
    CascadeMux I__1560 (
            .O(N__9588),
            .I(N__9582));
    CascadeBuf I__1559 (
            .O(N__9585),
            .I(N__9579));
    CascadeBuf I__1558 (
            .O(N__9582),
            .I(N__9576));
    CascadeMux I__1557 (
            .O(N__9579),
            .I(N__9573));
    CascadeMux I__1556 (
            .O(N__9576),
            .I(N__9570));
    CascadeBuf I__1555 (
            .O(N__9573),
            .I(N__9567));
    CascadeBuf I__1554 (
            .O(N__9570),
            .I(N__9564));
    CascadeMux I__1553 (
            .O(N__9567),
            .I(N__9561));
    CascadeMux I__1552 (
            .O(N__9564),
            .I(N__9558));
    CascadeBuf I__1551 (
            .O(N__9561),
            .I(N__9555));
    CascadeBuf I__1550 (
            .O(N__9558),
            .I(N__9552));
    CascadeMux I__1549 (
            .O(N__9555),
            .I(N__9549));
    CascadeMux I__1548 (
            .O(N__9552),
            .I(N__9546));
    CascadeBuf I__1547 (
            .O(N__9549),
            .I(N__9543));
    CascadeBuf I__1546 (
            .O(N__9546),
            .I(N__9540));
    CascadeMux I__1545 (
            .O(N__9543),
            .I(N__9537));
    CascadeMux I__1544 (
            .O(N__9540),
            .I(N__9534));
    CascadeBuf I__1543 (
            .O(N__9537),
            .I(N__9531));
    CascadeBuf I__1542 (
            .O(N__9534),
            .I(N__9528));
    CascadeMux I__1541 (
            .O(N__9531),
            .I(N__9525));
    CascadeMux I__1540 (
            .O(N__9528),
            .I(N__9522));
    CascadeBuf I__1539 (
            .O(N__9525),
            .I(N__9519));
    CascadeBuf I__1538 (
            .O(N__9522),
            .I(N__9516));
    CascadeMux I__1537 (
            .O(N__9519),
            .I(N__9513));
    CascadeMux I__1536 (
            .O(N__9516),
            .I(N__9510));
    CascadeBuf I__1535 (
            .O(N__9513),
            .I(N__9507));
    CascadeBuf I__1534 (
            .O(N__9510),
            .I(N__9504));
    CascadeMux I__1533 (
            .O(N__9507),
            .I(N__9501));
    CascadeMux I__1532 (
            .O(N__9504),
            .I(N__9498));
    CascadeBuf I__1531 (
            .O(N__9501),
            .I(N__9495));
    CascadeBuf I__1530 (
            .O(N__9498),
            .I(N__9492));
    CascadeMux I__1529 (
            .O(N__9495),
            .I(N__9489));
    CascadeMux I__1528 (
            .O(N__9492),
            .I(N__9486));
    CascadeBuf I__1527 (
            .O(N__9489),
            .I(N__9483));
    CascadeBuf I__1526 (
            .O(N__9486),
            .I(N__9480));
    CascadeMux I__1525 (
            .O(N__9483),
            .I(N__9477));
    CascadeMux I__1524 (
            .O(N__9480),
            .I(N__9474));
    CascadeBuf I__1523 (
            .O(N__9477),
            .I(N__9471));
    CascadeBuf I__1522 (
            .O(N__9474),
            .I(N__9468));
    CascadeMux I__1521 (
            .O(N__9471),
            .I(N__9465));
    CascadeMux I__1520 (
            .O(N__9468),
            .I(N__9462));
    CascadeBuf I__1519 (
            .O(N__9465),
            .I(N__9459));
    CascadeBuf I__1518 (
            .O(N__9462),
            .I(N__9456));
    CascadeMux I__1517 (
            .O(N__9459),
            .I(N__9453));
    CascadeMux I__1516 (
            .O(N__9456),
            .I(N__9450));
    CascadeBuf I__1515 (
            .O(N__9453),
            .I(N__9447));
    CascadeBuf I__1514 (
            .O(N__9450),
            .I(N__9444));
    CascadeMux I__1513 (
            .O(N__9447),
            .I(N__9441));
    CascadeMux I__1512 (
            .O(N__9444),
            .I(N__9438));
    CascadeBuf I__1511 (
            .O(N__9441),
            .I(N__9435));
    CascadeBuf I__1510 (
            .O(N__9438),
            .I(N__9432));
    CascadeMux I__1509 (
            .O(N__9435),
            .I(N__9429));
    CascadeMux I__1508 (
            .O(N__9432),
            .I(N__9426));
    CascadeBuf I__1507 (
            .O(N__9429),
            .I(N__9423));
    CascadeBuf I__1506 (
            .O(N__9426),
            .I(N__9420));
    CascadeMux I__1505 (
            .O(N__9423),
            .I(N__9417));
    CascadeMux I__1504 (
            .O(N__9420),
            .I(N__9414));
    InMux I__1503 (
            .O(N__9417),
            .I(N__9411));
    InMux I__1502 (
            .O(N__9414),
            .I(N__9408));
    LocalMux I__1501 (
            .O(N__9411),
            .I(N__9405));
    LocalMux I__1500 (
            .O(N__9408),
            .I(N__9402));
    Span12Mux_s11_h I__1499 (
            .O(N__9405),
            .I(N__9399));
    Span12Mux_s8_h I__1498 (
            .O(N__9402),
            .I(N__9396));
    Span12Mux_v I__1497 (
            .O(N__9399),
            .I(N__9391));
    Span12Mux_v I__1496 (
            .O(N__9396),
            .I(N__9391));
    Odrv12 I__1495 (
            .O(N__9391),
            .I(n23));
    InMux I__1494 (
            .O(N__9388),
            .I(N__9385));
    LocalMux I__1493 (
            .O(N__9385),
            .I(N__9381));
    InMux I__1492 (
            .O(N__9384),
            .I(N__9378));
    Span4Mux_v I__1491 (
            .O(N__9381),
            .I(N__9375));
    LocalMux I__1490 (
            .O(N__9378),
            .I(\transmit_module.n384 ));
    Odrv4 I__1489 (
            .O(N__9375),
            .I(\transmit_module.n384 ));
    IoInMux I__1488 (
            .O(N__9370),
            .I(N__9367));
    LocalMux I__1487 (
            .O(N__9367),
            .I(N__9363));
    InMux I__1486 (
            .O(N__9366),
            .I(N__9359));
    Span12Mux_s9_h I__1485 (
            .O(N__9363),
            .I(N__9355));
    InMux I__1484 (
            .O(N__9362),
            .I(N__9352));
    LocalMux I__1483 (
            .O(N__9359),
            .I(N__9349));
    InMux I__1482 (
            .O(N__9358),
            .I(N__9346));
    Odrv12 I__1481 (
            .O(N__9355),
            .I(DEBUG_c_4));
    LocalMux I__1480 (
            .O(N__9352),
            .I(DEBUG_c_4));
    Odrv12 I__1479 (
            .O(N__9349),
            .I(DEBUG_c_4));
    LocalMux I__1478 (
            .O(N__9346),
            .I(DEBUG_c_4));
    CascadeMux I__1477 (
            .O(N__9337),
            .I(N__9333));
    CascadeMux I__1476 (
            .O(N__9336),
            .I(N__9330));
    CascadeBuf I__1475 (
            .O(N__9333),
            .I(N__9327));
    CascadeBuf I__1474 (
            .O(N__9330),
            .I(N__9324));
    CascadeMux I__1473 (
            .O(N__9327),
            .I(N__9321));
    CascadeMux I__1472 (
            .O(N__9324),
            .I(N__9318));
    CascadeBuf I__1471 (
            .O(N__9321),
            .I(N__9315));
    CascadeBuf I__1470 (
            .O(N__9318),
            .I(N__9312));
    CascadeMux I__1469 (
            .O(N__9315),
            .I(N__9309));
    CascadeMux I__1468 (
            .O(N__9312),
            .I(N__9306));
    CascadeBuf I__1467 (
            .O(N__9309),
            .I(N__9303));
    CascadeBuf I__1466 (
            .O(N__9306),
            .I(N__9300));
    CascadeMux I__1465 (
            .O(N__9303),
            .I(N__9297));
    CascadeMux I__1464 (
            .O(N__9300),
            .I(N__9294));
    CascadeBuf I__1463 (
            .O(N__9297),
            .I(N__9291));
    CascadeBuf I__1462 (
            .O(N__9294),
            .I(N__9288));
    CascadeMux I__1461 (
            .O(N__9291),
            .I(N__9285));
    CascadeMux I__1460 (
            .O(N__9288),
            .I(N__9282));
    CascadeBuf I__1459 (
            .O(N__9285),
            .I(N__9279));
    CascadeBuf I__1458 (
            .O(N__9282),
            .I(N__9276));
    CascadeMux I__1457 (
            .O(N__9279),
            .I(N__9273));
    CascadeMux I__1456 (
            .O(N__9276),
            .I(N__9270));
    CascadeBuf I__1455 (
            .O(N__9273),
            .I(N__9267));
    CascadeBuf I__1454 (
            .O(N__9270),
            .I(N__9264));
    CascadeMux I__1453 (
            .O(N__9267),
            .I(N__9261));
    CascadeMux I__1452 (
            .O(N__9264),
            .I(N__9258));
    CascadeBuf I__1451 (
            .O(N__9261),
            .I(N__9255));
    CascadeBuf I__1450 (
            .O(N__9258),
            .I(N__9252));
    CascadeMux I__1449 (
            .O(N__9255),
            .I(N__9249));
    CascadeMux I__1448 (
            .O(N__9252),
            .I(N__9246));
    CascadeBuf I__1447 (
            .O(N__9249),
            .I(N__9243));
    CascadeBuf I__1446 (
            .O(N__9246),
            .I(N__9240));
    CascadeMux I__1445 (
            .O(N__9243),
            .I(N__9237));
    CascadeMux I__1444 (
            .O(N__9240),
            .I(N__9234));
    CascadeBuf I__1443 (
            .O(N__9237),
            .I(N__9231));
    CascadeBuf I__1442 (
            .O(N__9234),
            .I(N__9228));
    CascadeMux I__1441 (
            .O(N__9231),
            .I(N__9225));
    CascadeMux I__1440 (
            .O(N__9228),
            .I(N__9222));
    CascadeBuf I__1439 (
            .O(N__9225),
            .I(N__9219));
    CascadeBuf I__1438 (
            .O(N__9222),
            .I(N__9216));
    CascadeMux I__1437 (
            .O(N__9219),
            .I(N__9213));
    CascadeMux I__1436 (
            .O(N__9216),
            .I(N__9210));
    CascadeBuf I__1435 (
            .O(N__9213),
            .I(N__9207));
    CascadeBuf I__1434 (
            .O(N__9210),
            .I(N__9204));
    CascadeMux I__1433 (
            .O(N__9207),
            .I(N__9201));
    CascadeMux I__1432 (
            .O(N__9204),
            .I(N__9198));
    CascadeBuf I__1431 (
            .O(N__9201),
            .I(N__9195));
    CascadeBuf I__1430 (
            .O(N__9198),
            .I(N__9192));
    CascadeMux I__1429 (
            .O(N__9195),
            .I(N__9189));
    CascadeMux I__1428 (
            .O(N__9192),
            .I(N__9186));
    CascadeBuf I__1427 (
            .O(N__9189),
            .I(N__9183));
    CascadeBuf I__1426 (
            .O(N__9186),
            .I(N__9180));
    CascadeMux I__1425 (
            .O(N__9183),
            .I(N__9177));
    CascadeMux I__1424 (
            .O(N__9180),
            .I(N__9174));
    CascadeBuf I__1423 (
            .O(N__9177),
            .I(N__9171));
    CascadeBuf I__1422 (
            .O(N__9174),
            .I(N__9168));
    CascadeMux I__1421 (
            .O(N__9171),
            .I(N__9165));
    CascadeMux I__1420 (
            .O(N__9168),
            .I(N__9162));
    CascadeBuf I__1419 (
            .O(N__9165),
            .I(N__9159));
    CascadeBuf I__1418 (
            .O(N__9162),
            .I(N__9156));
    CascadeMux I__1417 (
            .O(N__9159),
            .I(N__9153));
    CascadeMux I__1416 (
            .O(N__9156),
            .I(N__9150));
    InMux I__1415 (
            .O(N__9153),
            .I(N__9147));
    InMux I__1414 (
            .O(N__9150),
            .I(N__9144));
    LocalMux I__1413 (
            .O(N__9147),
            .I(N__9141));
    LocalMux I__1412 (
            .O(N__9144),
            .I(N__9138));
    Span12Mux_h I__1411 (
            .O(N__9141),
            .I(N__9133));
    Span12Mux_h I__1410 (
            .O(N__9138),
            .I(N__9133));
    Span12Mux_v I__1409 (
            .O(N__9133),
            .I(N__9130));
    Odrv12 I__1408 (
            .O(N__9130),
            .I(n24));
    InMux I__1407 (
            .O(N__9127),
            .I(N__9123));
    InMux I__1406 (
            .O(N__9126),
            .I(N__9120));
    LocalMux I__1405 (
            .O(N__9123),
            .I(N__9117));
    LocalMux I__1404 (
            .O(N__9120),
            .I(\transmit_module.n386 ));
    Odrv12 I__1403 (
            .O(N__9117),
            .I(\transmit_module.n386 ));
    IoInMux I__1402 (
            .O(N__9112),
            .I(N__9109));
    LocalMux I__1401 (
            .O(N__9109),
            .I(N__9106));
    Span4Mux_s1_h I__1400 (
            .O(N__9106),
            .I(N__9103));
    Sp12to4 I__1399 (
            .O(N__9103),
            .I(N__9099));
    InMux I__1398 (
            .O(N__9102),
            .I(N__9096));
    Span12Mux_v I__1397 (
            .O(N__9099),
            .I(N__9093));
    LocalMux I__1396 (
            .O(N__9096),
            .I(N__9089));
    Span12Mux_h I__1395 (
            .O(N__9093),
            .I(N__9085));
    InMux I__1394 (
            .O(N__9092),
            .I(N__9082));
    Span4Mux_v I__1393 (
            .O(N__9089),
            .I(N__9079));
    InMux I__1392 (
            .O(N__9088),
            .I(N__9076));
    Odrv12 I__1391 (
            .O(N__9085),
            .I(DEBUG_c_2));
    LocalMux I__1390 (
            .O(N__9082),
            .I(DEBUG_c_2));
    Odrv4 I__1389 (
            .O(N__9079),
            .I(DEBUG_c_2));
    LocalMux I__1388 (
            .O(N__9076),
            .I(DEBUG_c_2));
    CascadeMux I__1387 (
            .O(N__9067),
            .I(N__9064));
    CascadeBuf I__1386 (
            .O(N__9064),
            .I(N__9061));
    CascadeMux I__1385 (
            .O(N__9061),
            .I(N__9057));
    CascadeMux I__1384 (
            .O(N__9060),
            .I(N__9054));
    CascadeBuf I__1383 (
            .O(N__9057),
            .I(N__9051));
    CascadeBuf I__1382 (
            .O(N__9054),
            .I(N__9048));
    CascadeMux I__1381 (
            .O(N__9051),
            .I(N__9045));
    CascadeMux I__1380 (
            .O(N__9048),
            .I(N__9042));
    CascadeBuf I__1379 (
            .O(N__9045),
            .I(N__9039));
    CascadeBuf I__1378 (
            .O(N__9042),
            .I(N__9036));
    CascadeMux I__1377 (
            .O(N__9039),
            .I(N__9033));
    CascadeMux I__1376 (
            .O(N__9036),
            .I(N__9030));
    CascadeBuf I__1375 (
            .O(N__9033),
            .I(N__9027));
    CascadeBuf I__1374 (
            .O(N__9030),
            .I(N__9024));
    CascadeMux I__1373 (
            .O(N__9027),
            .I(N__9021));
    CascadeMux I__1372 (
            .O(N__9024),
            .I(N__9018));
    CascadeBuf I__1371 (
            .O(N__9021),
            .I(N__9015));
    CascadeBuf I__1370 (
            .O(N__9018),
            .I(N__9012));
    CascadeMux I__1369 (
            .O(N__9015),
            .I(N__9009));
    CascadeMux I__1368 (
            .O(N__9012),
            .I(N__9006));
    CascadeBuf I__1367 (
            .O(N__9009),
            .I(N__9003));
    CascadeBuf I__1366 (
            .O(N__9006),
            .I(N__9000));
    CascadeMux I__1365 (
            .O(N__9003),
            .I(N__8997));
    CascadeMux I__1364 (
            .O(N__9000),
            .I(N__8994));
    CascadeBuf I__1363 (
            .O(N__8997),
            .I(N__8991));
    CascadeBuf I__1362 (
            .O(N__8994),
            .I(N__8988));
    CascadeMux I__1361 (
            .O(N__8991),
            .I(N__8985));
    CascadeMux I__1360 (
            .O(N__8988),
            .I(N__8982));
    CascadeBuf I__1359 (
            .O(N__8985),
            .I(N__8979));
    CascadeBuf I__1358 (
            .O(N__8982),
            .I(N__8976));
    CascadeMux I__1357 (
            .O(N__8979),
            .I(N__8973));
    CascadeMux I__1356 (
            .O(N__8976),
            .I(N__8970));
    CascadeBuf I__1355 (
            .O(N__8973),
            .I(N__8967));
    CascadeBuf I__1354 (
            .O(N__8970),
            .I(N__8964));
    CascadeMux I__1353 (
            .O(N__8967),
            .I(N__8961));
    CascadeMux I__1352 (
            .O(N__8964),
            .I(N__8958));
    CascadeBuf I__1351 (
            .O(N__8961),
            .I(N__8955));
    CascadeBuf I__1350 (
            .O(N__8958),
            .I(N__8952));
    CascadeMux I__1349 (
            .O(N__8955),
            .I(N__8949));
    CascadeMux I__1348 (
            .O(N__8952),
            .I(N__8946));
    CascadeBuf I__1347 (
            .O(N__8949),
            .I(N__8943));
    CascadeBuf I__1346 (
            .O(N__8946),
            .I(N__8940));
    CascadeMux I__1345 (
            .O(N__8943),
            .I(N__8937));
    CascadeMux I__1344 (
            .O(N__8940),
            .I(N__8934));
    CascadeBuf I__1343 (
            .O(N__8937),
            .I(N__8931));
    CascadeBuf I__1342 (
            .O(N__8934),
            .I(N__8928));
    CascadeMux I__1341 (
            .O(N__8931),
            .I(N__8925));
    CascadeMux I__1340 (
            .O(N__8928),
            .I(N__8922));
    CascadeBuf I__1339 (
            .O(N__8925),
            .I(N__8919));
    CascadeBuf I__1338 (
            .O(N__8922),
            .I(N__8916));
    CascadeMux I__1337 (
            .O(N__8919),
            .I(N__8913));
    CascadeMux I__1336 (
            .O(N__8916),
            .I(N__8910));
    CascadeBuf I__1335 (
            .O(N__8913),
            .I(N__8907));
    CascadeBuf I__1334 (
            .O(N__8910),
            .I(N__8904));
    CascadeMux I__1333 (
            .O(N__8907),
            .I(N__8901));
    CascadeMux I__1332 (
            .O(N__8904),
            .I(N__8898));
    CascadeBuf I__1331 (
            .O(N__8901),
            .I(N__8895));
    CascadeBuf I__1330 (
            .O(N__8898),
            .I(N__8892));
    CascadeMux I__1329 (
            .O(N__8895),
            .I(N__8889));
    CascadeMux I__1328 (
            .O(N__8892),
            .I(N__8886));
    InMux I__1327 (
            .O(N__8889),
            .I(N__8883));
    CascadeBuf I__1326 (
            .O(N__8886),
            .I(N__8880));
    LocalMux I__1325 (
            .O(N__8883),
            .I(N__8877));
    CascadeMux I__1324 (
            .O(N__8880),
            .I(N__8874));
    Span4Mux_h I__1323 (
            .O(N__8877),
            .I(N__8871));
    InMux I__1322 (
            .O(N__8874),
            .I(N__8868));
    Span4Mux_h I__1321 (
            .O(N__8871),
            .I(N__8865));
    LocalMux I__1320 (
            .O(N__8868),
            .I(N__8862));
    Sp12to4 I__1319 (
            .O(N__8865),
            .I(N__8859));
    Sp12to4 I__1318 (
            .O(N__8862),
            .I(N__8856));
    Span12Mux_s9_v I__1317 (
            .O(N__8859),
            .I(N__8851));
    Span12Mux_s9_v I__1316 (
            .O(N__8856),
            .I(N__8851));
    Odrv12 I__1315 (
            .O(N__8851),
            .I(n26));
    InMux I__1314 (
            .O(N__8848),
            .I(N__8843));
    InMux I__1313 (
            .O(N__8847),
            .I(N__8840));
    InMux I__1312 (
            .O(N__8846),
            .I(N__8837));
    LocalMux I__1311 (
            .O(N__8843),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    LocalMux I__1310 (
            .O(N__8840),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    LocalMux I__1309 (
            .O(N__8837),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    InMux I__1308 (
            .O(N__8830),
            .I(N__8827));
    LocalMux I__1307 (
            .O(N__8827),
            .I(\receive_module.rx_counter.n10_adj_570 ));
    CascadeMux I__1306 (
            .O(N__8824),
            .I(N__8821));
    InMux I__1305 (
            .O(N__8821),
            .I(N__8816));
    InMux I__1304 (
            .O(N__8820),
            .I(N__8813));
    InMux I__1303 (
            .O(N__8819),
            .I(N__8810));
    LocalMux I__1302 (
            .O(N__8816),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    LocalMux I__1301 (
            .O(N__8813),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    LocalMux I__1300 (
            .O(N__8810),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    IoInMux I__1299 (
            .O(N__8803),
            .I(N__8800));
    LocalMux I__1298 (
            .O(N__8800),
            .I(N__8797));
    IoSpan4Mux I__1297 (
            .O(N__8797),
            .I(N__8794));
    Sp12to4 I__1296 (
            .O(N__8794),
            .I(N__8791));
    Span12Mux_s9_v I__1295 (
            .O(N__8791),
            .I(N__8787));
    InMux I__1294 (
            .O(N__8790),
            .I(N__8784));
    Odrv12 I__1293 (
            .O(N__8787),
            .I(LED_c));
    LocalMux I__1292 (
            .O(N__8784),
            .I(LED_c));
    InMux I__1291 (
            .O(N__8779),
            .I(\transmit_module.n2743 ));
    InMux I__1290 (
            .O(N__8776),
            .I(\transmit_module.n2744 ));
    InMux I__1289 (
            .O(N__8773),
            .I(\transmit_module.n2745 ));
    InMux I__1288 (
            .O(N__8770),
            .I(\transmit_module.n2746 ));
    InMux I__1287 (
            .O(N__8767),
            .I(bfn_15_18_0_));
    InMux I__1286 (
            .O(N__8764),
            .I(\transmit_module.n2748 ));
    InMux I__1285 (
            .O(N__8761),
            .I(\transmit_module.n2749 ));
    InMux I__1284 (
            .O(N__8758),
            .I(\transmit_module.n2750 ));
    InMux I__1283 (
            .O(N__8755),
            .I(\transmit_module.n2751 ));
    InMux I__1282 (
            .O(N__8752),
            .I(N__8747));
    InMux I__1281 (
            .O(N__8751),
            .I(N__8744));
    InMux I__1280 (
            .O(N__8750),
            .I(N__8741));
    LocalMux I__1279 (
            .O(N__8747),
            .I(N__8738));
    LocalMux I__1278 (
            .O(N__8744),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__1277 (
            .O(N__8741),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    Odrv4 I__1276 (
            .O(N__8738),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    InMux I__1275 (
            .O(N__8731),
            .I(N__8728));
    LocalMux I__1274 (
            .O(N__8728),
            .I(\transmit_module.video_signal_controller.n3183 ));
    CascadeMux I__1273 (
            .O(N__8725),
            .I(N__8721));
    CascadeMux I__1272 (
            .O(N__8724),
            .I(N__8718));
    InMux I__1271 (
            .O(N__8721),
            .I(N__8714));
    InMux I__1270 (
            .O(N__8718),
            .I(N__8711));
    InMux I__1269 (
            .O(N__8717),
            .I(N__8708));
    LocalMux I__1268 (
            .O(N__8714),
            .I(N__8705));
    LocalMux I__1267 (
            .O(N__8711),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    LocalMux I__1266 (
            .O(N__8708),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    Odrv4 I__1265 (
            .O(N__8705),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    InMux I__1264 (
            .O(N__8698),
            .I(N__8695));
    LocalMux I__1263 (
            .O(N__8695),
            .I(\transmit_module.video_signal_controller.n6 ));
    CascadeMux I__1262 (
            .O(N__8692),
            .I(N__8688));
    InMux I__1261 (
            .O(N__8691),
            .I(N__8683));
    InMux I__1260 (
            .O(N__8688),
            .I(N__8680));
    InMux I__1259 (
            .O(N__8687),
            .I(N__8677));
    InMux I__1258 (
            .O(N__8686),
            .I(N__8674));
    LocalMux I__1257 (
            .O(N__8683),
            .I(N__8671));
    LocalMux I__1256 (
            .O(N__8680),
            .I(N__8668));
    LocalMux I__1255 (
            .O(N__8677),
            .I(N__8665));
    LocalMux I__1254 (
            .O(N__8674),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__1253 (
            .O(N__8671),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__1252 (
            .O(N__8668),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__1251 (
            .O(N__8665),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    InMux I__1250 (
            .O(N__8656),
            .I(N__8650));
    InMux I__1249 (
            .O(N__8655),
            .I(N__8647));
    InMux I__1248 (
            .O(N__8654),
            .I(N__8644));
    InMux I__1247 (
            .O(N__8653),
            .I(N__8641));
    LocalMux I__1246 (
            .O(N__8650),
            .I(N__8636));
    LocalMux I__1245 (
            .O(N__8647),
            .I(N__8636));
    LocalMux I__1244 (
            .O(N__8644),
            .I(N__8633));
    LocalMux I__1243 (
            .O(N__8641),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    Odrv4 I__1242 (
            .O(N__8636),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    Odrv4 I__1241 (
            .O(N__8633),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    CascadeMux I__1240 (
            .O(N__8626),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_558_cascade_ ));
    InMux I__1239 (
            .O(N__8623),
            .I(N__8620));
    LocalMux I__1238 (
            .O(N__8620),
            .I(\transmit_module.video_signal_controller.n18 ));
    CascadeMux I__1237 (
            .O(N__8617),
            .I(VGA_VISIBLE_cascade_));
    CascadeMux I__1236 (
            .O(N__8614),
            .I(N__8610));
    InMux I__1235 (
            .O(N__8613),
            .I(N__8607));
    InMux I__1234 (
            .O(N__8610),
            .I(N__8604));
    LocalMux I__1233 (
            .O(N__8607),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    LocalMux I__1232 (
            .O(N__8604),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    InMux I__1231 (
            .O(N__8599),
            .I(\transmit_module.n2740 ));
    InMux I__1230 (
            .O(N__8596),
            .I(\transmit_module.n2741 ));
    InMux I__1229 (
            .O(N__8593),
            .I(\transmit_module.n2742 ));
    InMux I__1228 (
            .O(N__8590),
            .I(bfn_15_11_0_));
    CascadeMux I__1227 (
            .O(N__8587),
            .I(N__8583));
    InMux I__1226 (
            .O(N__8586),
            .I(N__8580));
    InMux I__1225 (
            .O(N__8583),
            .I(N__8577));
    LocalMux I__1224 (
            .O(N__8580),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    LocalMux I__1223 (
            .O(N__8577),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    InMux I__1222 (
            .O(N__8572),
            .I(\receive_module.rx_counter.n2753 ));
    InMux I__1221 (
            .O(N__8569),
            .I(N__8565));
    InMux I__1220 (
            .O(N__8568),
            .I(N__8562));
    LocalMux I__1219 (
            .O(N__8565),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    LocalMux I__1218 (
            .O(N__8562),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    InMux I__1217 (
            .O(N__8557),
            .I(\receive_module.rx_counter.n2754 ));
    InMux I__1216 (
            .O(N__8554),
            .I(N__8550));
    InMux I__1215 (
            .O(N__8553),
            .I(N__8547));
    LocalMux I__1214 (
            .O(N__8550),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    LocalMux I__1213 (
            .O(N__8547),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    InMux I__1212 (
            .O(N__8542),
            .I(\receive_module.rx_counter.n2755 ));
    InMux I__1211 (
            .O(N__8539),
            .I(N__8535));
    InMux I__1210 (
            .O(N__8538),
            .I(N__8532));
    LocalMux I__1209 (
            .O(N__8535),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    LocalMux I__1208 (
            .O(N__8532),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    InMux I__1207 (
            .O(N__8527),
            .I(\receive_module.rx_counter.n2756 ));
    InMux I__1206 (
            .O(N__8524),
            .I(\receive_module.rx_counter.n2757 ));
    SRMux I__1205 (
            .O(N__8521),
            .I(N__8518));
    LocalMux I__1204 (
            .O(N__8518),
            .I(N__8515));
    Span4Mux_h I__1203 (
            .O(N__8515),
            .I(N__8512));
    Odrv4 I__1202 (
            .O(N__8512),
            .I(\receive_module.rx_counter.n2227 ));
    IoInMux I__1201 (
            .O(N__8509),
            .I(N__8506));
    LocalMux I__1200 (
            .O(N__8506),
            .I(N__8503));
    IoSpan4Mux I__1199 (
            .O(N__8503),
            .I(N__8499));
    IoInMux I__1198 (
            .O(N__8502),
            .I(N__8495));
    Span4Mux_s2_v I__1197 (
            .O(N__8499),
            .I(N__8492));
    IoInMux I__1196 (
            .O(N__8498),
            .I(N__8489));
    LocalMux I__1195 (
            .O(N__8495),
            .I(N__8486));
    Span4Mux_v I__1194 (
            .O(N__8492),
            .I(N__8483));
    LocalMux I__1193 (
            .O(N__8489),
            .I(N__8480));
    Span4Mux_s2_v I__1192 (
            .O(N__8486),
            .I(N__8477));
    Sp12to4 I__1191 (
            .O(N__8483),
            .I(N__8472));
    Span12Mux_s2_h I__1190 (
            .O(N__8480),
            .I(N__8472));
    Span4Mux_h I__1189 (
            .O(N__8477),
            .I(N__8469));
    Span12Mux_v I__1188 (
            .O(N__8472),
            .I(N__8466));
    Sp12to4 I__1187 (
            .O(N__8469),
            .I(N__8463));
    Span12Mux_h I__1186 (
            .O(N__8466),
            .I(N__8460));
    Span12Mux_s9_v I__1185 (
            .O(N__8463),
            .I(N__8457));
    Odrv12 I__1184 (
            .O(N__8460),
            .I(n1955));
    Odrv12 I__1183 (
            .O(N__8457),
            .I(n1955));
    InMux I__1182 (
            .O(N__8452),
            .I(N__8449));
    LocalMux I__1181 (
            .O(N__8449),
            .I(N__8446));
    Span4Mux_h I__1180 (
            .O(N__8446),
            .I(N__8443));
    Odrv4 I__1179 (
            .O(N__8443),
            .I(TX_DATA_2));
    IoInMux I__1178 (
            .O(N__8440),
            .I(N__8437));
    LocalMux I__1177 (
            .O(N__8437),
            .I(N__8434));
    IoSpan4Mux I__1176 (
            .O(N__8434),
            .I(N__8430));
    IoInMux I__1175 (
            .O(N__8433),
            .I(N__8426));
    IoSpan4Mux I__1174 (
            .O(N__8430),
            .I(N__8423));
    IoInMux I__1173 (
            .O(N__8429),
            .I(N__8420));
    LocalMux I__1172 (
            .O(N__8426),
            .I(N__8417));
    Span4Mux_s3_v I__1171 (
            .O(N__8423),
            .I(N__8414));
    LocalMux I__1170 (
            .O(N__8420),
            .I(N__8411));
    Span12Mux_s5_v I__1169 (
            .O(N__8417),
            .I(N__8408));
    Sp12to4 I__1168 (
            .O(N__8414),
            .I(N__8405));
    Span12Mux_s2_h I__1167 (
            .O(N__8411),
            .I(N__8402));
    Span12Mux_v I__1166 (
            .O(N__8408),
            .I(N__8399));
    Span12Mux_s10_v I__1165 (
            .O(N__8405),
            .I(N__8394));
    Span12Mux_h I__1164 (
            .O(N__8402),
            .I(N__8394));
    Odrv12 I__1163 (
            .O(N__8399),
            .I(n1953));
    Odrv12 I__1162 (
            .O(N__8394),
            .I(n1953));
    CascadeMux I__1161 (
            .O(N__8389),
            .I(\line_buffer.n3031_cascade_ ));
    InMux I__1160 (
            .O(N__8386),
            .I(N__8383));
    LocalMux I__1159 (
            .O(N__8383),
            .I(N__8380));
    Odrv12 I__1158 (
            .O(N__8380),
            .I(\line_buffer.n3030 ));
    CascadeMux I__1157 (
            .O(N__8377),
            .I(\line_buffer.n3095_cascade_ ));
    InMux I__1156 (
            .O(N__8374),
            .I(N__8371));
    LocalMux I__1155 (
            .O(N__8371),
            .I(N__8368));
    Span4Mux_h I__1154 (
            .O(N__8368),
            .I(N__8365));
    Odrv4 I__1153 (
            .O(N__8365),
            .I(\line_buffer.n3040 ));
    InMux I__1152 (
            .O(N__8362),
            .I(N__8359));
    LocalMux I__1151 (
            .O(N__8359),
            .I(N__8356));
    Span4Mux_v I__1150 (
            .O(N__8356),
            .I(N__8353));
    Span4Mux_h I__1149 (
            .O(N__8353),
            .I(N__8350));
    Span4Mux_h I__1148 (
            .O(N__8350),
            .I(N__8347));
    Odrv4 I__1147 (
            .O(N__8347),
            .I(\line_buffer.n625 ));
    InMux I__1146 (
            .O(N__8344),
            .I(N__8341));
    LocalMux I__1145 (
            .O(N__8341),
            .I(N__8338));
    Span4Mux_v I__1144 (
            .O(N__8338),
            .I(N__8335));
    Sp12to4 I__1143 (
            .O(N__8335),
            .I(N__8332));
    Span12Mux_h I__1142 (
            .O(N__8332),
            .I(N__8329));
    Span12Mux_v I__1141 (
            .O(N__8329),
            .I(N__8326));
    Odrv12 I__1140 (
            .O(N__8326),
            .I(\line_buffer.n617 ));
    InMux I__1139 (
            .O(N__8323),
            .I(N__8320));
    LocalMux I__1138 (
            .O(N__8320),
            .I(N__8317));
    Odrv12 I__1137 (
            .O(N__8317),
            .I(\line_buffer.n3089 ));
    CascadeMux I__1136 (
            .O(N__8314),
            .I(\line_buffer.n3092_cascade_ ));
    InMux I__1135 (
            .O(N__8311),
            .I(N__8308));
    LocalMux I__1134 (
            .O(N__8308),
            .I(\line_buffer.n3146 ));
    InMux I__1133 (
            .O(N__8305),
            .I(N__8302));
    LocalMux I__1132 (
            .O(N__8302),
            .I(N__8299));
    Span12Mux_h I__1131 (
            .O(N__8299),
            .I(N__8296));
    Odrv12 I__1130 (
            .O(N__8296),
            .I(\line_buffer.n626 ));
    InMux I__1129 (
            .O(N__8293),
            .I(N__8290));
    LocalMux I__1128 (
            .O(N__8290),
            .I(N__8287));
    Span4Mux_h I__1127 (
            .O(N__8287),
            .I(N__8284));
    Span4Mux_h I__1126 (
            .O(N__8284),
            .I(N__8281));
    Sp12to4 I__1125 (
            .O(N__8281),
            .I(N__8278));
    Odrv12 I__1124 (
            .O(N__8278),
            .I(\line_buffer.n618 ));
    InMux I__1123 (
            .O(N__8275),
            .I(N__8272));
    LocalMux I__1122 (
            .O(N__8272),
            .I(N__8269));
    Odrv12 I__1121 (
            .O(N__8269),
            .I(\line_buffer.n3039 ));
    CascadeMux I__1120 (
            .O(N__8266),
            .I(\receive_module.rx_counter.n10_adj_570_cascade_ ));
    InMux I__1119 (
            .O(N__8263),
            .I(N__8258));
    InMux I__1118 (
            .O(N__8262),
            .I(N__8255));
    InMux I__1117 (
            .O(N__8261),
            .I(N__8252));
    LocalMux I__1116 (
            .O(N__8258),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__1115 (
            .O(N__8255),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__1114 (
            .O(N__8252),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    InMux I__1113 (
            .O(N__8245),
            .I(N__8240));
    InMux I__1112 (
            .O(N__8244),
            .I(N__8235));
    InMux I__1111 (
            .O(N__8243),
            .I(N__8235));
    LocalMux I__1110 (
            .O(N__8240),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__1109 (
            .O(N__8235),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    InMux I__1108 (
            .O(N__8230),
            .I(N__8227));
    LocalMux I__1107 (
            .O(N__8227),
            .I(\transmit_module.X_DELTA_PATTERN_1 ));
    InMux I__1106 (
            .O(N__8224),
            .I(N__8221));
    LocalMux I__1105 (
            .O(N__8221),
            .I(\transmit_module.X_DELTA_PATTERN_2 ));
    InMux I__1104 (
            .O(N__8218),
            .I(N__8215));
    LocalMux I__1103 (
            .O(N__8215),
            .I(\transmit_module.X_DELTA_PATTERN_6 ));
    InMux I__1102 (
            .O(N__8212),
            .I(N__8209));
    LocalMux I__1101 (
            .O(N__8209),
            .I(\transmit_module.X_DELTA_PATTERN_5 ));
    InMux I__1100 (
            .O(N__8206),
            .I(N__8203));
    LocalMux I__1099 (
            .O(N__8203),
            .I(\transmit_module.X_DELTA_PATTERN_4 ));
    InMux I__1098 (
            .O(N__8200),
            .I(N__8197));
    LocalMux I__1097 (
            .O(N__8197),
            .I(\transmit_module.X_DELTA_PATTERN_3 ));
    InMux I__1096 (
            .O(N__8194),
            .I(N__8191));
    LocalMux I__1095 (
            .O(N__8191),
            .I(N__8188));
    Odrv12 I__1094 (
            .O(N__8188),
            .I(\line_buffer.n755 ));
    InMux I__1093 (
            .O(N__8185),
            .I(N__8182));
    LocalMux I__1092 (
            .O(N__8182),
            .I(N__8179));
    Span12Mux_h I__1091 (
            .O(N__8179),
            .I(N__8176));
    Span12Mux_v I__1090 (
            .O(N__8176),
            .I(N__8173));
    Odrv12 I__1089 (
            .O(N__8173),
            .I(\line_buffer.n747 ));
    InMux I__1088 (
            .O(N__8170),
            .I(\transmit_module.video_signal_controller.n2778 ));
    InMux I__1087 (
            .O(N__8167),
            .I(\transmit_module.video_signal_controller.n2779 ));
    InMux I__1086 (
            .O(N__8164),
            .I(\transmit_module.video_signal_controller.n2780 ));
    InMux I__1085 (
            .O(N__8161),
            .I(\transmit_module.video_signal_controller.n2781 ));
    SRMux I__1084 (
            .O(N__8158),
            .I(N__8154));
    SRMux I__1083 (
            .O(N__8157),
            .I(N__8150));
    LocalMux I__1082 (
            .O(N__8154),
            .I(N__8147));
    CEMux I__1081 (
            .O(N__8153),
            .I(N__8144));
    LocalMux I__1080 (
            .O(N__8150),
            .I(N__8141));
    Span4Mux_h I__1079 (
            .O(N__8147),
            .I(N__8138));
    LocalMux I__1078 (
            .O(N__8144),
            .I(n2147));
    Odrv4 I__1077 (
            .O(N__8141),
            .I(n2147));
    Odrv4 I__1076 (
            .O(N__8138),
            .I(n2147));
    SRMux I__1075 (
            .O(N__8131),
            .I(N__8128));
    LocalMux I__1074 (
            .O(N__8128),
            .I(\transmit_module.video_signal_controller.n2262 ));
    InMux I__1073 (
            .O(N__8125),
            .I(N__8121));
    InMux I__1072 (
            .O(N__8124),
            .I(N__8118));
    LocalMux I__1071 (
            .O(N__8121),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    LocalMux I__1070 (
            .O(N__8118),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    CascadeMux I__1069 (
            .O(N__8113),
            .I(\transmit_module.video_signal_controller.n3022_cascade_ ));
    InMux I__1068 (
            .O(N__8110),
            .I(N__8105));
    InMux I__1067 (
            .O(N__8109),
            .I(N__8102));
    InMux I__1066 (
            .O(N__8108),
            .I(N__8098));
    LocalMux I__1065 (
            .O(N__8105),
            .I(N__8093));
    LocalMux I__1064 (
            .O(N__8102),
            .I(N__8093));
    InMux I__1063 (
            .O(N__8101),
            .I(N__8090));
    LocalMux I__1062 (
            .O(N__8098),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    Odrv4 I__1061 (
            .O(N__8093),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    LocalMux I__1060 (
            .O(N__8090),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    InMux I__1059 (
            .O(N__8083),
            .I(N__8076));
    InMux I__1058 (
            .O(N__8082),
            .I(N__8073));
    InMux I__1057 (
            .O(N__8081),
            .I(N__8068));
    InMux I__1056 (
            .O(N__8080),
            .I(N__8068));
    InMux I__1055 (
            .O(N__8079),
            .I(N__8065));
    LocalMux I__1054 (
            .O(N__8076),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1053 (
            .O(N__8073),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1052 (
            .O(N__8068),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1051 (
            .O(N__8065),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    CascadeMux I__1050 (
            .O(N__8056),
            .I(N__8053));
    InMux I__1049 (
            .O(N__8053),
            .I(N__8046));
    InMux I__1048 (
            .O(N__8052),
            .I(N__8043));
    InMux I__1047 (
            .O(N__8051),
            .I(N__8036));
    InMux I__1046 (
            .O(N__8050),
            .I(N__8036));
    InMux I__1045 (
            .O(N__8049),
            .I(N__8036));
    LocalMux I__1044 (
            .O(N__8046),
            .I(N__8033));
    LocalMux I__1043 (
            .O(N__8043),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__1042 (
            .O(N__8036),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    Odrv4 I__1041 (
            .O(N__8033),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    InMux I__1040 (
            .O(N__8026),
            .I(N__8019));
    InMux I__1039 (
            .O(N__8025),
            .I(N__8016));
    InMux I__1038 (
            .O(N__8024),
            .I(N__8011));
    InMux I__1037 (
            .O(N__8023),
            .I(N__8011));
    InMux I__1036 (
            .O(N__8022),
            .I(N__8008));
    LocalMux I__1035 (
            .O(N__8019),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1034 (
            .O(N__8016),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1033 (
            .O(N__8011),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1032 (
            .O(N__8008),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    InMux I__1031 (
            .O(N__7999),
            .I(N__7994));
    InMux I__1030 (
            .O(N__7998),
            .I(N__7989));
    InMux I__1029 (
            .O(N__7997),
            .I(N__7989));
    LocalMux I__1028 (
            .O(N__7994),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1027 (
            .O(N__7989),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    InMux I__1026 (
            .O(N__7984),
            .I(N__7979));
    InMux I__1025 (
            .O(N__7983),
            .I(N__7976));
    InMux I__1024 (
            .O(N__7982),
            .I(N__7973));
    LocalMux I__1023 (
            .O(N__7979),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1022 (
            .O(N__7976),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1021 (
            .O(N__7973),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    InMux I__1020 (
            .O(N__7966),
            .I(N__7963));
    LocalMux I__1019 (
            .O(N__7963),
            .I(\transmit_module.X_DELTA_PATTERN_15 ));
    InMux I__1018 (
            .O(N__7960),
            .I(N__7957));
    LocalMux I__1017 (
            .O(N__7957),
            .I(\transmit_module.X_DELTA_PATTERN_14 ));
    InMux I__1016 (
            .O(N__7954),
            .I(N__7951));
    LocalMux I__1015 (
            .O(N__7951),
            .I(N__7948));
    Odrv12 I__1014 (
            .O(N__7948),
            .I(\line_buffer.n754 ));
    InMux I__1013 (
            .O(N__7945),
            .I(N__7942));
    LocalMux I__1012 (
            .O(N__7942),
            .I(N__7939));
    Span12Mux_h I__1011 (
            .O(N__7939),
            .I(N__7936));
    Span12Mux_v I__1010 (
            .O(N__7936),
            .I(N__7933));
    Odrv12 I__1009 (
            .O(N__7933),
            .I(\line_buffer.n746 ));
    InMux I__1008 (
            .O(N__7930),
            .I(N__7927));
    LocalMux I__1007 (
            .O(N__7927),
            .I(N__7924));
    Span12Mux_v I__1006 (
            .O(N__7924),
            .I(N__7921));
    Span12Mux_h I__1005 (
            .O(N__7921),
            .I(N__7918));
    Odrv12 I__1004 (
            .O(N__7918),
            .I(\line_buffer.n682 ));
    CascadeMux I__1003 (
            .O(N__7915),
            .I(\line_buffer.n3143_cascade_ ));
    InMux I__1002 (
            .O(N__7912),
            .I(N__7909));
    LocalMux I__1001 (
            .O(N__7909),
            .I(N__7906));
    Span4Mux_v I__1000 (
            .O(N__7906),
            .I(N__7903));
    Span4Mux_h I__999 (
            .O(N__7903),
            .I(N__7900));
    Span4Mux_v I__998 (
            .O(N__7900),
            .I(N__7897));
    Span4Mux_v I__997 (
            .O(N__7897),
            .I(N__7894));
    Odrv4 I__996 (
            .O(N__7894),
            .I(\line_buffer.n690 ));
    InMux I__995 (
            .O(N__7891),
            .I(N__7888));
    LocalMux I__994 (
            .O(N__7888),
            .I(N__7885));
    Span4Mux_h I__993 (
            .O(N__7885),
            .I(N__7882));
    Span4Mux_h I__992 (
            .O(N__7882),
            .I(N__7879));
    Odrv4 I__991 (
            .O(N__7879),
            .I(\line_buffer.n694 ));
    CascadeMux I__990 (
            .O(N__7876),
            .I(N__7873));
    InMux I__989 (
            .O(N__7873),
            .I(N__7870));
    LocalMux I__988 (
            .O(N__7870),
            .I(N__7867));
    Span12Mux_v I__987 (
            .O(N__7867),
            .I(N__7864));
    Span12Mux_v I__986 (
            .O(N__7864),
            .I(N__7861));
    Span12Mux_h I__985 (
            .O(N__7861),
            .I(N__7858));
    Odrv12 I__984 (
            .O(N__7858),
            .I(\line_buffer.n686 ));
    InMux I__983 (
            .O(N__7855),
            .I(N__7852));
    LocalMux I__982 (
            .O(N__7852),
            .I(\line_buffer.n3101 ));
    InMux I__981 (
            .O(N__7849),
            .I(N__7846));
    LocalMux I__980 (
            .O(N__7846),
            .I(N__7843));
    Span4Mux_h I__979 (
            .O(N__7843),
            .I(N__7840));
    Span4Mux_h I__978 (
            .O(N__7840),
            .I(N__7837));
    Span4Mux_v I__977 (
            .O(N__7837),
            .I(N__7834));
    Odrv4 I__976 (
            .O(N__7834),
            .I(\line_buffer.n691 ));
    InMux I__975 (
            .O(N__7831),
            .I(N__7828));
    LocalMux I__974 (
            .O(N__7828),
            .I(N__7825));
    Span12Mux_h I__973 (
            .O(N__7825),
            .I(N__7822));
    Odrv12 I__972 (
            .O(N__7822),
            .I(\line_buffer.n683 ));
    InMux I__971 (
            .O(N__7819),
            .I(N__7816));
    LocalMux I__970 (
            .O(N__7816),
            .I(N__7813));
    Span4Mux_h I__969 (
            .O(N__7813),
            .I(N__7810));
    Span4Mux_h I__968 (
            .O(N__7810),
            .I(N__7807));
    Odrv4 I__967 (
            .O(N__7807),
            .I(\line_buffer.n722 ));
    InMux I__966 (
            .O(N__7804),
            .I(N__7801));
    LocalMux I__965 (
            .O(N__7801),
            .I(N__7798));
    Span4Mux_v I__964 (
            .O(N__7798),
            .I(N__7795));
    Span4Mux_h I__963 (
            .O(N__7795),
            .I(N__7792));
    Span4Mux_h I__962 (
            .O(N__7792),
            .I(N__7789));
    Odrv4 I__961 (
            .O(N__7789),
            .I(\line_buffer.n714 ));
    InMux I__960 (
            .O(N__7786),
            .I(bfn_14_14_0_));
    InMux I__959 (
            .O(N__7783),
            .I(\transmit_module.video_signal_controller.n2776 ));
    InMux I__958 (
            .O(N__7780),
            .I(\transmit_module.video_signal_controller.n2777 ));
    InMux I__957 (
            .O(N__7777),
            .I(bfn_13_16_0_));
    InMux I__956 (
            .O(N__7774),
            .I(\transmit_module.video_signal_controller.n2774 ));
    InMux I__955 (
            .O(N__7771),
            .I(\transmit_module.video_signal_controller.n2775 ));
    InMux I__954 (
            .O(N__7768),
            .I(N__7765));
    LocalMux I__953 (
            .O(N__7765),
            .I(\transmit_module.X_DELTA_PATTERN_13 ));
    InMux I__952 (
            .O(N__7762),
            .I(N__7759));
    LocalMux I__951 (
            .O(N__7759),
            .I(\transmit_module.X_DELTA_PATTERN_10 ));
    InMux I__950 (
            .O(N__7756),
            .I(N__7753));
    LocalMux I__949 (
            .O(N__7753),
            .I(\transmit_module.X_DELTA_PATTERN_12 ));
    InMux I__948 (
            .O(N__7750),
            .I(N__7747));
    LocalMux I__947 (
            .O(N__7747),
            .I(\transmit_module.X_DELTA_PATTERN_11 ));
    InMux I__946 (
            .O(N__7744),
            .I(N__7741));
    LocalMux I__945 (
            .O(N__7741),
            .I(\transmit_module.X_DELTA_PATTERN_7 ));
    InMux I__944 (
            .O(N__7738),
            .I(N__7734));
    CascadeMux I__943 (
            .O(N__7737),
            .I(N__7729));
    LocalMux I__942 (
            .O(N__7734),
            .I(N__7726));
    InMux I__941 (
            .O(N__7733),
            .I(N__7723));
    InMux I__940 (
            .O(N__7732),
            .I(N__7720));
    InMux I__939 (
            .O(N__7729),
            .I(N__7717));
    Odrv4 I__938 (
            .O(N__7726),
            .I(Y_0));
    LocalMux I__937 (
            .O(N__7723),
            .I(Y_0));
    LocalMux I__936 (
            .O(N__7720),
            .I(Y_0));
    LocalMux I__935 (
            .O(N__7717),
            .I(Y_0));
    InMux I__934 (
            .O(N__7708),
            .I(N__7705));
    LocalMux I__933 (
            .O(N__7705),
            .I(N__7699));
    InMux I__932 (
            .O(N__7704),
            .I(N__7696));
    InMux I__931 (
            .O(N__7703),
            .I(N__7693));
    InMux I__930 (
            .O(N__7702),
            .I(N__7690));
    Odrv4 I__929 (
            .O(N__7699),
            .I(Y_1));
    LocalMux I__928 (
            .O(N__7696),
            .I(Y_1));
    LocalMux I__927 (
            .O(N__7693),
            .I(Y_1));
    LocalMux I__926 (
            .O(N__7690),
            .I(Y_1));
    CascadeMux I__925 (
            .O(N__7681),
            .I(n5_cascade_));
    InMux I__924 (
            .O(N__7678),
            .I(N__7675));
    LocalMux I__923 (
            .O(N__7675),
            .I(n3009));
    InMux I__922 (
            .O(N__7672),
            .I(N__7668));
    InMux I__921 (
            .O(N__7671),
            .I(N__7665));
    LocalMux I__920 (
            .O(N__7668),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    LocalMux I__919 (
            .O(N__7665),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    InMux I__918 (
            .O(N__7660),
            .I(bfn_13_15_0_));
    InMux I__917 (
            .O(N__7657),
            .I(N__7653));
    InMux I__916 (
            .O(N__7656),
            .I(N__7650));
    LocalMux I__915 (
            .O(N__7653),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__914 (
            .O(N__7650),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    InMux I__913 (
            .O(N__7645),
            .I(\transmit_module.video_signal_controller.n2766 ));
    InMux I__912 (
            .O(N__7642),
            .I(N__7638));
    InMux I__911 (
            .O(N__7641),
            .I(N__7635));
    LocalMux I__910 (
            .O(N__7638),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__909 (
            .O(N__7635),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    InMux I__908 (
            .O(N__7630),
            .I(\transmit_module.video_signal_controller.n2767 ));
    InMux I__907 (
            .O(N__7627),
            .I(N__7622));
    InMux I__906 (
            .O(N__7626),
            .I(N__7619));
    InMux I__905 (
            .O(N__7625),
            .I(N__7616));
    LocalMux I__904 (
            .O(N__7622),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__903 (
            .O(N__7619),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__902 (
            .O(N__7616),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    InMux I__901 (
            .O(N__7609),
            .I(\transmit_module.video_signal_controller.n2768 ));
    InMux I__900 (
            .O(N__7606),
            .I(N__7600));
    InMux I__899 (
            .O(N__7605),
            .I(N__7593));
    InMux I__898 (
            .O(N__7604),
            .I(N__7593));
    InMux I__897 (
            .O(N__7603),
            .I(N__7593));
    LocalMux I__896 (
            .O(N__7600),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__895 (
            .O(N__7593),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    InMux I__894 (
            .O(N__7588),
            .I(\transmit_module.video_signal_controller.n2769 ));
    InMux I__893 (
            .O(N__7585),
            .I(\transmit_module.video_signal_controller.n2770 ));
    InMux I__892 (
            .O(N__7582),
            .I(\transmit_module.video_signal_controller.n2771 ));
    InMux I__891 (
            .O(N__7579),
            .I(\transmit_module.video_signal_controller.n2772 ));
    InMux I__890 (
            .O(N__7576),
            .I(N__7573));
    LocalMux I__889 (
            .O(N__7573),
            .I(\transmit_module.X_DELTA_PATTERN_9 ));
    InMux I__888 (
            .O(N__7570),
            .I(N__7567));
    LocalMux I__887 (
            .O(N__7567),
            .I(\transmit_module.X_DELTA_PATTERN_8 ));
    InMux I__886 (
            .O(N__7564),
            .I(N__7561));
    LocalMux I__885 (
            .O(N__7561),
            .I(N__7558));
    Span12Mux_v I__884 (
            .O(N__7558),
            .I(N__7555));
    Odrv12 I__883 (
            .O(N__7555),
            .I(\line_buffer.n758 ));
    InMux I__882 (
            .O(N__7552),
            .I(N__7549));
    LocalMux I__881 (
            .O(N__7549),
            .I(N__7546));
    Span4Mux_v I__880 (
            .O(N__7546),
            .I(N__7543));
    Odrv4 I__879 (
            .O(N__7543),
            .I(\line_buffer.n750 ));
    CEMux I__878 (
            .O(N__7540),
            .I(N__7536));
    CEMux I__877 (
            .O(N__7539),
            .I(N__7533));
    LocalMux I__876 (
            .O(N__7536),
            .I(\receive_module.n2152 ));
    LocalMux I__875 (
            .O(N__7533),
            .I(\receive_module.n2152 ));
    InMux I__874 (
            .O(N__7528),
            .I(N__7525));
    LocalMux I__873 (
            .O(N__7525),
            .I(N__7520));
    InMux I__872 (
            .O(N__7524),
            .I(N__7515));
    InMux I__871 (
            .O(N__7523),
            .I(N__7515));
    Span4Mux_v I__870 (
            .O(N__7520),
            .I(N__7512));
    LocalMux I__869 (
            .O(N__7515),
            .I(N__7509));
    Span4Mux_h I__868 (
            .O(N__7512),
            .I(N__7506));
    Span4Mux_v I__867 (
            .O(N__7509),
            .I(N__7503));
    Span4Mux_h I__866 (
            .O(N__7506),
            .I(N__7500));
    Sp12to4 I__865 (
            .O(N__7503),
            .I(N__7497));
    Sp12to4 I__864 (
            .O(N__7500),
            .I(N__7492));
    Span12Mux_h I__863 (
            .O(N__7497),
            .I(N__7492));
    Odrv12 I__862 (
            .O(N__7492),
            .I(TVP_HSYNC_c));
    InMux I__861 (
            .O(N__7489),
            .I(N__7486));
    LocalMux I__860 (
            .O(N__7486),
            .I(\receive_module.old_HS ));
    InMux I__859 (
            .O(N__7483),
            .I(N__7480));
    LocalMux I__858 (
            .O(N__7480),
            .I(\transmit_module.video_signal_controller.n2484 ));
    InMux I__857 (
            .O(N__7477),
            .I(N__7471));
    InMux I__856 (
            .O(N__7476),
            .I(N__7468));
    InMux I__855 (
            .O(N__7475),
            .I(N__7463));
    InMux I__854 (
            .O(N__7474),
            .I(N__7463));
    LocalMux I__853 (
            .O(N__7471),
            .I(N__7460));
    LocalMux I__852 (
            .O(N__7468),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__851 (
            .O(N__7463),
            .I(\receive_module.rx_counter.Y_5 ));
    Odrv4 I__850 (
            .O(N__7460),
            .I(\receive_module.rx_counter.Y_5 ));
    CascadeMux I__849 (
            .O(N__7453),
            .I(n2147_cascade_));
    InMux I__848 (
            .O(N__7450),
            .I(N__7444));
    InMux I__847 (
            .O(N__7449),
            .I(N__7441));
    InMux I__846 (
            .O(N__7448),
            .I(N__7436));
    InMux I__845 (
            .O(N__7447),
            .I(N__7436));
    LocalMux I__844 (
            .O(N__7444),
            .I(N__7433));
    LocalMux I__843 (
            .O(N__7441),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__842 (
            .O(N__7436),
            .I(\receive_module.rx_counter.Y_6 ));
    Odrv4 I__841 (
            .O(N__7433),
            .I(\receive_module.rx_counter.Y_6 ));
    InMux I__840 (
            .O(N__7426),
            .I(N__7420));
    InMux I__839 (
            .O(N__7425),
            .I(N__7417));
    InMux I__838 (
            .O(N__7424),
            .I(N__7412));
    InMux I__837 (
            .O(N__7423),
            .I(N__7412));
    LocalMux I__836 (
            .O(N__7420),
            .I(N__7409));
    LocalMux I__835 (
            .O(N__7417),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__834 (
            .O(N__7412),
            .I(\receive_module.rx_counter.Y_2 ));
    Odrv4 I__833 (
            .O(N__7409),
            .I(\receive_module.rx_counter.Y_2 ));
    InMux I__832 (
            .O(N__7402),
            .I(N__7396));
    InMux I__831 (
            .O(N__7401),
            .I(N__7393));
    InMux I__830 (
            .O(N__7400),
            .I(N__7390));
    InMux I__829 (
            .O(N__7399),
            .I(N__7387));
    LocalMux I__828 (
            .O(N__7396),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__827 (
            .O(N__7393),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__826 (
            .O(N__7390),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__825 (
            .O(N__7387),
            .I(\receive_module.rx_counter.Y_8 ));
    CascadeMux I__824 (
            .O(N__7378),
            .I(\receive_module.rx_counter.n6_cascade_ ));
    InMux I__823 (
            .O(N__7375),
            .I(N__7369));
    InMux I__822 (
            .O(N__7374),
            .I(N__7366));
    InMux I__821 (
            .O(N__7373),
            .I(N__7361));
    InMux I__820 (
            .O(N__7372),
            .I(N__7361));
    LocalMux I__819 (
            .O(N__7369),
            .I(N__7358));
    LocalMux I__818 (
            .O(N__7366),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__817 (
            .O(N__7361),
            .I(\receive_module.rx_counter.Y_3 ));
    Odrv4 I__816 (
            .O(N__7358),
            .I(\receive_module.rx_counter.Y_3 ));
    InMux I__815 (
            .O(N__7351),
            .I(N__7348));
    LocalMux I__814 (
            .O(N__7348),
            .I(N__7345));
    Span12Mux_v I__813 (
            .O(N__7345),
            .I(N__7342));
    Odrv12 I__812 (
            .O(N__7342),
            .I(\line_buffer.n723 ));
    InMux I__811 (
            .O(N__7339),
            .I(N__7336));
    LocalMux I__810 (
            .O(N__7336),
            .I(N__7333));
    Span12Mux_h I__809 (
            .O(N__7333),
            .I(N__7330));
    Odrv12 I__808 (
            .O(N__7330),
            .I(\line_buffer.n715 ));
    CascadeMux I__807 (
            .O(N__7327),
            .I(N__7324));
    InMux I__806 (
            .O(N__7324),
            .I(N__7321));
    LocalMux I__805 (
            .O(N__7321),
            .I(\transmit_module.video_signal_controller.n2972 ));
    InMux I__804 (
            .O(N__7318),
            .I(N__7315));
    LocalMux I__803 (
            .O(N__7315),
            .I(\transmit_module.video_signal_controller.n3014 ));
    CascadeMux I__802 (
            .O(N__7312),
            .I(\transmit_module.video_signal_controller.n3186_cascade_ ));
    IoInMux I__801 (
            .O(N__7309),
            .I(N__7306));
    LocalMux I__800 (
            .O(N__7306),
            .I(N__7303));
    Span4Mux_s3_h I__799 (
            .O(N__7303),
            .I(N__7300));
    Sp12to4 I__798 (
            .O(N__7300),
            .I(N__7297));
    Span12Mux_v I__797 (
            .O(N__7297),
            .I(N__7294));
    Odrv12 I__796 (
            .O(N__7294),
            .I(ADV_HSYNC_c));
    InMux I__795 (
            .O(N__7291),
            .I(N__7288));
    LocalMux I__794 (
            .O(N__7288),
            .I(\transmit_module.video_signal_controller.n12 ));
    CascadeMux I__793 (
            .O(N__7285),
            .I(\transmit_module.video_signal_controller.n3182_cascade_ ));
    InMux I__792 (
            .O(N__7282),
            .I(N__7279));
    LocalMux I__791 (
            .O(N__7279),
            .I(\transmit_module.video_signal_controller.n8 ));
    InMux I__790 (
            .O(N__7276),
            .I(\receive_module.rx_counter.n2759 ));
    InMux I__789 (
            .O(N__7273),
            .I(\receive_module.rx_counter.n2760 ));
    InMux I__788 (
            .O(N__7270),
            .I(\receive_module.rx_counter.n2761 ));
    InMux I__787 (
            .O(N__7267),
            .I(\receive_module.rx_counter.n2762 ));
    InMux I__786 (
            .O(N__7264),
            .I(\receive_module.rx_counter.n2763 ));
    InMux I__785 (
            .O(N__7261),
            .I(\receive_module.rx_counter.n2764 ));
    InMux I__784 (
            .O(N__7258),
            .I(bfn_12_13_0_));
    InMux I__783 (
            .O(N__7255),
            .I(N__7252));
    LocalMux I__782 (
            .O(N__7252),
            .I(N__7246));
    InMux I__781 (
            .O(N__7251),
            .I(N__7243));
    InMux I__780 (
            .O(N__7250),
            .I(N__7238));
    InMux I__779 (
            .O(N__7249),
            .I(N__7238));
    Odrv4 I__778 (
            .O(N__7246),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__777 (
            .O(N__7243),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__776 (
            .O(N__7238),
            .I(\receive_module.rx_counter.Y_7 ));
    InMux I__775 (
            .O(N__7231),
            .I(N__7225));
    InMux I__774 (
            .O(N__7230),
            .I(N__7222));
    InMux I__773 (
            .O(N__7229),
            .I(N__7217));
    InMux I__772 (
            .O(N__7228),
            .I(N__7217));
    LocalMux I__771 (
            .O(N__7225),
            .I(N__7214));
    LocalMux I__770 (
            .O(N__7222),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__769 (
            .O(N__7217),
            .I(\receive_module.rx_counter.Y_4 ));
    Odrv4 I__768 (
            .O(N__7214),
            .I(\receive_module.rx_counter.Y_4 ));
    CascadeMux I__767 (
            .O(N__7207),
            .I(\receive_module.rx_counter.n4_cascade_ ));
    CascadeMux I__766 (
            .O(N__7204),
            .I(\receive_module.rx_counter.n2986_cascade_ ));
    CascadeMux I__765 (
            .O(N__7201),
            .I(\receive_module.rx_counter.n2989_cascade_ ));
    InMux I__764 (
            .O(N__7198),
            .I(N__7195));
    LocalMux I__763 (
            .O(N__7195),
            .I(\receive_module.rx_counter.n31_adj_572 ));
    InMux I__762 (
            .O(N__7192),
            .I(N__7189));
    LocalMux I__761 (
            .O(N__7189),
            .I(\receive_module.rx_counter.n7 ));
    InMux I__760 (
            .O(N__7186),
            .I(N__7183));
    LocalMux I__759 (
            .O(N__7183),
            .I(\receive_module.rx_counter.n3166 ));
    CascadeMux I__758 (
            .O(N__7180),
            .I(\receive_module.rx_counter.n2978_cascade_ ));
    InMux I__757 (
            .O(N__7177),
            .I(N__7174));
    LocalMux I__756 (
            .O(N__7174),
            .I(\receive_module.rx_counter.n4_adj_571 ));
    InMux I__755 (
            .O(N__7171),
            .I(bfn_12_12_0_));
    InMux I__754 (
            .O(N__7168),
            .I(\receive_module.rx_counter.n2758 ));
    InMux I__753 (
            .O(N__7165),
            .I(N__7161));
    InMux I__752 (
            .O(N__7164),
            .I(N__7158));
    LocalMux I__751 (
            .O(N__7161),
            .I(\receive_module.rx_counter.X_3 ));
    LocalMux I__750 (
            .O(N__7158),
            .I(\receive_module.rx_counter.X_3 ));
    InMux I__749 (
            .O(N__7153),
            .I(\receive_module.rx_counter.n2784 ));
    InMux I__748 (
            .O(N__7150),
            .I(N__7146));
    InMux I__747 (
            .O(N__7149),
            .I(N__7143));
    LocalMux I__746 (
            .O(N__7146),
            .I(\receive_module.rx_counter.X_4 ));
    LocalMux I__745 (
            .O(N__7143),
            .I(\receive_module.rx_counter.X_4 ));
    InMux I__744 (
            .O(N__7138),
            .I(\receive_module.rx_counter.n2785 ));
    InMux I__743 (
            .O(N__7135),
            .I(N__7131));
    InMux I__742 (
            .O(N__7134),
            .I(N__7128));
    LocalMux I__741 (
            .O(N__7131),
            .I(\receive_module.rx_counter.X_5 ));
    LocalMux I__740 (
            .O(N__7128),
            .I(\receive_module.rx_counter.X_5 ));
    InMux I__739 (
            .O(N__7123),
            .I(\receive_module.rx_counter.n2786 ));
    InMux I__738 (
            .O(N__7120),
            .I(N__7115));
    InMux I__737 (
            .O(N__7119),
            .I(N__7110));
    InMux I__736 (
            .O(N__7118),
            .I(N__7110));
    LocalMux I__735 (
            .O(N__7115),
            .I(\receive_module.rx_counter.X_6 ));
    LocalMux I__734 (
            .O(N__7110),
            .I(\receive_module.rx_counter.X_6 ));
    InMux I__733 (
            .O(N__7105),
            .I(\receive_module.rx_counter.n2787 ));
    InMux I__732 (
            .O(N__7102),
            .I(N__7095));
    InMux I__731 (
            .O(N__7101),
            .I(N__7095));
    InMux I__730 (
            .O(N__7100),
            .I(N__7092));
    LocalMux I__729 (
            .O(N__7095),
            .I(N__7089));
    LocalMux I__728 (
            .O(N__7092),
            .I(\receive_module.rx_counter.X_7 ));
    Odrv4 I__727 (
            .O(N__7089),
            .I(\receive_module.rx_counter.X_7 ));
    InMux I__726 (
            .O(N__7084),
            .I(\receive_module.rx_counter.n2788 ));
    InMux I__725 (
            .O(N__7081),
            .I(N__7077));
    InMux I__724 (
            .O(N__7080),
            .I(N__7074));
    LocalMux I__723 (
            .O(N__7077),
            .I(N__7071));
    LocalMux I__722 (
            .O(N__7074),
            .I(\receive_module.rx_counter.X_8 ));
    Odrv4 I__721 (
            .O(N__7071),
            .I(\receive_module.rx_counter.X_8 ));
    InMux I__720 (
            .O(N__7066),
            .I(bfn_10_15_0_));
    InMux I__719 (
            .O(N__7063),
            .I(\receive_module.rx_counter.n2790 ));
    InMux I__718 (
            .O(N__7060),
            .I(N__7056));
    InMux I__717 (
            .O(N__7059),
            .I(N__7053));
    LocalMux I__716 (
            .O(N__7056),
            .I(N__7050));
    LocalMux I__715 (
            .O(N__7053),
            .I(\receive_module.rx_counter.X_9 ));
    Odrv4 I__714 (
            .O(N__7050),
            .I(\receive_module.rx_counter.X_9 ));
    SRMux I__713 (
            .O(N__7045),
            .I(N__7041));
    SRMux I__712 (
            .O(N__7044),
            .I(N__7038));
    LocalMux I__711 (
            .O(N__7041),
            .I(N__7035));
    LocalMux I__710 (
            .O(N__7038),
            .I(N__7032));
    Sp12to4 I__709 (
            .O(N__7035),
            .I(N__7029));
    Span4Mux_v I__708 (
            .O(N__7032),
            .I(N__7026));
    Odrv12 I__707 (
            .O(N__7029),
            .I(n3184));
    Odrv4 I__706 (
            .O(N__7026),
            .I(n3184));
    InMux I__705 (
            .O(N__7021),
            .I(N__7018));
    LocalMux I__704 (
            .O(N__7018),
            .I(N__7015));
    Span4Mux_v I__703 (
            .O(N__7015),
            .I(N__7012));
    Odrv4 I__702 (
            .O(N__7012),
            .I(\line_buffer.n759 ));
    InMux I__701 (
            .O(N__7009),
            .I(N__7006));
    LocalMux I__700 (
            .O(N__7006),
            .I(N__7003));
    Span4Mux_v I__699 (
            .O(N__7003),
            .I(N__7000));
    Odrv4 I__698 (
            .O(N__7000),
            .I(\line_buffer.n751 ));
    CascadeMux I__697 (
            .O(N__6997),
            .I(\receive_module.rx_counter.n2975_cascade_ ));
    SRMux I__696 (
            .O(N__6994),
            .I(N__6989));
    SRMux I__695 (
            .O(N__6993),
            .I(N__6986));
    SRMux I__694 (
            .O(N__6992),
            .I(N__6982));
    LocalMux I__693 (
            .O(N__6989),
            .I(N__6977));
    LocalMux I__692 (
            .O(N__6986),
            .I(N__6977));
    SRMux I__691 (
            .O(N__6985),
            .I(N__6974));
    LocalMux I__690 (
            .O(N__6982),
            .I(N__6971));
    Span4Mux_v I__689 (
            .O(N__6977),
            .I(N__6966));
    LocalMux I__688 (
            .O(N__6974),
            .I(N__6966));
    Span4Mux_v I__687 (
            .O(N__6971),
            .I(N__6963));
    Span4Mux_v I__686 (
            .O(N__6966),
            .I(N__6960));
    Span4Mux_v I__685 (
            .O(N__6963),
            .I(N__6957));
    Span4Mux_v I__684 (
            .O(N__6960),
            .I(N__6952));
    Span4Mux_v I__683 (
            .O(N__6957),
            .I(N__6952));
    Odrv4 I__682 (
            .O(N__6952),
            .I(\line_buffer.n698 ));
    InMux I__681 (
            .O(N__6949),
            .I(N__6946));
    LocalMux I__680 (
            .O(N__6946),
            .I(\receive_module.rx_counter.n2900 ));
    CascadeMux I__679 (
            .O(N__6943),
            .I(\receive_module.rx_counter.n2900_cascade_ ));
    InMux I__678 (
            .O(N__6940),
            .I(N__6937));
    LocalMux I__677 (
            .O(N__6937),
            .I(\receive_module.rx_counter.n2943 ));
    InMux I__676 (
            .O(N__6934),
            .I(N__6931));
    LocalMux I__675 (
            .O(N__6931),
            .I(\receive_module.rx_counter.n10 ));
    InMux I__674 (
            .O(N__6928),
            .I(bfn_10_14_0_));
    InMux I__673 (
            .O(N__6925),
            .I(N__6922));
    LocalMux I__672 (
            .O(N__6922),
            .I(\receive_module.rx_counter.n9 ));
    InMux I__671 (
            .O(N__6919),
            .I(\receive_module.rx_counter.n2782 ));
    InMux I__670 (
            .O(N__6916),
            .I(N__6913));
    LocalMux I__669 (
            .O(N__6913),
            .I(\receive_module.rx_counter.n8 ));
    InMux I__668 (
            .O(N__6910),
            .I(\receive_module.rx_counter.n2783 ));
    InMux I__667 (
            .O(N__6907),
            .I(N__6904));
    LocalMux I__666 (
            .O(N__6904),
            .I(N__6901));
    Span4Mux_s2_v I__665 (
            .O(N__6901),
            .I(N__6897));
    InMux I__664 (
            .O(N__6900),
            .I(N__6894));
    Span4Mux_v I__663 (
            .O(N__6897),
            .I(N__6889));
    LocalMux I__662 (
            .O(N__6894),
            .I(N__6889));
    Span4Mux_v I__661 (
            .O(N__6889),
            .I(N__6885));
    InMux I__660 (
            .O(N__6888),
            .I(N__6882));
    Span4Mux_v I__659 (
            .O(N__6885),
            .I(N__6876));
    LocalMux I__658 (
            .O(N__6882),
            .I(N__6876));
    InMux I__657 (
            .O(N__6881),
            .I(N__6873));
    Span4Mux_v I__656 (
            .O(N__6876),
            .I(N__6868));
    LocalMux I__655 (
            .O(N__6873),
            .I(N__6868));
    Span4Mux_v I__654 (
            .O(N__6868),
            .I(N__6863));
    InMux I__653 (
            .O(N__6867),
            .I(N__6860));
    InMux I__652 (
            .O(N__6866),
            .I(N__6857));
    Span4Mux_v I__651 (
            .O(N__6863),
            .I(N__6852));
    LocalMux I__650 (
            .O(N__6860),
            .I(N__6852));
    LocalMux I__649 (
            .O(N__6857),
            .I(N__6849));
    Span4Mux_h I__648 (
            .O(N__6852),
            .I(N__6845));
    Span4Mux_h I__647 (
            .O(N__6849),
            .I(N__6842));
    InMux I__646 (
            .O(N__6848),
            .I(N__6839));
    Span4Mux_h I__645 (
            .O(N__6845),
            .I(N__6836));
    Span4Mux_v I__644 (
            .O(N__6842),
            .I(N__6832));
    LocalMux I__643 (
            .O(N__6839),
            .I(N__6829));
    Span4Mux_h I__642 (
            .O(N__6836),
            .I(N__6826));
    InMux I__641 (
            .O(N__6835),
            .I(N__6823));
    Span4Mux_v I__640 (
            .O(N__6832),
            .I(N__6818));
    Span4Mux_h I__639 (
            .O(N__6829),
            .I(N__6818));
    Span4Mux_h I__638 (
            .O(N__6826),
            .I(N__6813));
    LocalMux I__637 (
            .O(N__6823),
            .I(N__6813));
    Span4Mux_v I__636 (
            .O(N__6818),
            .I(N__6810));
    Span4Mux_h I__635 (
            .O(N__6813),
            .I(N__6807));
    Span4Mux_v I__634 (
            .O(N__6810),
            .I(N__6804));
    Span4Mux_v I__633 (
            .O(N__6807),
            .I(N__6801));
    Odrv4 I__632 (
            .O(N__6804),
            .I(TVP_VIDEO_c_2));
    Odrv4 I__631 (
            .O(N__6801),
            .I(TVP_VIDEO_c_2));
    SRMux I__630 (
            .O(N__6796),
            .I(N__6792));
    SRMux I__629 (
            .O(N__6795),
            .I(N__6789));
    LocalMux I__628 (
            .O(N__6792),
            .I(N__6785));
    LocalMux I__627 (
            .O(N__6789),
            .I(N__6782));
    SRMux I__626 (
            .O(N__6788),
            .I(N__6779));
    Span4Mux_v I__625 (
            .O(N__6785),
            .I(N__6776));
    Span4Mux_v I__624 (
            .O(N__6782),
            .I(N__6771));
    LocalMux I__623 (
            .O(N__6779),
            .I(N__6771));
    Span4Mux_v I__622 (
            .O(N__6776),
            .I(N__6768));
    Span4Mux_v I__621 (
            .O(N__6771),
            .I(N__6765));
    Span4Mux_v I__620 (
            .O(N__6768),
            .I(N__6759));
    Span4Mux_h I__619 (
            .O(N__6765),
            .I(N__6759));
    SRMux I__618 (
            .O(N__6764),
            .I(N__6756));
    Odrv4 I__617 (
            .O(N__6759),
            .I(\line_buffer.n730 ));
    LocalMux I__616 (
            .O(N__6756),
            .I(\line_buffer.n730 ));
    SRMux I__615 (
            .O(N__6751),
            .I(N__6748));
    LocalMux I__614 (
            .O(N__6748),
            .I(N__6743));
    SRMux I__613 (
            .O(N__6747),
            .I(N__6740));
    SRMux I__612 (
            .O(N__6746),
            .I(N__6737));
    Span4Mux_v I__611 (
            .O(N__6743),
            .I(N__6733));
    LocalMux I__610 (
            .O(N__6740),
            .I(N__6728));
    LocalMux I__609 (
            .O(N__6737),
            .I(N__6728));
    SRMux I__608 (
            .O(N__6736),
            .I(N__6725));
    Span4Mux_h I__607 (
            .O(N__6733),
            .I(N__6722));
    Span4Mux_v I__606 (
            .O(N__6728),
            .I(N__6717));
    LocalMux I__605 (
            .O(N__6725),
            .I(N__6717));
    Sp12to4 I__604 (
            .O(N__6722),
            .I(N__6714));
    Span4Mux_v I__603 (
            .O(N__6717),
            .I(N__6711));
    Span12Mux_h I__602 (
            .O(N__6714),
            .I(N__6708));
    Span4Mux_v I__601 (
            .O(N__6711),
            .I(N__6705));
    Odrv12 I__600 (
            .O(N__6708),
            .I(\line_buffer.n632 ));
    Odrv4 I__599 (
            .O(N__6705),
            .I(\line_buffer.n632 ));
    SRMux I__598 (
            .O(N__6700),
            .I(N__6697));
    LocalMux I__597 (
            .O(N__6697),
            .I(N__6693));
    SRMux I__596 (
            .O(N__6696),
            .I(N__6688));
    Span4Mux_v I__595 (
            .O(N__6693),
            .I(N__6685));
    SRMux I__594 (
            .O(N__6692),
            .I(N__6682));
    SRMux I__593 (
            .O(N__6691),
            .I(N__6679));
    LocalMux I__592 (
            .O(N__6688),
            .I(N__6676));
    Span4Mux_v I__591 (
            .O(N__6685),
            .I(N__6671));
    LocalMux I__590 (
            .O(N__6682),
            .I(N__6671));
    LocalMux I__589 (
            .O(N__6679),
            .I(N__6668));
    Span4Mux_v I__588 (
            .O(N__6676),
            .I(N__6663));
    Span4Mux_v I__587 (
            .O(N__6671),
            .I(N__6663));
    Span4Mux_h I__586 (
            .O(N__6668),
            .I(N__6660));
    Odrv4 I__585 (
            .O(N__6663),
            .I(\line_buffer.n762 ));
    Odrv4 I__584 (
            .O(N__6660),
            .I(\line_buffer.n762 ));
    InMux I__583 (
            .O(N__6655),
            .I(N__6651));
    InMux I__582 (
            .O(N__6654),
            .I(N__6648));
    LocalMux I__581 (
            .O(N__6651),
            .I(N__6641));
    LocalMux I__580 (
            .O(N__6648),
            .I(N__6641));
    InMux I__579 (
            .O(N__6647),
            .I(N__6638));
    InMux I__578 (
            .O(N__6646),
            .I(N__6635));
    Span4Mux_v I__577 (
            .O(N__6641),
            .I(N__6627));
    LocalMux I__576 (
            .O(N__6638),
            .I(N__6627));
    LocalMux I__575 (
            .O(N__6635),
            .I(N__6627));
    InMux I__574 (
            .O(N__6634),
            .I(N__6623));
    Span4Mux_v I__573 (
            .O(N__6627),
            .I(N__6620));
    InMux I__572 (
            .O(N__6626),
            .I(N__6617));
    LocalMux I__571 (
            .O(N__6623),
            .I(N__6614));
    Span4Mux_v I__570 (
            .O(N__6620),
            .I(N__6609));
    LocalMux I__569 (
            .O(N__6617),
            .I(N__6609));
    Span4Mux_v I__568 (
            .O(N__6614),
            .I(N__6604));
    Span4Mux_v I__567 (
            .O(N__6609),
            .I(N__6601));
    InMux I__566 (
            .O(N__6608),
            .I(N__6598));
    InMux I__565 (
            .O(N__6607),
            .I(N__6595));
    Sp12to4 I__564 (
            .O(N__6604),
            .I(N__6592));
    Span4Mux_h I__563 (
            .O(N__6601),
            .I(N__6589));
    LocalMux I__562 (
            .O(N__6598),
            .I(N__6586));
    LocalMux I__561 (
            .O(N__6595),
            .I(N__6583));
    Span12Mux_h I__560 (
            .O(N__6592),
            .I(N__6580));
    Span4Mux_h I__559 (
            .O(N__6589),
            .I(N__6577));
    Span4Mux_h I__558 (
            .O(N__6586),
            .I(N__6574));
    Span4Mux_h I__557 (
            .O(N__6583),
            .I(N__6571));
    Span12Mux_v I__556 (
            .O(N__6580),
            .I(N__6566));
    Sp12to4 I__555 (
            .O(N__6577),
            .I(N__6566));
    IoSpan4Mux I__554 (
            .O(N__6574),
            .I(N__6563));
    Span4Mux_h I__553 (
            .O(N__6571),
            .I(N__6560));
    Span12Mux_v I__552 (
            .O(N__6566),
            .I(N__6557));
    IoSpan4Mux I__551 (
            .O(N__6563),
            .I(N__6554));
    Span4Mux_h I__550 (
            .O(N__6560),
            .I(N__6551));
    Odrv12 I__549 (
            .O(N__6557),
            .I(TVP_VIDEO_c_8));
    Odrv4 I__548 (
            .O(N__6554),
            .I(TVP_VIDEO_c_8));
    Odrv4 I__547 (
            .O(N__6551),
            .I(TVP_VIDEO_c_8));
    InMux I__546 (
            .O(N__6544),
            .I(N__6540));
    InMux I__545 (
            .O(N__6543),
            .I(N__6537));
    LocalMux I__544 (
            .O(N__6540),
            .I(N__6531));
    LocalMux I__543 (
            .O(N__6537),
            .I(N__6531));
    InMux I__542 (
            .O(N__6536),
            .I(N__6528));
    Span4Mux_v I__541 (
            .O(N__6531),
            .I(N__6523));
    LocalMux I__540 (
            .O(N__6528),
            .I(N__6523));
    Span4Mux_v I__539 (
            .O(N__6523),
            .I(N__6518));
    InMux I__538 (
            .O(N__6522),
            .I(N__6515));
    InMux I__537 (
            .O(N__6521),
            .I(N__6511));
    Span4Mux_v I__536 (
            .O(N__6518),
            .I(N__6506));
    LocalMux I__535 (
            .O(N__6515),
            .I(N__6506));
    InMux I__534 (
            .O(N__6514),
            .I(N__6503));
    LocalMux I__533 (
            .O(N__6511),
            .I(N__6500));
    Span4Mux_h I__532 (
            .O(N__6506),
            .I(N__6497));
    LocalMux I__531 (
            .O(N__6503),
            .I(N__6494));
    Span12Mux_s11_h I__530 (
            .O(N__6500),
            .I(N__6490));
    Sp12to4 I__529 (
            .O(N__6497),
            .I(N__6487));
    Span12Mux_s8_h I__528 (
            .O(N__6494),
            .I(N__6484));
    InMux I__527 (
            .O(N__6493),
            .I(N__6481));
    Span12Mux_h I__526 (
            .O(N__6490),
            .I(N__6478));
    Span12Mux_v I__525 (
            .O(N__6487),
            .I(N__6475));
    Span12Mux_v I__524 (
            .O(N__6484),
            .I(N__6472));
    LocalMux I__523 (
            .O(N__6481),
            .I(N__6469));
    Span12Mux_v I__522 (
            .O(N__6478),
            .I(N__6465));
    Span12Mux_h I__521 (
            .O(N__6475),
            .I(N__6462));
    Span12Mux_v I__520 (
            .O(N__6472),
            .I(N__6459));
    Span4Mux_h I__519 (
            .O(N__6469),
            .I(N__6456));
    InMux I__518 (
            .O(N__6468),
            .I(N__6453));
    Odrv12 I__517 (
            .O(N__6465),
            .I(TVP_VIDEO_c_9));
    Odrv12 I__516 (
            .O(N__6462),
            .I(TVP_VIDEO_c_9));
    Odrv12 I__515 (
            .O(N__6459),
            .I(TVP_VIDEO_c_9));
    Odrv4 I__514 (
            .O(N__6456),
            .I(TVP_VIDEO_c_9));
    LocalMux I__513 (
            .O(N__6453),
            .I(TVP_VIDEO_c_9));
    InMux I__512 (
            .O(N__6442),
            .I(N__6437));
    InMux I__511 (
            .O(N__6441),
            .I(N__6433));
    InMux I__510 (
            .O(N__6440),
            .I(N__6429));
    LocalMux I__509 (
            .O(N__6437),
            .I(N__6426));
    InMux I__508 (
            .O(N__6436),
            .I(N__6423));
    LocalMux I__507 (
            .O(N__6433),
            .I(N__6420));
    InMux I__506 (
            .O(N__6432),
            .I(N__6417));
    LocalMux I__505 (
            .O(N__6429),
            .I(N__6414));
    Span4Mux_h I__504 (
            .O(N__6426),
            .I(N__6411));
    LocalMux I__503 (
            .O(N__6423),
            .I(N__6408));
    Span4Mux_v I__502 (
            .O(N__6420),
            .I(N__6403));
    LocalMux I__501 (
            .O(N__6417),
            .I(N__6403));
    Span4Mux_v I__500 (
            .O(N__6414),
            .I(N__6399));
    Span4Mux_h I__499 (
            .O(N__6411),
            .I(N__6396));
    Span4Mux_h I__498 (
            .O(N__6408),
            .I(N__6393));
    Span4Mux_v I__497 (
            .O(N__6403),
            .I(N__6390));
    InMux I__496 (
            .O(N__6402),
            .I(N__6385));
    Sp12to4 I__495 (
            .O(N__6399),
            .I(N__6382));
    Sp12to4 I__494 (
            .O(N__6396),
            .I(N__6379));
    Span4Mux_h I__493 (
            .O(N__6393),
            .I(N__6376));
    Span4Mux_v I__492 (
            .O(N__6390),
            .I(N__6373));
    InMux I__491 (
            .O(N__6389),
            .I(N__6370));
    InMux I__490 (
            .O(N__6388),
            .I(N__6367));
    LocalMux I__489 (
            .O(N__6385),
            .I(N__6364));
    Span12Mux_h I__488 (
            .O(N__6382),
            .I(N__6359));
    Span12Mux_s9_v I__487 (
            .O(N__6379),
            .I(N__6359));
    Sp12to4 I__486 (
            .O(N__6376),
            .I(N__6356));
    Sp12to4 I__485 (
            .O(N__6373),
            .I(N__6351));
    LocalMux I__484 (
            .O(N__6370),
            .I(N__6351));
    LocalMux I__483 (
            .O(N__6367),
            .I(N__6348));
    Span4Mux_h I__482 (
            .O(N__6364),
            .I(N__6345));
    Span12Mux_v I__481 (
            .O(N__6359),
            .I(N__6342));
    Span12Mux_v I__480 (
            .O(N__6356),
            .I(N__6335));
    Span12Mux_h I__479 (
            .O(N__6351),
            .I(N__6335));
    Span12Mux_h I__478 (
            .O(N__6348),
            .I(N__6335));
    Span4Mux_h I__477 (
            .O(N__6345),
            .I(N__6332));
    Odrv12 I__476 (
            .O(N__6342),
            .I(TVP_VIDEO_c_7));
    Odrv12 I__475 (
            .O(N__6335),
            .I(TVP_VIDEO_c_7));
    Odrv4 I__474 (
            .O(N__6332),
            .I(TVP_VIDEO_c_7));
    InMux I__473 (
            .O(N__6325),
            .I(N__6321));
    InMux I__472 (
            .O(N__6324),
            .I(N__6318));
    LocalMux I__471 (
            .O(N__6321),
            .I(N__6315));
    LocalMux I__470 (
            .O(N__6318),
            .I(N__6311));
    Span4Mux_v I__469 (
            .O(N__6315),
            .I(N__6308));
    InMux I__468 (
            .O(N__6314),
            .I(N__6305));
    Span4Mux_v I__467 (
            .O(N__6311),
            .I(N__6301));
    Span4Mux_v I__466 (
            .O(N__6308),
            .I(N__6296));
    LocalMux I__465 (
            .O(N__6305),
            .I(N__6296));
    InMux I__464 (
            .O(N__6304),
            .I(N__6293));
    Span4Mux_v I__463 (
            .O(N__6301),
            .I(N__6290));
    Span4Mux_v I__462 (
            .O(N__6296),
            .I(N__6284));
    LocalMux I__461 (
            .O(N__6293),
            .I(N__6284));
    Span4Mux_v I__460 (
            .O(N__6290),
            .I(N__6280));
    InMux I__459 (
            .O(N__6289),
            .I(N__6277));
    Span4Mux_v I__458 (
            .O(N__6284),
            .I(N__6273));
    InMux I__457 (
            .O(N__6283),
            .I(N__6270));
    Span4Mux_v I__456 (
            .O(N__6280),
            .I(N__6265));
    LocalMux I__455 (
            .O(N__6277),
            .I(N__6265));
    InMux I__454 (
            .O(N__6276),
            .I(N__6262));
    Span4Mux_v I__453 (
            .O(N__6273),
            .I(N__6257));
    LocalMux I__452 (
            .O(N__6270),
            .I(N__6257));
    Span4Mux_v I__451 (
            .O(N__6265),
            .I(N__6252));
    LocalMux I__450 (
            .O(N__6262),
            .I(N__6252));
    Span4Mux_v I__449 (
            .O(N__6257),
            .I(N__6248));
    Span4Mux_v I__448 (
            .O(N__6252),
            .I(N__6245));
    InMux I__447 (
            .O(N__6251),
            .I(N__6242));
    Sp12to4 I__446 (
            .O(N__6248),
            .I(N__6239));
    Span4Mux_v I__445 (
            .O(N__6245),
            .I(N__6234));
    LocalMux I__444 (
            .O(N__6242),
            .I(N__6234));
    Span12Mux_h I__443 (
            .O(N__6239),
            .I(N__6231));
    Span4Mux_h I__442 (
            .O(N__6234),
            .I(N__6228));
    Odrv12 I__441 (
            .O(N__6231),
            .I(TVP_VIDEO_c_6));
    Odrv4 I__440 (
            .O(N__6228),
            .I(TVP_VIDEO_c_6));
    InMux I__439 (
            .O(N__6223),
            .I(N__6219));
    InMux I__438 (
            .O(N__6222),
            .I(N__6216));
    LocalMux I__437 (
            .O(N__6219),
            .I(N__6212));
    LocalMux I__436 (
            .O(N__6216),
            .I(N__6209));
    InMux I__435 (
            .O(N__6215),
            .I(N__6206));
    Sp12to4 I__434 (
            .O(N__6212),
            .I(N__6202));
    Span4Mux_h I__433 (
            .O(N__6209),
            .I(N__6199));
    LocalMux I__432 (
            .O(N__6206),
            .I(N__6196));
    InMux I__431 (
            .O(N__6205),
            .I(N__6192));
    Span12Mux_h I__430 (
            .O(N__6202),
            .I(N__6187));
    Span4Mux_h I__429 (
            .O(N__6199),
            .I(N__6184));
    Span4Mux_v I__428 (
            .O(N__6196),
            .I(N__6181));
    InMux I__427 (
            .O(N__6195),
            .I(N__6178));
    LocalMux I__426 (
            .O(N__6192),
            .I(N__6175));
    InMux I__425 (
            .O(N__6191),
            .I(N__6172));
    InMux I__424 (
            .O(N__6190),
            .I(N__6168));
    Span12Mux_v I__423 (
            .O(N__6187),
            .I(N__6163));
    Sp12to4 I__422 (
            .O(N__6184),
            .I(N__6163));
    Sp12to4 I__421 (
            .O(N__6181),
            .I(N__6160));
    LocalMux I__420 (
            .O(N__6178),
            .I(N__6157));
    Span12Mux_h I__419 (
            .O(N__6175),
            .I(N__6154));
    LocalMux I__418 (
            .O(N__6172),
            .I(N__6151));
    InMux I__417 (
            .O(N__6171),
            .I(N__6148));
    LocalMux I__416 (
            .O(N__6168),
            .I(N__6145));
    Span12Mux_v I__415 (
            .O(N__6163),
            .I(N__6140));
    Span12Mux_h I__414 (
            .O(N__6160),
            .I(N__6140));
    Span12Mux_h I__413 (
            .O(N__6157),
            .I(N__6137));
    Span12Mux_v I__412 (
            .O(N__6154),
            .I(N__6130));
    Span12Mux_h I__411 (
            .O(N__6151),
            .I(N__6130));
    LocalMux I__410 (
            .O(N__6148),
            .I(N__6130));
    Span4Mux_h I__409 (
            .O(N__6145),
            .I(N__6127));
    Span12Mux_h I__408 (
            .O(N__6140),
            .I(N__6122));
    Span12Mux_v I__407 (
            .O(N__6137),
            .I(N__6122));
    Span12Mux_h I__406 (
            .O(N__6130),
            .I(N__6117));
    Sp12to4 I__405 (
            .O(N__6127),
            .I(N__6117));
    Odrv12 I__404 (
            .O(N__6122),
            .I(TVP_VIDEO_c_3));
    Odrv12 I__403 (
            .O(N__6117),
            .I(TVP_VIDEO_c_3));
    InMux I__402 (
            .O(N__6112),
            .I(N__6108));
    InMux I__401 (
            .O(N__6111),
            .I(N__6105));
    LocalMux I__400 (
            .O(N__6108),
            .I(N__6102));
    LocalMux I__399 (
            .O(N__6105),
            .I(N__6098));
    Span4Mux_v I__398 (
            .O(N__6102),
            .I(N__6095));
    InMux I__397 (
            .O(N__6101),
            .I(N__6092));
    Span4Mux_v I__396 (
            .O(N__6098),
            .I(N__6089));
    Span4Mux_v I__395 (
            .O(N__6095),
            .I(N__6083));
    LocalMux I__394 (
            .O(N__6092),
            .I(N__6083));
    Span4Mux_v I__393 (
            .O(N__6089),
            .I(N__6079));
    InMux I__392 (
            .O(N__6088),
            .I(N__6076));
    Span4Mux_v I__391 (
            .O(N__6083),
            .I(N__6073));
    InMux I__390 (
            .O(N__6082),
            .I(N__6070));
    Span4Mux_v I__389 (
            .O(N__6079),
            .I(N__6064));
    LocalMux I__388 (
            .O(N__6076),
            .I(N__6064));
    Span4Mux_v I__387 (
            .O(N__6073),
            .I(N__6058));
    LocalMux I__386 (
            .O(N__6070),
            .I(N__6058));
    InMux I__385 (
            .O(N__6069),
            .I(N__6055));
    Span4Mux_v I__384 (
            .O(N__6064),
            .I(N__6052));
    InMux I__383 (
            .O(N__6063),
            .I(N__6049));
    Span4Mux_v I__382 (
            .O(N__6058),
            .I(N__6044));
    LocalMux I__381 (
            .O(N__6055),
            .I(N__6044));
    Span4Mux_v I__380 (
            .O(N__6052),
            .I(N__6039));
    LocalMux I__379 (
            .O(N__6049),
            .I(N__6039));
    Span4Mux_v I__378 (
            .O(N__6044),
            .I(N__6035));
    Span4Mux_v I__377 (
            .O(N__6039),
            .I(N__6032));
    InMux I__376 (
            .O(N__6038),
            .I(N__6029));
    Sp12to4 I__375 (
            .O(N__6035),
            .I(N__6026));
    Span4Mux_v I__374 (
            .O(N__6032),
            .I(N__6021));
    LocalMux I__373 (
            .O(N__6029),
            .I(N__6021));
    Span12Mux_h I__372 (
            .O(N__6026),
            .I(N__6018));
    Span4Mux_h I__371 (
            .O(N__6021),
            .I(N__6015));
    Odrv12 I__370 (
            .O(N__6018),
            .I(TVP_VIDEO_c_5));
    Odrv4 I__369 (
            .O(N__6015),
            .I(TVP_VIDEO_c_5));
    InMux I__368 (
            .O(N__6010),
            .I(N__6007));
    LocalMux I__367 (
            .O(N__6007),
            .I(N__6004));
    Span4Mux_v I__366 (
            .O(N__6004),
            .I(N__5998));
    InMux I__365 (
            .O(N__6003),
            .I(N__5995));
    InMux I__364 (
            .O(N__6002),
            .I(N__5991));
    InMux I__363 (
            .O(N__6001),
            .I(N__5987));
    Span4Mux_v I__362 (
            .O(N__5998),
            .I(N__5982));
    LocalMux I__361 (
            .O(N__5995),
            .I(N__5982));
    InMux I__360 (
            .O(N__5994),
            .I(N__5979));
    LocalMux I__359 (
            .O(N__5991),
            .I(N__5976));
    InMux I__358 (
            .O(N__5990),
            .I(N__5973));
    LocalMux I__357 (
            .O(N__5987),
            .I(N__5970));
    Span4Mux_v I__356 (
            .O(N__5982),
            .I(N__5965));
    LocalMux I__355 (
            .O(N__5979),
            .I(N__5965));
    Span4Mux_h I__354 (
            .O(N__5976),
            .I(N__5962));
    LocalMux I__353 (
            .O(N__5973),
            .I(N__5959));
    Span4Mux_s1_v I__352 (
            .O(N__5970),
            .I(N__5955));
    Span4Mux_v I__351 (
            .O(N__5965),
            .I(N__5952));
    Span4Mux_h I__350 (
            .O(N__5962),
            .I(N__5949));
    Span4Mux_h I__349 (
            .O(N__5959),
            .I(N__5946));
    InMux I__348 (
            .O(N__5958),
            .I(N__5943));
    Sp12to4 I__347 (
            .O(N__5955),
            .I(N__5940));
    Sp12to4 I__346 (
            .O(N__5952),
            .I(N__5937));
    Span4Mux_h I__345 (
            .O(N__5949),
            .I(N__5934));
    Span4Mux_v I__344 (
            .O(N__5946),
            .I(N__5931));
    LocalMux I__343 (
            .O(N__5943),
            .I(N__5928));
    Span12Mux_s10_h I__342 (
            .O(N__5940),
            .I(N__5924));
    Span12Mux_s9_h I__341 (
            .O(N__5937),
            .I(N__5921));
    Span4Mux_h I__340 (
            .O(N__5934),
            .I(N__5914));
    Span4Mux_v I__339 (
            .O(N__5931),
            .I(N__5914));
    Span4Mux_h I__338 (
            .O(N__5928),
            .I(N__5914));
    InMux I__337 (
            .O(N__5927),
            .I(N__5911));
    Span12Mux_v I__336 (
            .O(N__5924),
            .I(N__5908));
    Span12Mux_v I__335 (
            .O(N__5921),
            .I(N__5905));
    Span4Mux_v I__334 (
            .O(N__5914),
            .I(N__5902));
    LocalMux I__333 (
            .O(N__5911),
            .I(N__5899));
    Span12Mux_v I__332 (
            .O(N__5908),
            .I(N__5896));
    Span12Mux_h I__331 (
            .O(N__5905),
            .I(N__5893));
    Span4Mux_v I__330 (
            .O(N__5902),
            .I(N__5890));
    Span4Mux_h I__329 (
            .O(N__5899),
            .I(N__5887));
    Odrv12 I__328 (
            .O(N__5896),
            .I(TVP_VIDEO_c_4));
    Odrv12 I__327 (
            .O(N__5893),
            .I(TVP_VIDEO_c_4));
    Odrv4 I__326 (
            .O(N__5890),
            .I(TVP_VIDEO_c_4));
    Odrv4 I__325 (
            .O(N__5887),
            .I(TVP_VIDEO_c_4));
    INV INVADV_R__i2C (
            .O(INVADV_R__i2C_net),
            .I(N__17333));
    INV INVADV_R__i6C (
            .O(INVADV_R__i6C_net),
            .I(N__17196));
    INV INVADV_R__i3C (
            .O(INVADV_R__i3C_net),
            .I(N__17411));
    INV INVADV_R__i1C (
            .O(INVADV_R__i1C_net),
            .I(N__17495));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n2773 ),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\transmit_module.n2747 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(\receive_module.rx_counter.n2765 ),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\receive_module.rx_counter.n2789 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\receive_module.n2734 ),
            .carryinitout(bfn_18_15_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_9_13_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_9_13_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_LC_9_13_5  (
            .in0(N__18151),
            .in1(N__18070),
            .in2(N__17972),
            .in3(N__17780),
            .lcout(\line_buffer.n730 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1639_2_lut_3_lut_4_lut_LC_9_17_2 .C_ON=1'b0;
    defparam \line_buffer.i1639_2_lut_3_lut_4_lut_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1639_2_lut_3_lut_4_lut_LC_9_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \line_buffer.i1639_2_lut_3_lut_4_lut_LC_9_17_2  (
            .in0(N__17812),
            .in1(N__18139),
            .in2(N__17971),
            .in3(N__18068),
            .lcout(\line_buffer.n632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_9_17_7 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_9_17_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_9_17_7  (
            .in0(N__18069),
            .in1(N__17952),
            .in2(N__18149),
            .in3(N__17811),
            .lcout(\line_buffer.n762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1584_3_lut_LC_9_20_5 .C_ON=1'b0;
    defparam \line_buffer.i1584_3_lut_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1584_3_lut_LC_9_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i1584_3_lut_LC_9_20_5  (
            .in0(N__18474),
            .in1(N__7021),
            .in2(_gnd_net_),
            .in3(N__7009),
            .lcout(\line_buffer.n3028 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_LC_10_13_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_LC_10_13_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_LC_10_13_2  (
            .in0(N__7101),
            .in1(N__7118),
            .in2(_gnd_net_),
            .in3(N__6949),
            .lcout(),
            .ltout(\receive_module.rx_counter.n2975_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i38_4_lut_LC_10_13_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i38_4_lut_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i38_4_lut_LC_10_13_3 .LUT_INIT=16'b1010100010111001;
    LogicCell40 \receive_module.rx_counter.i38_4_lut_LC_10_13_3  (
            .in0(N__7060),
            .in1(N__7081),
            .in2(N__6997),
            .in3(N__6940),
            .lcout(\receive_module.rx_counter.n31_adj_572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_10_13_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_10_13_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_10_13_4  (
            .in0(N__18150),
            .in1(N__18067),
            .in2(N__17980),
            .in3(N__17762),
            .lcout(\line_buffer.n698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_adj_19_LC_10_13_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_adj_19_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_adj_19_LC_10_13_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_adj_19_LC_10_13_6  (
            .in0(N__7164),
            .in1(N__7134),
            .in2(_gnd_net_),
            .in3(N__7149),
            .lcout(\receive_module.rx_counter.n2900 ),
            .ltout(\receive_module.rx_counter.n2900_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1499_3_lut_LC_10_13_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1499_3_lut_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1499_3_lut_LC_10_13_7 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \receive_module.rx_counter.i1499_3_lut_LC_10_13_7  (
            .in0(N__7119),
            .in1(_gnd_net_),
            .in2(N__6943),
            .in3(N__7102),
            .lcout(\receive_module.rx_counter.n2943 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.X_284__i0_LC_10_14_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i0_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i0_LC_10_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i0_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__6934),
            .in2(_gnd_net_),
            .in3(N__6928),
            .lcout(\receive_module.rx_counter.n10 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\receive_module.rx_counter.n2782 ),
            .clk(N__16101),
            .ce(),
            .sr(N__7044));
    defparam \receive_module.rx_counter.X_284__i1_LC_10_14_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i1_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i1_LC_10_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i1_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__6925),
            .in2(_gnd_net_),
            .in3(N__6919),
            .lcout(\receive_module.rx_counter.n9 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2782 ),
            .carryout(\receive_module.rx_counter.n2783 ),
            .clk(N__16101),
            .ce(),
            .sr(N__7044));
    defparam \receive_module.rx_counter.X_284__i2_LC_10_14_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i2_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i2_LC_10_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i2_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__6916),
            .in2(_gnd_net_),
            .in3(N__6910),
            .lcout(\receive_module.rx_counter.n8 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2783 ),
            .carryout(\receive_module.rx_counter.n2784 ),
            .clk(N__16101),
            .ce(),
            .sr(N__7044));
    defparam \receive_module.rx_counter.X_284__i3_LC_10_14_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i3_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i3_LC_10_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i3_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__7165),
            .in2(_gnd_net_),
            .in3(N__7153),
            .lcout(\receive_module.rx_counter.X_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2784 ),
            .carryout(\receive_module.rx_counter.n2785 ),
            .clk(N__16101),
            .ce(),
            .sr(N__7044));
    defparam \receive_module.rx_counter.X_284__i4_LC_10_14_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i4_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i4_LC_10_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i4_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__7150),
            .in2(_gnd_net_),
            .in3(N__7138),
            .lcout(\receive_module.rx_counter.X_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2785 ),
            .carryout(\receive_module.rx_counter.n2786 ),
            .clk(N__16101),
            .ce(),
            .sr(N__7044));
    defparam \receive_module.rx_counter.X_284__i5_LC_10_14_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i5_LC_10_14_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i5_LC_10_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i5_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__7135),
            .in2(_gnd_net_),
            .in3(N__7123),
            .lcout(\receive_module.rx_counter.X_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2786 ),
            .carryout(\receive_module.rx_counter.n2787 ),
            .clk(N__16101),
            .ce(),
            .sr(N__7044));
    defparam \receive_module.rx_counter.X_284__i6_LC_10_14_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i6_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i6_LC_10_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i6_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__7120),
            .in2(_gnd_net_),
            .in3(N__7105),
            .lcout(\receive_module.rx_counter.X_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2787 ),
            .carryout(\receive_module.rx_counter.n2788 ),
            .clk(N__16101),
            .ce(),
            .sr(N__7044));
    defparam \receive_module.rx_counter.X_284__i7_LC_10_14_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i7_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i7_LC_10_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i7_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__7100),
            .in2(_gnd_net_),
            .in3(N__7084),
            .lcout(\receive_module.rx_counter.X_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2788 ),
            .carryout(\receive_module.rx_counter.n2789 ),
            .clk(N__16101),
            .ce(),
            .sr(N__7044));
    defparam \receive_module.rx_counter.X_284__i8_LC_10_15_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_284__i8_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i8_LC_10_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i8_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__7080),
            .in2(_gnd_net_),
            .in3(N__7066),
            .lcout(\receive_module.rx_counter.X_8 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\receive_module.rx_counter.n2790 ),
            .clk(N__16103),
            .ce(),
            .sr(N__7045));
    defparam \receive_module.rx_counter.X_284__i9_LC_10_15_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.X_284__i9_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_284__i9_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_284__i9_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__7059),
            .in2(_gnd_net_),
            .in3(N__7063),
            .lcout(\receive_module.rx_counter.X_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16103),
            .ce(),
            .sr(N__7045));
    defparam i27_1_lut_rep_20_LC_11_12_3.C_ON=1'b0;
    defparam i27_1_lut_rep_20_LC_11_12_3.SEQ_MODE=4'b0000;
    defparam i27_1_lut_rep_20_LC_11_12_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 i27_1_lut_rep_20_LC_11_12_3 (
            .in0(N__7528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n3184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_LC_11_13_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_LC_11_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__7372),
            .in2(_gnd_net_),
            .in3(N__7228),
            .lcout(),
            .ltout(\receive_module.rx_counter.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_adj_17_LC_11_13_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_adj_17_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_adj_17_LC_11_13_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_adj_17_LC_11_13_1  (
            .in0(N__7732),
            .in1(N__7702),
            .in2(N__7207),
            .in3(N__7423),
            .lcout(),
            .ltout(\receive_module.rx_counter.n2986_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i4_4_lut_adj_18_LC_11_13_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i4_4_lut_adj_18_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i4_4_lut_adj_18_LC_11_13_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \receive_module.rx_counter.i4_4_lut_adj_18_LC_11_13_2  (
            .in0(N__7475),
            .in1(N__7192),
            .in2(N__7204),
            .in3(N__7400),
            .lcout(),
            .ltout(\receive_module.rx_counter.n2989_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_adj_20_LC_11_13_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_adj_20_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_adj_20_LC_11_13_3 .LUT_INIT=16'b1111111110001111;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_adj_20_LC_11_13_3  (
            .in0(N__7250),
            .in1(N__7177),
            .in2(N__7201),
            .in3(N__7198),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_2_lut_LC_11_13_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_LC_11_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__7447),
            .in2(_gnd_net_),
            .in3(N__7249),
            .lcout(\receive_module.rx_counter.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_rep_2_2_lut_LC_11_13_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_rep_2_2_lut_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_rep_2_2_lut_LC_11_13_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \receive_module.rx_counter.i1_rep_2_2_lut_LC_11_13_5  (
            .in0(N__7448),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7474),
            .lcout(\receive_module.rx_counter.n3166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_LC_11_13_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_LC_11_13_6 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_LC_11_13_6  (
            .in0(N__7424),
            .in1(N__7703),
            .in2(N__7737),
            .in3(N__7373),
            .lcout(),
            .ltout(\receive_module.rx_counter.n2978_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_4_lut_LC_11_13_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_4_lut_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_4_lut_LC_11_13_7 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \receive_module.rx_counter.i1_4_lut_LC_11_13_7  (
            .in0(N__7229),
            .in1(N__7186),
            .in2(N__7180),
            .in3(N__7399),
            .lcout(\receive_module.rx_counter.n4_adj_571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.Y__i0_LC_12_12_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i0_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i0_LC_12_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i0_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__7733),
            .in2(_gnd_net_),
            .in3(N__7171),
            .lcout(Y_0),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\receive_module.rx_counter.n2758 ),
            .clk(N__16092),
            .ce(N__7539),
            .sr(N__15979));
    defparam \receive_module.rx_counter.Y__i1_LC_12_12_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i1_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i1_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i1_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__7704),
            .in2(_gnd_net_),
            .in3(N__7168),
            .lcout(Y_1),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2758 ),
            .carryout(\receive_module.rx_counter.n2759 ),
            .clk(N__16092),
            .ce(N__7539),
            .sr(N__15979));
    defparam \receive_module.rx_counter.Y__i2_LC_12_12_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i2_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i2_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i2_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__7425),
            .in2(_gnd_net_),
            .in3(N__7276),
            .lcout(\receive_module.rx_counter.Y_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2759 ),
            .carryout(\receive_module.rx_counter.n2760 ),
            .clk(N__16092),
            .ce(N__7539),
            .sr(N__15979));
    defparam \receive_module.rx_counter.Y__i3_LC_12_12_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i3_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i3_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i3_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__7374),
            .in2(_gnd_net_),
            .in3(N__7273),
            .lcout(\receive_module.rx_counter.Y_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2760 ),
            .carryout(\receive_module.rx_counter.n2761 ),
            .clk(N__16092),
            .ce(N__7539),
            .sr(N__15979));
    defparam \receive_module.rx_counter.Y__i4_LC_12_12_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i4_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i4_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i4_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__7230),
            .in2(_gnd_net_),
            .in3(N__7270),
            .lcout(\receive_module.rx_counter.Y_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2761 ),
            .carryout(\receive_module.rx_counter.n2762 ),
            .clk(N__16092),
            .ce(N__7539),
            .sr(N__15979));
    defparam \receive_module.rx_counter.Y__i5_LC_12_12_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i5_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i5_LC_12_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i5_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__7476),
            .in2(_gnd_net_),
            .in3(N__7267),
            .lcout(\receive_module.rx_counter.Y_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2762 ),
            .carryout(\receive_module.rx_counter.n2763 ),
            .clk(N__16092),
            .ce(N__7539),
            .sr(N__15979));
    defparam \receive_module.rx_counter.Y__i6_LC_12_12_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i6_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i6_LC_12_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i6_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__7449),
            .in2(_gnd_net_),
            .in3(N__7264),
            .lcout(\receive_module.rx_counter.Y_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2763 ),
            .carryout(\receive_module.rx_counter.n2764 ),
            .clk(N__16092),
            .ce(N__7539),
            .sr(N__15979));
    defparam \receive_module.rx_counter.Y__i7_LC_12_12_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i7_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i7_LC_12_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i7_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__7251),
            .in2(_gnd_net_),
            .in3(N__7261),
            .lcout(\receive_module.rx_counter.Y_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2764 ),
            .carryout(\receive_module.rx_counter.n2765 ),
            .clk(N__16092),
            .ce(N__7539),
            .sr(N__15979));
    defparam \receive_module.rx_counter.Y__i8_LC_12_13_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.Y__i8_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i8_LC_12_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i8_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__7401),
            .in2(_gnd_net_),
            .in3(N__7258),
            .lcout(\receive_module.rx_counter.Y_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16096),
            .ce(N__7540),
            .sr(N__15964));
    defparam \transmit_module.video_signal_controller.i1570_4_lut_LC_12_14_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1570_4_lut_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1570_4_lut_LC_12_14_1 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \transmit_module.video_signal_controller.i1570_4_lut_LC_12_14_1  (
            .in0(N__8656),
            .in1(N__8691),
            .in2(N__7327),
            .in3(N__8026),
            .lcout(\transmit_module.video_signal_controller.n3014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_21_LC_12_14_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_21_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_21_LC_12_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_21_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__7255),
            .in2(_gnd_net_),
            .in3(N__7231),
            .lcout(),
            .ltout(\receive_module.rx_counter.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i4_4_lut_adj_22_LC_12_14_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i4_4_lut_adj_22_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i4_4_lut_adj_22_LC_12_14_7 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \receive_module.rx_counter.i4_4_lut_adj_22_LC_12_14_7  (
            .in0(N__7426),
            .in1(N__7402),
            .in2(N__7378),
            .in3(N__7375),
            .lcout(n3009),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i3_3_lut_LC_12_15_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i3_3_lut_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i3_3_lut_LC_12_15_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i3_3_lut_LC_12_15_0  (
            .in0(N__7641),
            .in1(N__7625),
            .in2(_gnd_net_),
            .in3(N__7603),
            .lcout(\transmit_module.video_signal_controller.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1596_3_lut_LC_12_15_1 .C_ON=1'b0;
    defparam \line_buffer.i1596_3_lut_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1596_3_lut_LC_12_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i1596_3_lut_LC_12_15_1  (
            .in0(N__18441),
            .in1(N__7351),
            .in2(_gnd_net_),
            .in3(N__7339),
            .lcout(\line_buffer.n3040 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_2  (
            .in0(N__8050),
            .in1(N__7604),
            .in2(_gnd_net_),
            .in3(N__8081),
            .lcout(\transmit_module.video_signal_controller.n2972 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_12_15_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_12_15_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_12_15_3  (
            .in0(N__8024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8083),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_HS_48_LC_12_15_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_HS_48_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_HS_48_LC_12_15_4 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \transmit_module.video_signal_controller.VGA_HS_48_LC_12_15_4  (
            .in0(N__7291),
            .in1(N__7318),
            .in2(N__7312),
            .in3(N__8110),
            .lcout(ADV_HSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17491),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i541_3_lut_LC_12_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i541_3_lut_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i541_3_lut_LC_12_15_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \transmit_module.video_signal_controller.i541_3_lut_LC_12_15_5  (
            .in0(N__7605),
            .in1(N__7627),
            .in2(_gnd_net_),
            .in3(N__8051),
            .lcout(\transmit_module.video_signal_controller.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_18_3_lut_LC_12_15_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_18_3_lut_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_18_3_lut_LC_12_15_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_18_3_lut_LC_12_15_6  (
            .in0(N__8049),
            .in1(N__8080),
            .in2(_gnd_net_),
            .in3(N__8023),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3182_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1127_4_lut_LC_12_15_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1127_4_lut_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1127_4_lut_LC_12_15_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \transmit_module.video_signal_controller.i1127_4_lut_LC_12_15_7  (
            .in0(N__7671),
            .in1(N__7656),
            .in2(N__7285),
            .in3(N__7282),
            .lcout(\transmit_module.video_signal_controller.n2484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_12_17_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_12_17_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_12_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i9_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7762),
            .lcout(\transmit_module.X_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17424),
            .ce(N__9961),
            .sr(N__14404));
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_12_17_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_12_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_12_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i8_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7576),
            .lcout(\transmit_module.X_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17424),
            .ce(N__9961),
            .sr(N__14404));
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_12_17_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_12_17_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_12_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i7_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7570),
            .lcout(\transmit_module.X_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17424),
            .ce(N__9961),
            .sr(N__14404));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1661_LC_12_20_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1661_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1661_LC_12_20_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1661_LC_12_20_2  (
            .in0(N__18440),
            .in1(N__7564),
            .in2(N__15809),
            .in3(N__7552),
            .lcout(\line_buffer.n3101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i297_3_lut_3_lut_3_lut_LC_13_12_2 .C_ON=1'b0;
    defparam \receive_module.i297_3_lut_3_lut_3_lut_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.i297_3_lut_3_lut_3_lut_LC_13_12_2 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \receive_module.i297_3_lut_3_lut_3_lut_LC_13_12_2  (
            .in0(N__7523),
            .in1(N__7489),
            .in2(_gnd_net_),
            .in3(N__16471),
            .lcout(\receive_module.n2152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_HS_48_LC_13_12_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_HS_48_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_HS_48_LC_13_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receive_module.rx_counter.old_HS_48_LC_13_12_4  (
            .in0(N__7524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.old_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16089),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1145_4_lut_LC_13_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1145_4_lut_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1145_4_lut_LC_13_14_2 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \transmit_module.video_signal_controller.i1145_4_lut_LC_13_14_2  (
            .in0(N__8655),
            .in1(N__7483),
            .in2(N__8692),
            .in3(N__8109),
            .lcout(n2147),
            .ltout(n2147_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_3_lut_LC_13_14_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_3_lut_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_3_lut_LC_13_14_3 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \receive_module.rx_counter.i1_3_lut_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__7477),
            .in2(N__7453),
            .in3(N__7450),
            .lcout(),
            .ltout(n5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1642_4_lut_LC_13_14_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1642_4_lut_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1642_4_lut_LC_13_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \transmit_module.video_signal_controller.i1642_4_lut_LC_13_14_4  (
            .in0(N__7738),
            .in1(N__7708),
            .in2(N__7681),
            .in3(N__7678),
            .lcout(\transmit_module.video_signal_controller.n2262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i1_LC_13_15_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i1_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i1_LC_13_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i1_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__7672),
            .in2(_gnd_net_),
            .in3(N__7660),
            .lcout(\transmit_module.video_signal_controller.VGA_X_0 ),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\transmit_module.video_signal_controller.n2766 ),
            .clk(N__17516),
            .ce(),
            .sr(N__8158));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i2_LC_13_15_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i2_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i2_LC_13_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i2_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__7657),
            .in2(_gnd_net_),
            .in3(N__7645),
            .lcout(\transmit_module.video_signal_controller.VGA_X_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2766 ),
            .carryout(\transmit_module.video_signal_controller.n2767 ),
            .clk(N__17516),
            .ce(),
            .sr(N__8158));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i3_LC_13_15_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i3_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i3_LC_13_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i3_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__7642),
            .in2(_gnd_net_),
            .in3(N__7630),
            .lcout(\transmit_module.video_signal_controller.VGA_X_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2767 ),
            .carryout(\transmit_module.video_signal_controller.n2768 ),
            .clk(N__17516),
            .ce(),
            .sr(N__8158));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i4_LC_13_15_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i4_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i4_LC_13_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i4_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__7626),
            .in2(_gnd_net_),
            .in3(N__7609),
            .lcout(\transmit_module.video_signal_controller.VGA_X_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2768 ),
            .carryout(\transmit_module.video_signal_controller.n2769 ),
            .clk(N__17516),
            .ce(),
            .sr(N__8158));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i5_LC_13_15_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i5_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i5_LC_13_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i5_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__7606),
            .in2(_gnd_net_),
            .in3(N__7588),
            .lcout(\transmit_module.video_signal_controller.VGA_X_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2769 ),
            .carryout(\transmit_module.video_signal_controller.n2770 ),
            .clk(N__17516),
            .ce(),
            .sr(N__8158));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i6_LC_13_15_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i6_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i6_LC_13_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i6_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__8052),
            .in2(_gnd_net_),
            .in3(N__7585),
            .lcout(\transmit_module.video_signal_controller.VGA_X_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2770 ),
            .carryout(\transmit_module.video_signal_controller.n2771 ),
            .clk(N__17516),
            .ce(),
            .sr(N__8158));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i7_LC_13_15_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i7_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i7_LC_13_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i7_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__8082),
            .in2(_gnd_net_),
            .in3(N__7582),
            .lcout(\transmit_module.video_signal_controller.VGA_X_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2771 ),
            .carryout(\transmit_module.video_signal_controller.n2772 ),
            .clk(N__17516),
            .ce(),
            .sr(N__8158));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i8_LC_13_15_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i8_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i8_LC_13_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i8_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(N__8025),
            .in2(_gnd_net_),
            .in3(N__7579),
            .lcout(\transmit_module.video_signal_controller.VGA_X_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2772 ),
            .carryout(\transmit_module.video_signal_controller.n2773 ),
            .clk(N__17516),
            .ce(),
            .sr(N__8158));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i9_LC_13_16_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i9_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i9_LC_13_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i9_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__8108),
            .in2(_gnd_net_),
            .in3(N__7777),
            .lcout(\transmit_module.video_signal_controller.VGA_X_8 ),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\transmit_module.video_signal_controller.n2774 ),
            .clk(N__17474),
            .ce(),
            .sr(N__8157));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i10_LC_13_16_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i10_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i10_LC_13_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i10_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__8686),
            .in2(_gnd_net_),
            .in3(N__7774),
            .lcout(\transmit_module.video_signal_controller.VGA_X_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2774 ),
            .carryout(\transmit_module.video_signal_controller.n2775 ),
            .clk(N__17474),
            .ce(),
            .sr(N__8157));
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i11_LC_13_16_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i11_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_288_289__i11_LC_13_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_288_289__i11_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__8653),
            .in2(_gnd_net_),
            .in3(N__7771),
            .lcout(\transmit_module.video_signal_controller.VGA_X_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17474),
            .ce(),
            .sr(N__8157));
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_13_17_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_13_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i12_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7768),
            .lcout(\transmit_module.X_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17423),
            .ce(N__9955),
            .sr(N__14413));
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_13_17_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_13_17_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_13_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i13_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7960),
            .lcout(\transmit_module.X_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17423),
            .ce(N__9955),
            .sr(N__14413));
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_13_17_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_13_17_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_13_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i15_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8613),
            .lcout(\transmit_module.X_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17423),
            .ce(N__9955),
            .sr(N__14413));
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_13_17_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_13_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i10_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7750),
            .lcout(\transmit_module.X_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17423),
            .ce(N__9955),
            .sr(N__14413));
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_13_17_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_13_17_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i11_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7756),
            .lcout(\transmit_module.X_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17423),
            .ce(N__9955),
            .sr(N__14413));
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_13_17_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_13_17_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_13_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i6_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7744),
            .lcout(\transmit_module.X_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17423),
            .ce(N__9955),
            .sr(N__14413));
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_13_17_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_13_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i14_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7966),
            .lcout(\transmit_module.X_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17423),
            .ce(N__9955),
            .sr(N__14413));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1696_LC_13_18_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1696_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1696_LC_13_18_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1696_LC_13_18_0  (
            .in0(N__18393),
            .in1(N__7954),
            .in2(N__15781),
            .in3(N__7945),
            .lcout(),
            .ltout(\line_buffer.n3143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3143_bdd_4_lut_LC_13_18_1 .C_ON=1'b0;
    defparam \line_buffer.n3143_bdd_4_lut_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3143_bdd_4_lut_LC_13_18_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \line_buffer.n3143_bdd_4_lut_LC_13_18_1  (
            .in0(N__7930),
            .in1(N__15745),
            .in2(N__7915),
            .in3(N__7912),
            .lcout(\line_buffer.n3146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3101_bdd_4_lut_LC_13_20_2 .C_ON=1'b0;
    defparam \line_buffer.n3101_bdd_4_lut_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3101_bdd_4_lut_LC_13_20_2 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3101_bdd_4_lut_LC_13_20_2  (
            .in0(N__7891),
            .in1(N__15772),
            .in2(N__7876),
            .in3(N__7855),
            .lcout(\line_buffer.n3104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1586_3_lut_LC_14_9_0 .C_ON=1'b0;
    defparam \line_buffer.i1586_3_lut_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1586_3_lut_LC_14_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i1586_3_lut_LC_14_9_0  (
            .in0(N__18471),
            .in1(N__7849),
            .in2(_gnd_net_),
            .in3(N__7831),
            .lcout(\line_buffer.n3030 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1656_LC_14_13_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1656_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1656_LC_14_13_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1656_LC_14_13_0  (
            .in0(N__18487),
            .in1(N__7819),
            .in2(N__15810),
            .in3(N__7804),
            .lcout(\line_buffer.n3089 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i1_LC_14_14_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i1_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i1_LC_14_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_286_287__i1_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__8124),
            .in2(_gnd_net_),
            .in3(N__7786),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_0 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\transmit_module.video_signal_controller.n2776 ),
            .clk(N__17496),
            .ce(N__8153),
            .sr(N__8131));
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i2_LC_14_14_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i2_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i2_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_286_287__i2_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__7999),
            .in2(_gnd_net_),
            .in3(N__7783),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2776 ),
            .carryout(\transmit_module.video_signal_controller.n2777 ),
            .clk(N__17496),
            .ce(N__8153),
            .sr(N__8131));
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i3_LC_14_14_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i3_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i3_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_286_287__i3_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__7983),
            .in2(_gnd_net_),
            .in3(N__7780),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2777 ),
            .carryout(\transmit_module.video_signal_controller.n2778 ),
            .clk(N__17496),
            .ce(N__8153),
            .sr(N__8131));
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i4_LC_14_14_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i4_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i4_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_286_287__i4_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__8717),
            .in2(_gnd_net_),
            .in3(N__8170),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2778 ),
            .carryout(\transmit_module.video_signal_controller.n2779 ),
            .clk(N__17496),
            .ce(N__8153),
            .sr(N__8131));
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i5_LC_14_14_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i5_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i5_LC_14_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_286_287__i5_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__8751),
            .in2(_gnd_net_),
            .in3(N__8167),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2779 ),
            .carryout(\transmit_module.video_signal_controller.n2780 ),
            .clk(N__17496),
            .ce(N__8153),
            .sr(N__8131));
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i6_LC_14_14_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i6_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i6_LC_14_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_286_287__i6_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__8263),
            .in2(_gnd_net_),
            .in3(N__8164),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n2780 ),
            .carryout(\transmit_module.video_signal_controller.n2781 ),
            .clk(N__17496),
            .ce(N__8153),
            .sr(N__8131));
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i7_LC_14_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i7_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_286_287__i7_LC_14_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_286_287__i7_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__8245),
            .in2(_gnd_net_),
            .in3(N__8161),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17496),
            .ce(N__8153),
            .sr(N__8131));
    defparam \transmit_module.video_signal_controller.i1578_3_lut_4_lut_LC_14_15_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1578_3_lut_4_lut_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1578_3_lut_4_lut_LC_14_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i1578_3_lut_4_lut_LC_14_15_0  (
            .in0(N__8244),
            .in1(N__8750),
            .in2(N__8724),
            .in3(N__8262),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3022_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VS_49_LC_14_15_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VS_49_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VS_49_LC_14_15_1 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VS_49_LC_14_15_1  (
            .in0(N__7998),
            .in1(N__8125),
            .in2(N__8113),
            .in3(N__7984),
            .lcout(ADV_VSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17490),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i511_2_lut_3_lut_4_lut_LC_14_15_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i511_2_lut_3_lut_4_lut_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i511_2_lut_3_lut_4_lut_LC_14_15_2 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \transmit_module.video_signal_controller.i511_2_lut_3_lut_4_lut_LC_14_15_2  (
            .in0(N__8101),
            .in1(N__8079),
            .in2(N__8056),
            .in3(N__8022),
            .lcout(\transmit_module.video_signal_controller.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i508_2_lut_LC_14_15_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i508_2_lut_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i508_2_lut_LC_14_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i508_2_lut_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__7997),
            .in2(_gnd_net_),
            .in3(N__7982),
            .lcout(\transmit_module.video_signal_controller.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_14_15_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_14_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__8261),
            .in2(_gnd_net_),
            .in3(N__8243),
            .lcout(\transmit_module.video_signal_controller.n3183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8230),
            .lcout(\transmit_module.X_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17436),
            .ce(N__9956),
            .sr(N__14440));
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_14_16_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_14_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i1_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8224),
            .lcout(\transmit_module.X_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17436),
            .ce(N__9956),
            .sr(N__14440));
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_14_16_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_14_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_14_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i2_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8200),
            .lcout(\transmit_module.X_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17436),
            .ce(N__9956),
            .sr(N__14440));
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_14_16_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_14_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i5_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8218),
            .lcout(\transmit_module.X_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17436),
            .ce(N__9956),
            .sr(N__14440));
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_14_16_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_14_16_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_14_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i4_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8212),
            .lcout(\transmit_module.X_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17436),
            .ce(N__9956),
            .sr(N__14440));
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_14_16_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_14_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i3_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8206),
            .lcout(\transmit_module.X_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17436),
            .ce(N__9956),
            .sr(N__14440));
    defparam \transmit_module.i1_2_lut_LC_14_17_3 .C_ON=1'b0;
    defparam \transmit_module.i1_2_lut_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1_2_lut_LC_14_17_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \transmit_module.i1_2_lut_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__14348),
            .in2(_gnd_net_),
            .in3(N__14131),
            .lcout(\transmit_module.n2200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1587_3_lut_LC_14_17_4 .C_ON=1'b0;
    defparam \line_buffer.i1587_3_lut_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1587_3_lut_LC_14_17_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i1587_3_lut_LC_14_17_4  (
            .in0(N__18386),
            .in1(N__8194),
            .in2(_gnd_net_),
            .in3(N__8185),
            .lcout(),
            .ltout(\line_buffer.n3031_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_1676_LC_14_17_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_1676_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_1676_LC_14_17_5 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_1676_LC_14_17_5  (
            .in0(N__17635),
            .in1(N__15723),
            .in2(N__8389),
            .in3(N__8386),
            .lcout(),
            .ltout(\line_buffer.n3095_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i3_LC_14_17_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i3_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i3_LC_14_17_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.dout_i3_LC_14_17_6  (
            .in0(N__17651),
            .in1(N__8275),
            .in2(N__8377),
            .in3(N__8374),
            .lcout(TX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17446),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_4 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \transmit_module.BRAM_ADDR__i7_LC_14_18_4  (
            .in0(N__14411),
            .in1(N__9897),
            .in2(N__9930),
            .in3(N__14172),
            .lcout(DEBUG_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17434),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i11_LC_14_18_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i11_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i11_LC_14_18_5 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \transmit_module.BRAM_ADDR__i11_LC_14_18_5  (
            .in0(N__14171),
            .in1(N__10634),
            .in2(N__10612),
            .in3(N__14412),
            .lcout(\transmit_module.TX_ADDR_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17434),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3089_bdd_4_lut_LC_14_19_3 .C_ON=1'b0;
    defparam \line_buffer.n3089_bdd_4_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3089_bdd_4_lut_LC_14_19_3 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \line_buffer.n3089_bdd_4_lut_LC_14_19_3  (
            .in0(N__8362),
            .in1(N__8344),
            .in2(N__15768),
            .in3(N__8323),
            .lcout(),
            .ltout(\line_buffer.n3092_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i2_LC_14_19_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i2_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i2_LC_14_19_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i2_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__17650),
            .in2(N__8314),
            .in3(N__8311),
            .lcout(TX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17412),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1595_3_lut_LC_14_21_3 .C_ON=1'b0;
    defparam \line_buffer.i1595_3_lut_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1595_3_lut_LC_14_21_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i1595_3_lut_LC_14_21_3  (
            .in0(N__8305),
            .in1(N__8293),
            .in2(_gnd_net_),
            .in3(N__18439),
            .lcout(\line_buffer.n3039 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i4_4_lut_LC_15_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i4_4_lut_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i4_4_lut_LC_15_10_1 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \receive_module.rx_counter.i4_4_lut_LC_15_10_1  (
            .in0(N__8538),
            .in1(N__8553),
            .in2(N__8587),
            .in3(N__8568),
            .lcout(\receive_module.rx_counter.n10_adj_570 ),
            .ltout(\receive_module.rx_counter.n10_adj_570_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i873_2_lut_4_lut_LC_15_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i873_2_lut_4_lut_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i873_2_lut_4_lut_LC_15_10_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \receive_module.rx_counter.i873_2_lut_4_lut_LC_15_10_2  (
            .in0(N__8846),
            .in1(N__8819),
            .in2(N__8266),
            .in3(N__10334),
            .lcout(\receive_module.rx_counter.n2227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i0_LC_15_11_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i0_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i0_LC_15_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_285__i0_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__8820),
            .in2(_gnd_net_),
            .in3(N__8590),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_0 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\receive_module.rx_counter.n2753 ),
            .clk(N__16084),
            .ce(N__10341),
            .sr(N__8521));
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i1_LC_15_11_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i1_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i1_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_285__i1_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__8586),
            .in2(_gnd_net_),
            .in3(N__8572),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2753 ),
            .carryout(\receive_module.rx_counter.n2754 ),
            .clk(N__16084),
            .ce(N__10341),
            .sr(N__8521));
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i2_LC_15_11_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i2_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i2_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_285__i2_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__8569),
            .in2(_gnd_net_),
            .in3(N__8557),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2754 ),
            .carryout(\receive_module.rx_counter.n2755 ),
            .clk(N__16084),
            .ce(N__10341),
            .sr(N__8521));
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i3_LC_15_11_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i3_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i3_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_285__i3_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__8554),
            .in2(_gnd_net_),
            .in3(N__8542),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2755 ),
            .carryout(\receive_module.rx_counter.n2756 ),
            .clk(N__16084),
            .ce(N__10341),
            .sr(N__8521));
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i4_LC_15_11_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i4_LC_15_11_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i4_LC_15_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_285__i4_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__8539),
            .in2(_gnd_net_),
            .in3(N__8527),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n2756 ),
            .carryout(\receive_module.rx_counter.n2757 ),
            .clk(N__16084),
            .ce(N__10341),
            .sr(N__8521));
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i5_LC_15_11_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i5_LC_15_11_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_285__i5_LC_15_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_285__i5_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__8848),
            .in2(_gnd_net_),
            .in3(N__8524),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16084),
            .ce(N__10341),
            .sr(N__8521));
    defparam \receive_module.i24_1_lut_rep_21_LC_15_13_3 .C_ON=1'b0;
    defparam \receive_module.i24_1_lut_rep_21_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.i24_1_lut_rep_21_LC_15_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \receive_module.i24_1_lut_rep_21_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16386),
            .lcout(\receive_module.n3185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ADV_R__i1_LC_15_14_1.C_ON=1'b0;
    defparam ADV_R__i1_LC_15_14_1.SEQ_MODE=4'b1000;
    defparam ADV_R__i1_LC_15_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i1_LC_15_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12220),
            .lcout(n1955),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__14184));
    defparam ADV_R__i3_LC_15_15_7.C_ON=1'b0;
    defparam ADV_R__i3_LC_15_15_7.SEQ_MODE=4'b1000;
    defparam ADV_R__i3_LC_15_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i3_LC_15_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8452),
            .lcout(n1953),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i3C_net),
            .ce(),
            .sr(N__14130));
    defparam \transmit_module.BRAM_ADDR__i5_LC_15_16_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i5_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i5_LC_15_16_1 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \transmit_module.BRAM_ADDR__i5_LC_15_16_1  (
            .in0(N__9384),
            .in1(N__9362),
            .in2(N__14360),
            .in3(N__14140),
            .lcout(DEBUG_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17435),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_15_16_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_15_16_3 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_LC_15_16_3  (
            .in0(N__8752),
            .in1(N__8731),
            .in2(N__8725),
            .in3(N__8698),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.VGA_VISIBLE_N_558_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1636_4_lut_4_lut_LC_15_16_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1636_4_lut_4_lut_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1636_4_lut_4_lut_LC_15_16_4 .LUT_INIT=16'b1100111110011111;
    LogicCell40 \transmit_module.video_signal_controller.i1636_4_lut_4_lut_LC_15_16_4  (
            .in0(N__8687),
            .in1(N__8654),
            .in2(N__8626),
            .in3(N__8623),
            .lcout(VGA_VISIBLE),
            .ltout(VGA_VISIBLE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i3_LC_15_16_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i3_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i3_LC_15_16_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \transmit_module.BRAM_ADDR__i3_LC_15_16_5  (
            .in0(N__14296),
            .in1(N__9126),
            .in2(N__8617),
            .in3(N__9092),
            .lcout(DEBUG_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17435),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_16_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_16_7 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \transmit_module.BRAM_ADDR__i6_LC_15_16_7  (
            .in0(N__9657),
            .in1(N__9626),
            .in2(N__14361),
            .in3(N__14141),
            .lcout(DEBUG_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17435),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_2_lut_LC_15_17_0 .C_ON=1'b1;
    defparam \transmit_module.add_15_2_lut_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_2_lut_LC_15_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_2_lut_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__14206),
            .in2(N__8614),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n388 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\transmit_module.n2740 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_3_lut_LC_15_17_1 .C_ON=1'b1;
    defparam \transmit_module.add_15_3_lut_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_3_lut_LC_15_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_3_lut_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__12085),
            .in2(_gnd_net_),
            .in3(N__8599),
            .lcout(\transmit_module.n387 ),
            .ltout(),
            .carryin(\transmit_module.n2740 ),
            .carryout(\transmit_module.n2741 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_4_lut_LC_15_17_2 .C_ON=1'b1;
    defparam \transmit_module.add_15_4_lut_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_4_lut_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_4_lut_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__9088),
            .in2(_gnd_net_),
            .in3(N__8596),
            .lcout(\transmit_module.n386 ),
            .ltout(),
            .carryin(\transmit_module.n2741 ),
            .carryout(\transmit_module.n2742 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_5_lut_LC_15_17_3 .C_ON=1'b1;
    defparam \transmit_module.add_15_5_lut_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_5_lut_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_5_lut_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__11530),
            .in2(_gnd_net_),
            .in3(N__8593),
            .lcout(\transmit_module.n385 ),
            .ltout(),
            .carryin(\transmit_module.n2742 ),
            .carryout(\transmit_module.n2743 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_6_lut_LC_15_17_4 .C_ON=1'b1;
    defparam \transmit_module.add_15_6_lut_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_6_lut_LC_15_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_6_lut_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__9358),
            .in2(_gnd_net_),
            .in3(N__8779),
            .lcout(\transmit_module.n384 ),
            .ltout(),
            .carryin(\transmit_module.n2743 ),
            .carryout(\transmit_module.n2744 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_7_lut_LC_15_17_5 .C_ON=1'b1;
    defparam \transmit_module.add_15_7_lut_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_7_lut_LC_15_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_7_lut_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__9622),
            .in2(_gnd_net_),
            .in3(N__8776),
            .lcout(\transmit_module.n383 ),
            .ltout(),
            .carryin(\transmit_module.n2744 ),
            .carryout(\transmit_module.n2745 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_8_lut_LC_15_17_6 .C_ON=1'b1;
    defparam \transmit_module.add_15_8_lut_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_8_lut_LC_15_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_8_lut_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9929),
            .in3(N__8773),
            .lcout(\transmit_module.n382 ),
            .ltout(),
            .carryin(\transmit_module.n2745 ),
            .carryout(\transmit_module.n2746 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_9_lut_LC_15_17_7 .C_ON=1'b1;
    defparam \transmit_module.add_15_9_lut_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_9_lut_LC_15_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_9_lut_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__11833),
            .in2(_gnd_net_),
            .in3(N__8770),
            .lcout(\transmit_module.n381 ),
            .ltout(),
            .carryin(\transmit_module.n2746 ),
            .carryout(\transmit_module.n2747 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_10_lut_LC_15_18_0 .C_ON=1'b1;
    defparam \transmit_module.add_15_10_lut_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_10_lut_LC_15_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_10_lut_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__10880),
            .in2(_gnd_net_),
            .in3(N__8767),
            .lcout(\transmit_module.n380 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\transmit_module.n2748 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_11_lut_LC_15_18_1 .C_ON=1'b1;
    defparam \transmit_module.add_15_11_lut_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_11_lut_LC_15_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_11_lut_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10902),
            .in3(N__8764),
            .lcout(\transmit_module.n379 ),
            .ltout(),
            .carryin(\transmit_module.n2748 ),
            .carryout(\transmit_module.n2749 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_15_12_lut_LC_15_18_2 .C_ON=1'b1;
    defparam \transmit_module.add_15_12_lut_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_15_12_lut_LC_15_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_15_12_lut_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10635),
            .in3(N__8761),
            .lcout(\transmit_module.n378 ),
            .ltout(),
            .carryin(\transmit_module.n2749 ),
            .carryout(\transmit_module.n2750 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_18_3 .C_ON=1'b1;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_18_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__18385),
            .in2(_gnd_net_),
            .in3(N__8758),
            .lcout(TX_ADDR_11),
            .ltout(),
            .carryin(\transmit_module.n2750 ),
            .carryout(\transmit_module.n2751 ),
            .clk(N__17330),
            .ce(N__9960),
            .sr(N__14445));
    defparam \transmit_module.BRAM_ADDR__rep_1_i1_LC_15_18_4 .C_ON=1'b1;
    defparam \transmit_module.BRAM_ADDR__rep_1_i1_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i1_LC_15_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i1_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__15719),
            .in2(_gnd_net_),
            .in3(N__8755),
            .lcout(TX_ADDR_12),
            .ltout(),
            .carryin(\transmit_module.n2751 ),
            .carryout(\transmit_module.n2752 ),
            .clk(N__17330),
            .ce(N__9960),
            .sr(N__14445));
    defparam \transmit_module.BRAM_ADDR__rep_1_i2_LC_15_18_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__rep_1_i2_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i2_LC_15_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i2_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__17649),
            .in2(_gnd_net_),
            .in3(N__9964),
            .lcout(TX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17330),
            .ce(N__9960),
            .sr(N__14445));
    defparam \transmit_module.i1056_4_lut_LC_15_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1056_4_lut_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1056_4_lut_LC_15_19_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1056_4_lut_LC_15_19_0  (
            .in0(N__9922),
            .in1(N__9898),
            .in2(N__14425),
            .in3(N__14164),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1057_4_lut_LC_15_19_2 .C_ON=1'b0;
    defparam \transmit_module.i1057_4_lut_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1057_4_lut_LC_15_19_2 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \transmit_module.i1057_4_lut_LC_15_19_2  (
            .in0(N__9658),
            .in1(N__9630),
            .in2(N__14427),
            .in3(N__14166),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1058_4_lut_LC_15_19_4 .C_ON=1'b0;
    defparam \transmit_module.i1058_4_lut_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1058_4_lut_LC_15_19_4 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \transmit_module.i1058_4_lut_LC_15_19_4  (
            .in0(N__9388),
            .in1(N__9366),
            .in2(N__14426),
            .in3(N__14165),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i9_LC_15_19_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i9_LC_15_19_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i9_LC_15_19_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i9_LC_15_19_5  (
            .in0(N__14167),
            .in1(N__14384),
            .in2(N__10864),
            .in3(N__10882),
            .lcout(\transmit_module.TX_ADDR_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17332),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1060_4_lut_LC_15_23_2 .C_ON=1'b0;
    defparam \transmit_module.i1060_4_lut_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1060_4_lut_LC_15_23_2 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \transmit_module.i1060_4_lut_LC_15_23_2  (
            .in0(N__9127),
            .in1(N__9102),
            .in2(N__14444),
            .in3(N__14185),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.PULSE_1HZ_46_LC_16_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.PULSE_1HZ_46_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.PULSE_1HZ_46_LC_16_10_0 .LUT_INIT=16'b1101111100100000;
    LogicCell40 \receive_module.rx_counter.PULSE_1HZ_46_LC_16_10_0  (
            .in0(N__8847),
            .in1(N__8830),
            .in2(N__8824),
            .in3(N__8790),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16080),
            .ce(N__10345),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_VS_49_LC_16_11_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_VS_49_LC_16_11_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_VS_49_LC_16_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receive_module.rx_counter.old_VS_49_LC_16_11_1  (
            .in0(N__16406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.old_VS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16082),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i141_2_lut_2_lut_LC_16_11_6 .C_ON=1'b0;
    defparam \receive_module.i141_2_lut_2_lut_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.i141_2_lut_2_lut_LC_16_11_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \receive_module.i141_2_lut_2_lut_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__10351),
            .in2(_gnd_net_),
            .in3(N__16405),
            .lcout(\receive_module.n252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ADV_R__i6_LC_16_15_2.C_ON=1'b0;
    defparam ADV_R__i6_LC_16_15_2.SEQ_MODE=4'b1000;
    defparam ADV_R__i6_LC_16_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i6_LC_16_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14803),
            .lcout(n1950),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i6C_net),
            .ce(),
            .sr(N__14101));
    defparam \transmit_module.BRAM_ADDR__i4_LC_16_16_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i4_LC_16_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i4_LC_16_16_6 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \transmit_module.BRAM_ADDR__i4_LC_16_16_6  (
            .in0(N__11571),
            .in1(N__14398),
            .in2(N__11541),
            .in3(N__14139),
            .lcout(DEBUG_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17331),
            .ce(),
            .sr(_gnd_net_));
    defparam ADV_R__i2_LC_16_17_0.C_ON=1'b0;
    defparam ADV_R__i2_LC_16_17_0.SEQ_MODE=4'b1000;
    defparam ADV_R__i2_LC_16_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i2_LC_16_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11194),
            .lcout(n1954),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14102));
    defparam ADV_R__i4_LC_16_17_3.C_ON=1'b0;
    defparam ADV_R__i4_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam ADV_R__i4_LC_16_17_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 ADV_R__i4_LC_16_17_3 (
            .in0(N__10207),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n1952),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14102));
    defparam ADV_R__i5_LC_16_17_4.C_ON=1'b0;
    defparam ADV_R__i5_LC_16_17_4.SEQ_MODE=4'b1000;
    defparam ADV_R__i5_LC_16_17_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 ADV_R__i5_LC_16_17_4 (
            .in0(N__17602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n1951),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14102));
    defparam ADV_R__i7_LC_16_17_6.C_ON=1'b0;
    defparam ADV_R__i7_LC_16_17_6.SEQ_MODE=4'b1000;
    defparam ADV_R__i7_LC_16_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i7_LC_16_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10375),
            .lcout(n1949),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14102));
    defparam ADV_R__i8_LC_16_17_7.C_ON=1'b0;
    defparam ADV_R__i8_LC_16_17_7.SEQ_MODE=4'b1000;
    defparam ADV_R__i8_LC_16_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i8_LC_16_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11284),
            .lcout(ADV_B_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14102));
    defparam \transmit_module.BRAM_ADDR__i2_LC_16_18_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i2_LC_16_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i2_LC_16_18_1 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \transmit_module.BRAM_ADDR__i2_LC_16_18_1  (
            .in0(N__14173),
            .in1(N__12114),
            .in2(N__14436),
            .in3(N__12093),
            .lcout(DEBUG_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17329),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i1_LC_16_18_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i1_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i1_LC_16_18_4 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \transmit_module.BRAM_ADDR__i1_LC_16_18_4  (
            .in0(N__14466),
            .in1(N__14174),
            .in2(N__14219),
            .in3(N__14402),
            .lcout(DEBUG_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17329),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i8_LC_16_18_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i8_LC_16_18_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i8_LC_16_18_6 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \transmit_module.BRAM_ADDR__i8_LC_16_18_6  (
            .in0(N__11835),
            .in1(N__14175),
            .in2(N__11811),
            .in3(N__14403),
            .lcout(DEBUG_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17329),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1053_4_lut_LC_16_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1053_4_lut_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1053_4_lut_LC_16_19_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1053_4_lut_LC_16_19_0  (
            .in0(N__14180),
            .in1(N__10898),
            .in2(N__14434),
            .in3(N__10911),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i10_LC_16_19_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i10_LC_16_19_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i10_LC_16_19_1 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \transmit_module.BRAM_ADDR__i10_LC_16_19_1  (
            .in0(N__10912),
            .in1(N__14397),
            .in2(N__10903),
            .in3(N__14182),
            .lcout(\transmit_module.TX_ADDR_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17195),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1054_4_lut_LC_16_19_4 .C_ON=1'b0;
    defparam \transmit_module.i1054_4_lut_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1054_4_lut_LC_16_19_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1054_4_lut_LC_16_19_4  (
            .in0(N__14181),
            .in1(N__10881),
            .in2(N__14435),
            .in3(N__10860),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1052_4_lut_LC_16_19_7 .C_ON=1'b0;
    defparam \transmit_module.i1052_4_lut_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1052_4_lut_LC_16_19_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1052_4_lut_LC_16_19_7  (
            .in0(N__10639),
            .in1(N__10608),
            .in2(N__14424),
            .in3(N__14179),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i6_LC_16_20_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i6_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i6_LC_16_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i6_LC_16_20_6  (
            .in0(N__17668),
            .in1(N__10384),
            .in2(_gnd_net_),
            .in3(N__12679),
            .lcout(TX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17249),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_0.C_ON=1'b0;
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_0 (
            .in0(N__16129),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_TVP_CLK_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i1632_2_lut_rep_17_LC_17_14_5 .C_ON=1'b0;
    defparam \receive_module.i1632_2_lut_rep_17_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.i1632_2_lut_rep_17_LC_17_14_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \receive_module.i1632_2_lut_rep_17_LC_17_14_5  (
            .in0(N__17861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16432),
            .lcout(\receive_module.n3181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i9_LC_17_15_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i9_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i9_LC_17_15_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \receive_module.BRAM_ADDR__i9_LC_17_15_2  (
            .in0(N__17869),
            .in1(N__16445),
            .in2(N__14506),
            .in3(N__14530),
            .lcout(RX_ADDR_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16087),
            .ce(),
            .sr(N__15965));
    defparam \receive_module.BRAM_ADDR__i8_LC_17_15_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i8_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i8_LC_17_15_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \receive_module.BRAM_ADDR__i8_LC_17_15_3  (
            .in0(N__12775),
            .in1(N__12751),
            .in2(N__16470),
            .in3(N__17868),
            .lcout(RX_ADDR_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16087),
            .ce(),
            .sr(N__15965));
    defparam \receive_module.BRAM_ADDR__i7_LC_17_15_4 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i7_LC_17_15_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i7_LC_17_15_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \receive_module.BRAM_ADDR__i7_LC_17_15_4  (
            .in0(N__17867),
            .in1(N__12997),
            .in2(N__16481),
            .in3(N__13021),
            .lcout(RX_ADDR_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16087),
            .ce(),
            .sr(N__15965));
    defparam \receive_module.BRAM_ADDR__i5_LC_17_15_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i5_LC_17_15_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i5_LC_17_15_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \receive_module.BRAM_ADDR__i5_LC_17_15_6  (
            .in0(N__17866),
            .in1(N__16444),
            .in2(N__13274),
            .in3(N__13246),
            .lcout(RX_ADDR_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16087),
            .ce(),
            .sr(N__15965));
    defparam \receive_module.BRAM_ADDR__i0_LC_17_15_7 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i0_LC_17_15_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i0_LC_17_15_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \receive_module.BRAM_ADDR__i0_LC_17_15_7  (
            .in0(N__16443),
            .in1(N__13507),
            .in2(N__13544),
            .in3(N__17865),
            .lcout(RX_ADDR_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16087),
            .ce(),
            .sr(N__15965));
    defparam \line_buffer.n3137_bdd_4_lut_LC_17_16_6 .C_ON=1'b0;
    defparam \line_buffer.n3137_bdd_4_lut_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3137_bdd_4_lut_LC_17_16_6 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3137_bdd_4_lut_LC_17_16_6  (
            .in0(N__11239),
            .in1(N__15777),
            .in2(N__11218),
            .in3(N__12172),
            .lcout(),
            .ltout(\line_buffer.n3140_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i1_LC_17_16_7 .C_ON=1'b0;
    defparam \line_buffer.dout_i1_LC_17_16_7 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i1_LC_17_16_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \line_buffer.dout_i1_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__17684),
            .in2(N__11197),
            .in3(N__11134),
            .lcout(TX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17419),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1666_LC_17_17_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1666_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1666_LC_17_17_3 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1666_LC_17_17_3  (
            .in0(N__18470),
            .in1(N__11188),
            .in2(N__15830),
            .in3(N__11179),
            .lcout(),
            .ltout(\line_buffer.n3107_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3107_bdd_4_lut_LC_17_17_4 .C_ON=1'b0;
    defparam \line_buffer.n3107_bdd_4_lut_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3107_bdd_4_lut_LC_17_17_4 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \line_buffer.n3107_bdd_4_lut_LC_17_17_4  (
            .in0(N__11161),
            .in1(N__11149),
            .in2(N__11137),
            .in3(N__15808),
            .lcout(\line_buffer.n3110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1691_LC_17_17_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1691_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1691_LC_17_17_6 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1691_LC_17_17_6  (
            .in0(N__18469),
            .in1(N__12208),
            .in2(N__12193),
            .in3(N__15807),
            .lcout(\line_buffer.n3137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_19_0 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_19_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_19_0  (
            .in0(N__18137),
            .in1(N__18046),
            .in2(N__17979),
            .in3(N__17878),
            .lcout(\line_buffer.n761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1061_4_lut_LC_17_19_1 .C_ON=1'b0;
    defparam \transmit_module.i1061_4_lut_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1061_4_lut_LC_17_19_1 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \transmit_module.i1061_4_lut_LC_17_19_1  (
            .in0(N__12118),
            .in1(N__12086),
            .in2(N__14443),
            .in3(N__14178),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1055_4_lut_LC_17_19_3 .C_ON=1'b0;
    defparam \transmit_module.i1055_4_lut_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1055_4_lut_LC_17_19_3 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1055_4_lut_LC_17_19_3  (
            .in0(N__11834),
            .in1(N__11812),
            .in2(N__14441),
            .in3(N__14176),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1059_4_lut_LC_17_19_7 .C_ON=1'b0;
    defparam \transmit_module.i1059_4_lut_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1059_4_lut_LC_17_19_7 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \transmit_module.i1059_4_lut_LC_17_19_7  (
            .in0(N__11575),
            .in1(N__11540),
            .in2(N__14442),
            .in3(N__14177),
            .lcout(n25_adj_573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_1681_LC_17_20_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_1681_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_1681_LC_17_20_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_1681_LC_17_20_3  (
            .in0(N__15776),
            .in1(N__11296),
            .in2(N__17685),
            .in3(N__13753),
            .lcout(),
            .ltout(\line_buffer.n3125_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i7_LC_17_20_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i7_LC_17_20_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i7_LC_17_20_4 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \line_buffer.dout_i7_LC_17_20_4  (
            .in0(N__12640),
            .in1(N__17672),
            .in2(N__11287),
            .in3(N__11245),
            .lcout(TX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17337),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1599_3_lut_LC_17_20_7 .C_ON=1'b0;
    defparam \line_buffer.i1599_3_lut_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1599_3_lut_LC_17_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i1599_3_lut_LC_17_20_7  (
            .in0(N__11275),
            .in1(N__11260),
            .in2(_gnd_net_),
            .in3(N__18450),
            .lcout(\line_buffer.n3043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_21_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_21_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_21_1  (
            .in0(N__18451),
            .in1(N__12742),
            .in2(N__15812),
            .in3(N__12727),
            .lcout(),
            .ltout(\line_buffer.n3161_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3161_bdd_4_lut_LC_17_21_2 .C_ON=1'b0;
    defparam \line_buffer.n3161_bdd_4_lut_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3161_bdd_4_lut_LC_17_21_2 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \line_buffer.n3161_bdd_4_lut_LC_17_21_2  (
            .in0(N__12712),
            .in1(N__12700),
            .in2(N__12682),
            .in3(N__15785),
            .lcout(\line_buffer.n3164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1598_3_lut_LC_17_23_1 .C_ON=1'b0;
    defparam \line_buffer.i1598_3_lut_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1598_3_lut_LC_17_23_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i1598_3_lut_LC_17_23_1  (
            .in0(N__12673),
            .in1(N__12658),
            .in2(_gnd_net_),
            .in3(N__18475),
            .lcout(\line_buffer.n3042 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_18_2_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_18_2_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_18_2_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_18_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3113_bdd_4_lut_LC_18_13_0 .C_ON=1'b0;
    defparam \line_buffer.n3113_bdd_4_lut_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3113_bdd_4_lut_LC_18_13_0 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.n3113_bdd_4_lut_LC_18_13_0  (
            .in0(N__15825),
            .in1(N__12343),
            .in2(N__12325),
            .in3(N__12271),
            .lcout(\line_buffer.n3116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1671_LC_18_13_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1671_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1671_LC_18_13_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1671_LC_18_13_4  (
            .in0(N__18477),
            .in1(N__12304),
            .in2(N__15836),
            .in3(N__12289),
            .lcout(\line_buffer.n3113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3119_bdd_4_lut_LC_18_13_5 .C_ON=1'b0;
    defparam \line_buffer.n3119_bdd_4_lut_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3119_bdd_4_lut_LC_18_13_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3119_bdd_4_lut_LC_18_13_5  (
            .in0(N__12265),
            .in1(N__15826),
            .in2(N__12247),
            .in3(N__13795),
            .lcout(),
            .ltout(\line_buffer.n3122_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i0_LC_18_13_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i0_LC_18_13_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i0_LC_18_13_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \line_buffer.dout_i0_LC_18_13_6  (
            .in0(N__17694),
            .in1(_gnd_net_),
            .in2(N__12229),
            .in3(N__12226),
            .lcout(TX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17497),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_2_lut_LC_18_14_0 .C_ON=1'b1;
    defparam \receive_module.add_12_2_lut_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_2_lut_LC_18_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_2_lut_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__13534),
            .in2(_gnd_net_),
            .in3(N__13501),
            .lcout(\receive_module.n136 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\receive_module.n2727 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_3_lut_LC_18_14_1 .C_ON=1'b1;
    defparam \receive_module.add_12_3_lut_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_3_lut_LC_18_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_3_lut_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__14873),
            .in2(_gnd_net_),
            .in3(N__13498),
            .lcout(\receive_module.n135 ),
            .ltout(),
            .carryin(\receive_module.n2727 ),
            .carryout(\receive_module.n2728 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_4_lut_LC_18_14_2 .C_ON=1'b1;
    defparam \receive_module.add_12_4_lut_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_4_lut_LC_18_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_4_lut_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__15119),
            .in2(_gnd_net_),
            .in3(N__13495),
            .lcout(\receive_module.n134 ),
            .ltout(),
            .carryin(\receive_module.n2728 ),
            .carryout(\receive_module.n2729 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_5_lut_LC_18_14_3 .C_ON=1'b1;
    defparam \receive_module.add_12_5_lut_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_5_lut_LC_18_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_5_lut_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__15356),
            .in2(_gnd_net_),
            .in3(N__13492),
            .lcout(\receive_module.n133 ),
            .ltout(),
            .carryin(\receive_module.n2729 ),
            .carryout(\receive_module.n2730 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_6_lut_LC_18_14_4 .C_ON=1'b1;
    defparam \receive_module.add_12_6_lut_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_6_lut_LC_18_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_6_lut_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__16763),
            .in2(_gnd_net_),
            .in3(N__13489),
            .lcout(\receive_module.n132 ),
            .ltout(),
            .carryin(\receive_module.n2730 ),
            .carryout(\receive_module.n2731 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_7_lut_LC_18_14_5 .C_ON=1'b1;
    defparam \receive_module.add_12_7_lut_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_7_lut_LC_18_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_7_lut_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__13265),
            .in2(_gnd_net_),
            .in3(N__13240),
            .lcout(\receive_module.n131 ),
            .ltout(),
            .carryin(\receive_module.n2731 ),
            .carryout(\receive_module.n2732 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_8_lut_LC_18_14_6 .C_ON=1'b1;
    defparam \receive_module.add_12_8_lut_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_8_lut_LC_18_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_8_lut_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__16523),
            .in2(_gnd_net_),
            .in3(N__13237),
            .lcout(\receive_module.n130 ),
            .ltout(),
            .carryin(\receive_module.n2732 ),
            .carryout(\receive_module.n2733 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_9_lut_LC_18_14_7 .C_ON=1'b1;
    defparam \receive_module.add_12_9_lut_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_9_lut_LC_18_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_9_lut_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__13022),
            .in2(_gnd_net_),
            .in3(N__12991),
            .lcout(\receive_module.n129 ),
            .ltout(),
            .carryin(\receive_module.n2733 ),
            .carryout(\receive_module.n2734 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_10_lut_LC_18_15_0 .C_ON=1'b1;
    defparam \receive_module.add_12_10_lut_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_10_lut_LC_18_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_10_lut_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__12776),
            .in2(_gnd_net_),
            .in3(N__12745),
            .lcout(\receive_module.n128 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\receive_module.n2735 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_11_lut_LC_18_15_1 .C_ON=1'b1;
    defparam \receive_module.add_12_11_lut_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_11_lut_LC_18_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_11_lut_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__14531),
            .in2(_gnd_net_),
            .in3(N__14497),
            .lcout(\receive_module.n127 ),
            .ltout(),
            .carryin(\receive_module.n2735 ),
            .carryout(\receive_module.n2736 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_12_lut_LC_18_15_2 .C_ON=1'b1;
    defparam \receive_module.add_12_12_lut_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_12_lut_LC_18_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_12_lut_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__16160),
            .in2(_gnd_net_),
            .in3(N__14494),
            .lcout(\receive_module.n126 ),
            .ltout(),
            .carryin(\receive_module.n2736 ),
            .carryout(\receive_module.n2737 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i11_LC_18_15_3 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i11_LC_18_15_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i11_LC_18_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i11_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__18007),
            .in2(_gnd_net_),
            .in3(N__14491),
            .lcout(RX_ADDR_11),
            .ltout(),
            .carryin(\receive_module.n2737 ),
            .carryout(\receive_module.n2738 ),
            .clk(N__16090),
            .ce(N__14482),
            .sr(N__15966));
    defparam \receive_module.BRAM_ADDR__i12_LC_18_15_4 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i12_LC_18_15_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i12_LC_18_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i12_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__18107),
            .in2(_gnd_net_),
            .in3(N__14488),
            .lcout(RX_ADDR_12),
            .ltout(),
            .carryin(\receive_module.n2738 ),
            .carryout(\receive_module.n2739 ),
            .clk(N__16090),
            .ce(N__14482),
            .sr(N__15966));
    defparam \receive_module.BRAM_ADDR__i13_LC_18_15_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i13_LC_18_15_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i13_LC_18_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i13_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__17925),
            .in2(_gnd_net_),
            .in3(N__14485),
            .lcout(RX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16090),
            .ce(N__14482),
            .sr(N__15966));
    defparam \transmit_module.i1096_4_lut_LC_18_19_5 .C_ON=1'b0;
    defparam \transmit_module.i1096_4_lut_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1096_4_lut_LC_18_19_5 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \transmit_module.i1096_4_lut_LC_18_19_5  (
            .in0(N__14470),
            .in1(N__14423),
            .in2(N__14229),
            .in3(N__14183),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1686_LC_18_19_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1686_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1686_LC_18_19_6 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1686_LC_18_19_6  (
            .in0(N__18448),
            .in1(N__15813),
            .in2(N__13834),
            .in3(N__13810),
            .lcout(\line_buffer.n3119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1583_3_lut_LC_18_21_3 .C_ON=1'b0;
    defparam \line_buffer.i1583_3_lut_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1583_3_lut_LC_18_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i1583_3_lut_LC_18_21_3  (
            .in0(N__18449),
            .in1(N__13783),
            .in2(_gnd_net_),
            .in3(N__13774),
            .lcout(\line_buffer.n3027 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1701_LC_19_13_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1701_LC_19_13_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1701_LC_19_13_3 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1701_LC_19_13_3  (
            .in0(N__15598),
            .in1(N__18476),
            .in2(N__15811),
            .in3(N__15583),
            .lcout(\line_buffer.n3149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i3_LC_19_15_1 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i3_LC_19_15_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i3_LC_19_15_1 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \receive_module.BRAM_ADDR__i3_LC_19_15_1  (
            .in0(N__15574),
            .in1(N__15355),
            .in2(N__16480),
            .in3(N__17872),
            .lcout(RX_ADDR_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16093),
            .ce(),
            .sr(N__15967));
    defparam \receive_module.BRAM_ADDR__i2_LC_19_15_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i2_LC_19_15_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i2_LC_19_15_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \receive_module.BRAM_ADDR__i2_LC_19_15_2  (
            .in0(N__17871),
            .in1(N__15118),
            .in2(N__15334),
            .in3(N__16466),
            .lcout(RX_ADDR_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16093),
            .ce(),
            .sr(N__15967));
    defparam \receive_module.BRAM_ADDR__i1_LC_19_15_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i1_LC_19_15_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i1_LC_19_15_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \receive_module.BRAM_ADDR__i1_LC_19_15_3  (
            .in0(N__15091),
            .in1(N__14872),
            .in2(N__16479),
            .in3(N__17870),
            .lcout(RX_ADDR_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16093),
            .ce(),
            .sr(N__15967));
    defparam \line_buffer.n3149_bdd_4_lut_LC_19_17_3 .C_ON=1'b0;
    defparam \line_buffer.n3149_bdd_4_lut_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3149_bdd_4_lut_LC_19_17_3 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3149_bdd_4_lut_LC_19_17_3  (
            .in0(N__14848),
            .in1(N__15835),
            .in2(N__14833),
            .in3(N__14815),
            .lcout(),
            .ltout(\line_buffer.n3152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i5_LC_19_17_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i5_LC_19_17_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i5_LC_19_17_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i5_LC_19_17_4  (
            .in0(_gnd_net_),
            .in1(N__17686),
            .in2(N__14806),
            .in3(N__15643),
            .lcout(TX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17453),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1580_3_lut_LC_20_9_3 .C_ON=1'b0;
    defparam \line_buffer.i1580_3_lut_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1580_3_lut_LC_20_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i1580_3_lut_LC_20_9_3  (
            .in0(N__18472),
            .in1(N__14791),
            .in2(_gnd_net_),
            .in3(N__14779),
            .lcout(\line_buffer.n3024 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1  (
            .in0(N__15837),
            .in1(N__18250),
            .in2(N__17695),
            .in3(N__14764),
            .lcout(),
            .ltout(\line_buffer.n3131_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i4_LC_20_13_2 .C_ON=1'b0;
    defparam \line_buffer.dout_i4_LC_20_13_2 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i4_LC_20_13_2 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \line_buffer.dout_i4_LC_20_13_2  (
            .in0(N__16981),
            .in1(N__15610),
            .in2(N__14752),
            .in3(N__17693),
            .lcout(TX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__17517),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1602_3_lut_LC_20_13_7 .C_ON=1'b0;
    defparam \line_buffer.i1602_3_lut_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1602_3_lut_LC_20_13_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \line_buffer.i1602_3_lut_LC_20_13_7  (
            .in0(N__18490),
            .in1(N__17014),
            .in2(_gnd_net_),
            .in3(N__16999),
            .lcout(\line_buffer.n3046 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i4_LC_20_14_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i4_LC_20_14_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i4_LC_20_14_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \receive_module.BRAM_ADDR__i4_LC_20_14_5  (
            .in0(N__16753),
            .in1(N__16975),
            .in2(N__16482),
            .in3(N__17873),
            .lcout(RX_ADDR_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16094),
            .ce(),
            .sr(N__15978));
    defparam \receive_module.BRAM_ADDR__i6_LC_20_14_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i6_LC_20_14_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i6_LC_20_14_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \receive_module.BRAM_ADDR__i6_LC_20_14_6  (
            .in0(N__17874),
            .in1(N__16513),
            .in2(N__16729),
            .in3(N__16475),
            .lcout(RX_ADDR_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16094),
            .ce(),
            .sr(N__15978));
    defparam \receive_module.BRAM_ADDR__i10_LC_20_15_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i10_LC_20_15_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i10_LC_20_15_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \receive_module.BRAM_ADDR__i10_LC_20_15_5  (
            .in0(N__16150),
            .in1(N__16492),
            .in2(N__16483),
            .in3(N__17875),
            .lcout(RX_ADDR_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16097),
            .ce(),
            .sr(N__15968));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1706_LC_20_17_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1706_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_1706_LC_20_17_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_1706_LC_20_17_0  (
            .in0(N__18488),
            .in1(N__15904),
            .in2(N__15838),
            .in3(N__15892),
            .lcout(),
            .ltout(\line_buffer.n3155_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3155_bdd_4_lut_LC_20_17_1 .C_ON=1'b0;
    defparam \line_buffer.n3155_bdd_4_lut_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3155_bdd_4_lut_LC_20_17_1 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.n3155_bdd_4_lut_LC_20_17_1  (
            .in0(N__15874),
            .in1(N__15856),
            .in2(N__15841),
            .in3(N__15834),
            .lcout(\line_buffer.n3158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1601_3_lut_LC_20_19_0 .C_ON=1'b0;
    defparam \line_buffer.i1601_3_lut_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1601_3_lut_LC_20_19_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i1601_3_lut_LC_20_19_0  (
            .in0(N__15637),
            .in1(N__15622),
            .in2(_gnd_net_),
            .in3(N__18473),
            .lcout(\line_buffer.n3045 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1581_3_lut_LC_21_13_0 .C_ON=1'b0;
    defparam \line_buffer.i1581_3_lut_LC_21_13_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1581_3_lut_LC_21_13_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i1581_3_lut_LC_21_13_0  (
            .in0(N__18489),
            .in1(N__18286),
            .in2(_gnd_net_),
            .in3(N__18271),
            .lcout(\line_buffer.n3025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_21_13_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_21_13_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_21_13_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_21_13_5  (
            .in0(N__18138),
            .in1(N__18047),
            .in2(N__17974),
            .in3(N__17857),
            .lcout(\line_buffer.n729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_22_13_2 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_22_13_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_22_13_2  (
            .in0(N__18135),
            .in1(N__18054),
            .in2(N__17973),
            .in3(N__17877),
            .lcout(\line_buffer.n697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_22_17_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_22_17_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_22_17_5  (
            .in0(N__18136),
            .in1(N__18055),
            .in2(N__17975),
            .in3(N__17876),
            .lcout(\line_buffer.n633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // main
