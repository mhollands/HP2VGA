// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 15 2018 02:00:41

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "main" view "INTERFACE"

module main (
    TVP_VIDEO,
    ADV_B,
    ADV_G,
    ADV_R,
    DEBUG,
    TVP_CLK,
    ADV_CLK,
    TVP_HSYNC,
    ADV_HSYNC,
    TVP_VSYNC,
    ADV_VSYNC,
    ADV_BLANK_N,
    LED,
    ADV_SYNC_N);

    input [9:0] TVP_VIDEO;
    output [7:0] ADV_B;
    output [7:0] ADV_G;
    output [7:0] ADV_R;
    inout [7:0] DEBUG;
    input TVP_CLK;
    output ADV_CLK;
    input TVP_HSYNC;
    output ADV_HSYNC;
    input TVP_VSYNC;
    output ADV_VSYNC;
    output ADV_BLANK_N;
    output LED;
    output ADV_SYNC_N;

    wire N__23675;
    wire N__23674;
    wire N__23673;
    wire N__23664;
    wire N__23663;
    wire N__23662;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23646;
    wire N__23645;
    wire N__23644;
    wire N__23637;
    wire N__23636;
    wire N__23635;
    wire N__23628;
    wire N__23627;
    wire N__23626;
    wire N__23619;
    wire N__23618;
    wire N__23617;
    wire N__23610;
    wire N__23609;
    wire N__23608;
    wire N__23601;
    wire N__23600;
    wire N__23599;
    wire N__23592;
    wire N__23591;
    wire N__23590;
    wire N__23583;
    wire N__23582;
    wire N__23581;
    wire N__23574;
    wire N__23573;
    wire N__23572;
    wire N__23565;
    wire N__23564;
    wire N__23563;
    wire N__23556;
    wire N__23555;
    wire N__23554;
    wire N__23547;
    wire N__23546;
    wire N__23545;
    wire N__23538;
    wire N__23537;
    wire N__23536;
    wire N__23529;
    wire N__23528;
    wire N__23527;
    wire N__23520;
    wire N__23519;
    wire N__23518;
    wire N__23511;
    wire N__23510;
    wire N__23509;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23493;
    wire N__23492;
    wire N__23491;
    wire N__23484;
    wire N__23483;
    wire N__23482;
    wire N__23475;
    wire N__23474;
    wire N__23473;
    wire N__23466;
    wire N__23465;
    wire N__23464;
    wire N__23457;
    wire N__23456;
    wire N__23455;
    wire N__23448;
    wire N__23447;
    wire N__23446;
    wire N__23439;
    wire N__23438;
    wire N__23437;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23421;
    wire N__23420;
    wire N__23419;
    wire N__23412;
    wire N__23411;
    wire N__23410;
    wire N__23403;
    wire N__23402;
    wire N__23401;
    wire N__23394;
    wire N__23393;
    wire N__23392;
    wire N__23385;
    wire N__23384;
    wire N__23383;
    wire N__23376;
    wire N__23375;
    wire N__23374;
    wire N__23367;
    wire N__23366;
    wire N__23365;
    wire N__23358;
    wire N__23357;
    wire N__23356;
    wire N__23349;
    wire N__23348;
    wire N__23347;
    wire N__23340;
    wire N__23339;
    wire N__23338;
    wire N__23331;
    wire N__23330;
    wire N__23329;
    wire N__23322;
    wire N__23321;
    wire N__23320;
    wire N__23313;
    wire N__23312;
    wire N__23311;
    wire N__23304;
    wire N__23303;
    wire N__23302;
    wire N__23295;
    wire N__23294;
    wire N__23293;
    wire N__23286;
    wire N__23285;
    wire N__23284;
    wire N__23277;
    wire N__23276;
    wire N__23275;
    wire N__23268;
    wire N__23267;
    wire N__23266;
    wire N__23259;
    wire N__23258;
    wire N__23257;
    wire N__23250;
    wire N__23249;
    wire N__23248;
    wire N__23241;
    wire N__23240;
    wire N__23239;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23143;
    wire N__23142;
    wire N__23141;
    wire N__23138;
    wire N__23137;
    wire N__23136;
    wire N__23135;
    wire N__23134;
    wire N__23133;
    wire N__23132;
    wire N__23131;
    wire N__23130;
    wire N__23129;
    wire N__23126;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23118;
    wire N__23117;
    wire N__23114;
    wire N__23109;
    wire N__23108;
    wire N__23107;
    wire N__23106;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23094;
    wire N__23093;
    wire N__23092;
    wire N__23091;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23025;
    wire N__23016;
    wire N__23013;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22986;
    wire N__22981;
    wire N__22970;
    wire N__22965;
    wire N__22960;
    wire N__22955;
    wire N__22946;
    wire N__22943;
    wire N__22934;
    wire N__22933;
    wire N__22932;
    wire N__22931;
    wire N__22930;
    wire N__22929;
    wire N__22928;
    wire N__22927;
    wire N__22926;
    wire N__22925;
    wire N__22922;
    wire N__22921;
    wire N__22920;
    wire N__22919;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22908;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22897;
    wire N__22896;
    wire N__22893;
    wire N__22892;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22873;
    wire N__22872;
    wire N__22867;
    wire N__22866;
    wire N__22865;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22850;
    wire N__22847;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22832;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22807;
    wire N__22802;
    wire N__22795;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22774;
    wire N__22765;
    wire N__22758;
    wire N__22753;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22686;
    wire N__22685;
    wire N__22684;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22672;
    wire N__22671;
    wire N__22668;
    wire N__22667;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22653;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22645;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22621;
    wire N__22620;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22608;
    wire N__22607;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22592;
    wire N__22591;
    wire N__22590;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22575;
    wire N__22574;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22557;
    wire N__22556;
    wire N__22555;
    wire N__22554;
    wire N__22551;
    wire N__22546;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22534;
    wire N__22533;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22516;
    wire N__22515;
    wire N__22512;
    wire N__22509;
    wire N__22508;
    wire N__22507;
    wire N__22506;
    wire N__22503;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22471;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22449;
    wire N__22446;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22432;
    wire N__22427;
    wire N__22422;
    wire N__22419;
    wire N__22414;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22374;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22159;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22151;
    wire N__22150;
    wire N__22149;
    wire N__22146;
    wire N__22145;
    wire N__22144;
    wire N__22143;
    wire N__22142;
    wire N__22141;
    wire N__22140;
    wire N__22139;
    wire N__22138;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22124;
    wire N__22123;
    wire N__22120;
    wire N__22119;
    wire N__22118;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22104;
    wire N__22103;
    wire N__22100;
    wire N__22099;
    wire N__22096;
    wire N__22095;
    wire N__22092;
    wire N__22091;
    wire N__22090;
    wire N__22089;
    wire N__22088;
    wire N__22087;
    wire N__22086;
    wire N__22085;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22077;
    wire N__22074;
    wire N__22073;
    wire N__22072;
    wire N__22071;
    wire N__22070;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22053;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22038;
    wire N__22037;
    wire N__22032;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21987;
    wire N__21984;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21959;
    wire N__21958;
    wire N__21957;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21943;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21926;
    wire N__21925;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21893;
    wire N__21888;
    wire N__21885;
    wire N__21880;
    wire N__21877;
    wire N__21876;
    wire N__21875;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21842;
    wire N__21839;
    wire N__21832;
    wire N__21829;
    wire N__21828;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21817;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21809;
    wire N__21808;
    wire N__21805;
    wire N__21804;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21786;
    wire N__21783;
    wire N__21782;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21765;
    wire N__21762;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21742;
    wire N__21735;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21723;
    wire N__21720;
    wire N__21715;
    wire N__21708;
    wire N__21703;
    wire N__21698;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21686;
    wire N__21685;
    wire N__21684;
    wire N__21683;
    wire N__21682;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21667;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21628;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21604;
    wire N__21593;
    wire N__21590;
    wire N__21585;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21559;
    wire N__21558;
    wire N__21557;
    wire N__21554;
    wire N__21553;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21518;
    wire N__21513;
    wire N__21510;
    wire N__21509;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21491;
    wire N__21490;
    wire N__21487;
    wire N__21480;
    wire N__21479;
    wire N__21476;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21447;
    wire N__21446;
    wire N__21439;
    wire N__21434;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21416;
    wire N__21413;
    wire N__21408;
    wire N__21405;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21371;
    wire N__21366;
    wire N__21361;
    wire N__21356;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21330;
    wire N__21325;
    wire N__21322;
    wire N__21317;
    wire N__21308;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21295;
    wire N__21292;
    wire N__21291;
    wire N__21290;
    wire N__21289;
    wire N__21288;
    wire N__21285;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21277;
    wire N__21276;
    wire N__21273;
    wire N__21272;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21261;
    wire N__21258;
    wire N__21257;
    wire N__21254;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21242;
    wire N__21235;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21176;
    wire N__21173;
    wire N__21168;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21093;
    wire N__21088;
    wire N__21083;
    wire N__21080;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21050;
    wire N__21047;
    wire N__21046;
    wire N__21045;
    wire N__21044;
    wire N__21043;
    wire N__21042;
    wire N__21041;
    wire N__21040;
    wire N__21039;
    wire N__21036;
    wire N__21035;
    wire N__21034;
    wire N__21033;
    wire N__21032;
    wire N__21031;
    wire N__21030;
    wire N__21029;
    wire N__21028;
    wire N__21027;
    wire N__21026;
    wire N__21025;
    wire N__21024;
    wire N__21023;
    wire N__21022;
    wire N__21021;
    wire N__21020;
    wire N__21019;
    wire N__21018;
    wire N__21017;
    wire N__21016;
    wire N__21015;
    wire N__21014;
    wire N__21013;
    wire N__21012;
    wire N__21011;
    wire N__21010;
    wire N__21009;
    wire N__21008;
    wire N__21007;
    wire N__21006;
    wire N__21005;
    wire N__21004;
    wire N__21003;
    wire N__21002;
    wire N__21001;
    wire N__21000;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20732;
    wire N__20729;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20717;
    wire N__20714;
    wire N__20713;
    wire N__20712;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20701;
    wire N__20700;
    wire N__20699;
    wire N__20698;
    wire N__20697;
    wire N__20696;
    wire N__20695;
    wire N__20694;
    wire N__20693;
    wire N__20692;
    wire N__20691;
    wire N__20690;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20684;
    wire N__20683;
    wire N__20682;
    wire N__20681;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20666;
    wire N__20665;
    wire N__20662;
    wire N__20661;
    wire N__20660;
    wire N__20657;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20620;
    wire N__20619;
    wire N__20618;
    wire N__20617;
    wire N__20614;
    wire N__20613;
    wire N__20610;
    wire N__20609;
    wire N__20606;
    wire N__20605;
    wire N__20602;
    wire N__20601;
    wire N__20600;
    wire N__20599;
    wire N__20598;
    wire N__20593;
    wire N__20588;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20577;
    wire N__20574;
    wire N__20573;
    wire N__20572;
    wire N__20569;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20557;
    wire N__20554;
    wire N__20545;
    wire N__20540;
    wire N__20537;
    wire N__20532;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20513;
    wire N__20512;
    wire N__20509;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20495;
    wire N__20492;
    wire N__20491;
    wire N__20490;
    wire N__20489;
    wire N__20486;
    wire N__20481;
    wire N__20476;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20431;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20395;
    wire N__20392;
    wire N__20385;
    wire N__20384;
    wire N__20383;
    wire N__20378;
    wire N__20369;
    wire N__20368;
    wire N__20367;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20349;
    wire N__20342;
    wire N__20337;
    wire N__20328;
    wire N__20315;
    wire N__20310;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20291;
    wire N__20284;
    wire N__20277;
    wire N__20270;
    wire N__20255;
    wire N__20254;
    wire N__20253;
    wire N__20252;
    wire N__20251;
    wire N__20250;
    wire N__20249;
    wire N__20246;
    wire N__20241;
    wire N__20240;
    wire N__20239;
    wire N__20238;
    wire N__20237;
    wire N__20236;
    wire N__20235;
    wire N__20234;
    wire N__20233;
    wire N__20232;
    wire N__20229;
    wire N__20222;
    wire N__20217;
    wire N__20212;
    wire N__20207;
    wire N__20206;
    wire N__20197;
    wire N__20196;
    wire N__20195;
    wire N__20194;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20180;
    wire N__20179;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20160;
    wire N__20157;
    wire N__20152;
    wire N__20147;
    wire N__20136;
    wire N__20129;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19913;
    wire N__19912;
    wire N__19907;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19841;
    wire N__19838;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19826;
    wire N__19823;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19811;
    wire N__19808;
    wire N__19807;
    wire N__19806;
    wire N__19803;
    wire N__19798;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19768;
    wire N__19765;
    wire N__19764;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19739;
    wire N__19738;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19730;
    wire N__19729;
    wire N__19728;
    wire N__19727;
    wire N__19724;
    wire N__19723;
    wire N__19722;
    wire N__19721;
    wire N__19716;
    wire N__19709;
    wire N__19708;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19693;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19674;
    wire N__19669;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19636;
    wire N__19635;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19623;
    wire N__19616;
    wire N__19615;
    wire N__19610;
    wire N__19609;
    wire N__19608;
    wire N__19607;
    wire N__19606;
    wire N__19605;
    wire N__19602;
    wire N__19597;
    wire N__19594;
    wire N__19593;
    wire N__19592;
    wire N__19591;
    wire N__19590;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19576;
    wire N__19569;
    wire N__19568;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19550;
    wire N__19549;
    wire N__19548;
    wire N__19547;
    wire N__19546;
    wire N__19545;
    wire N__19544;
    wire N__19543;
    wire N__19542;
    wire N__19537;
    wire N__19530;
    wire N__19525;
    wire N__19516;
    wire N__19507;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19478;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19262;
    wire N__19259;
    wire N__19258;
    wire N__19257;
    wire N__19254;
    wire N__19253;
    wire N__19252;
    wire N__19251;
    wire N__19250;
    wire N__19249;
    wire N__19246;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19228;
    wire N__19227;
    wire N__19226;
    wire N__19223;
    wire N__19222;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19207;
    wire N__19202;
    wire N__19197;
    wire N__19194;
    wire N__19189;
    wire N__19188;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19172;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19150;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19132;
    wire N__19129;
    wire N__19128;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18730;
    wire N__18727;
    wire N__18726;
    wire N__18725;
    wire N__18724;
    wire N__18721;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18713;
    wire N__18712;
    wire N__18709;
    wire N__18708;
    wire N__18707;
    wire N__18704;
    wire N__18703;
    wire N__18702;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18694;
    wire N__18693;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18613;
    wire N__18610;
    wire N__18603;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18584;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18459;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18438;
    wire N__18435;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17983;
    wire N__17982;
    wire N__17981;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17970;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17962;
    wire N__17959;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17943;
    wire N__17940;
    wire N__17939;
    wire N__17936;
    wire N__17931;
    wire N__17928;
    wire N__17925;
    wire N__17922;
    wire N__17919;
    wire N__17914;
    wire N__17913;
    wire N__17910;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17839;
    wire N__17838;
    wire N__17837;
    wire N__17836;
    wire N__17835;
    wire N__17834;
    wire N__17833;
    wire N__17832;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17808;
    wire N__17805;
    wire N__17802;
    wire N__17801;
    wire N__17792;
    wire N__17785;
    wire N__17774;
    wire N__17773;
    wire N__17772;
    wire N__17771;
    wire N__17770;
    wire N__17767;
    wire N__17762;
    wire N__17759;
    wire N__17758;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17731;
    wire N__17728;
    wire N__17723;
    wire N__17720;
    wire N__17715;
    wire N__17710;
    wire N__17707;
    wire N__17702;
    wire N__17699;
    wire N__17698;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17690;
    wire N__17687;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17675;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17661;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17645;
    wire N__17644;
    wire N__17643;
    wire N__17640;
    wire N__17639;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17601;
    wire N__17594;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17501;
    wire N__17498;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17464;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17368;
    wire N__17365;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17348;
    wire N__17347;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17317;
    wire N__17316;
    wire N__17315;
    wire N__17312;
    wire N__17307;
    wire N__17304;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17279;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16846;
    wire N__16843;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16721;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16700;
    wire N__16697;
    wire N__16692;
    wire N__16689;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16669;
    wire N__16668;
    wire N__16667;
    wire N__16664;
    wire N__16659;
    wire N__16656;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16621;
    wire N__16620;
    wire N__16619;
    wire N__16616;
    wire N__16611;
    wire N__16608;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16577;
    wire N__16576;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16568;
    wire N__16565;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16544;
    wire N__16543;
    wire N__16540;
    wire N__16539;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16471;
    wire N__16470;
    wire N__16467;
    wire N__16464;
    wire N__16463;
    wire N__16460;
    wire N__16455;
    wire N__16452;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16435;
    wire N__16432;
    wire N__16431;
    wire N__16428;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16393;
    wire N__16390;
    wire N__16389;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16377;
    wire N__16370;
    wire N__16367;
    wire N__16366;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16349;
    wire N__16346;
    wire N__16345;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16328;
    wire N__16325;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16313;
    wire N__16310;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16298;
    wire N__16295;
    wire N__16294;
    wire N__16293;
    wire N__16290;
    wire N__16285;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16265;
    wire N__16262;
    wire N__16261;
    wire N__16260;
    wire N__16259;
    wire N__16258;
    wire N__16255;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16221;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16213;
    wire N__16210;
    wire N__16209;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16194;
    wire N__16189;
    wire N__16186;
    wire N__16175;
    wire N__16174;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15976;
    wire N__15975;
    wire N__15972;
    wire N__15969;
    wire N__15966;
    wire N__15963;
    wire N__15960;
    wire N__15957;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15939;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15916;
    wire N__15915;
    wire N__15914;
    wire N__15913;
    wire N__15912;
    wire N__15911;
    wire N__15910;
    wire N__15909;
    wire N__15900;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15879;
    wire N__15876;
    wire N__15871;
    wire N__15868;
    wire N__15863;
    wire N__15860;
    wire N__15859;
    wire N__15856;
    wire N__15855;
    wire N__15854;
    wire N__15853;
    wire N__15848;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15840;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15829;
    wire N__15820;
    wire N__15817;
    wire N__15814;
    wire N__15811;
    wire N__15808;
    wire N__15805;
    wire N__15802;
    wire N__15797;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15766;
    wire N__15765;
    wire N__15764;
    wire N__15761;
    wire N__15760;
    wire N__15759;
    wire N__15756;
    wire N__15753;
    wire N__15752;
    wire N__15751;
    wire N__15748;
    wire N__15747;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15728;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15708;
    wire N__15701;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15665;
    wire N__15662;
    wire N__15661;
    wire N__15660;
    wire N__15659;
    wire N__15656;
    wire N__15649;
    wire N__15644;
    wire N__15641;
    wire N__15640;
    wire N__15639;
    wire N__15638;
    wire N__15635;
    wire N__15628;
    wire N__15623;
    wire N__15620;
    wire N__15619;
    wire N__15618;
    wire N__15615;
    wire N__15614;
    wire N__15611;
    wire N__15604;
    wire N__15599;
    wire N__15596;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15496;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15388;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15360;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15337;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15124;
    wire N__15121;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15113;
    wire N__15110;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15096;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14871;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14853;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14611;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14601;
    wire N__14598;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14382;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14364;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14130;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14112;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13899;
    wire N__13896;
    wire N__13893;
    wire N__13890;
    wire N__13887;
    wire N__13884;
    wire N__13881;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13837;
    wire N__13834;
    wire N__13831;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13657;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13642;
    wire N__13639;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13619;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13582;
    wire N__13579;
    wire N__13576;
    wire N__13571;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13559;
    wire N__13558;
    wire N__13555;
    wire N__13552;
    wire N__13547;
    wire N__13546;
    wire N__13543;
    wire N__13540;
    wire N__13535;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13523;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13498;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13468;
    wire N__13465;
    wire N__13462;
    wire N__13459;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13447;
    wire N__13444;
    wire N__13441;
    wire N__13438;
    wire N__13435;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13417;
    wire N__13414;
    wire N__13411;
    wire N__13408;
    wire N__13405;
    wire N__13402;
    wire N__13399;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13384;
    wire N__13381;
    wire N__13378;
    wire N__13375;
    wire N__13372;
    wire N__13369;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13357;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13324;
    wire N__13321;
    wire N__13318;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13291;
    wire N__13288;
    wire N__13285;
    wire N__13282;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13270;
    wire N__13269;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13219;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13192;
    wire N__13189;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13108;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13054;
    wire N__13051;
    wire N__13048;
    wire N__13045;
    wire N__13042;
    wire N__13039;
    wire N__13036;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13010;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12993;
    wire N__12990;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12965;
    wire N__12962;
    wire N__12959;
    wire N__12956;
    wire N__12955;
    wire N__12954;
    wire N__12953;
    wire N__12948;
    wire N__12943;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12931;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12916;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12880;
    wire N__12879;
    wire N__12878;
    wire N__12875;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12867;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12822;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12694;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12637;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12584;
    wire N__12581;
    wire N__12580;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12546;
    wire N__12543;
    wire N__12540;
    wire N__12535;
    wire N__12532;
    wire N__12529;
    wire N__12524;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12475;
    wire N__12470;
    wire N__12469;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12424;
    wire N__12421;
    wire N__12416;
    wire N__12413;
    wire N__12412;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12358;
    wire N__12353;
    wire N__12350;
    wire N__12349;
    wire N__12346;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12049;
    wire N__12046;
    wire N__12045;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12023;
    wire N__12020;
    wire N__12019;
    wire N__12018;
    wire N__12017;
    wire N__12016;
    wire N__12013;
    wire N__12012;
    wire N__12011;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11975;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11920;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11863;
    wire N__11860;
    wire N__11857;
    wire N__11854;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11767;
    wire N__11764;
    wire N__11761;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11683;
    wire N__11680;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11449;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11351;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11320;
    wire N__11319;
    wire N__11318;
    wire N__11317;
    wire N__11316;
    wire N__11315;
    wire N__11314;
    wire N__11313;
    wire N__11312;
    wire N__11311;
    wire N__11310;
    wire N__11309;
    wire N__11308;
    wire N__11305;
    wire N__11304;
    wire N__11303;
    wire N__11302;
    wire N__11301;
    wire N__11300;
    wire N__11299;
    wire N__11298;
    wire N__11287;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11259;
    wire N__11250;
    wire N__11245;
    wire N__11234;
    wire N__11231;
    wire N__11230;
    wire N__11227;
    wire N__11226;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11204;
    wire N__11201;
    wire N__11200;
    wire N__11199;
    wire N__11196;
    wire N__11193;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11177;
    wire N__11174;
    wire N__11173;
    wire N__11172;
    wire N__11169;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11134;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11118;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11104;
    wire N__11101;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11093;
    wire N__11090;
    wire N__11085;
    wire N__11082;
    wire N__11075;
    wire N__11074;
    wire N__11071;
    wire N__11070;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11058;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11007;
    wire N__11004;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10979;
    wire N__10978;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10970;
    wire N__10967;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10951;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10918;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10831;
    wire N__10828;
    wire N__10825;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10814;
    wire N__10811;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10774;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10766;
    wire N__10763;
    wire N__10758;
    wire N__10755;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10738;
    wire N__10733;
    wire N__10732;
    wire N__10731;
    wire N__10730;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10700;
    wire N__10699;
    wire N__10698;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10690;
    wire N__10687;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10606;
    wire N__10603;
    wire N__10600;
    wire N__10597;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10525;
    wire N__10522;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10345;
    wire N__10342;
    wire N__10339;
    wire N__10336;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10205;
    wire N__10204;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10183;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10166;
    wire N__10163;
    wire N__10162;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10112;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10100;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10075;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10009;
    wire N__10006;
    wire N__10005;
    wire N__10002;
    wire N__9997;
    wire N__9992;
    wire N__9991;
    wire N__9990;
    wire N__9987;
    wire N__9982;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9967;
    wire N__9966;
    wire N__9965;
    wire N__9962;
    wire N__9957;
    wire N__9954;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9940;
    wire N__9939;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9907;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9861;
    wire N__9856;
    wire N__9853;
    wire N__9852;
    wire N__9847;
    wire N__9844;
    wire N__9841;
    wire N__9838;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9815;
    wire N__9812;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9553;
    wire N__9552;
    wire N__9549;
    wire N__9544;
    wire N__9539;
    wire N__9538;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9507;
    wire N__9502;
    wire N__9499;
    wire N__9498;
    wire N__9493;
    wire N__9490;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9458;
    wire N__9455;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9439;
    wire N__9436;
    wire N__9433;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8759;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8751;
    wire N__8746;
    wire N__8743;
    wire N__8738;
    wire N__8737;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8722;
    wire N__8719;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8688;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8671;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8638;
    wire N__8637;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8626;
    wire N__8623;
    wire N__8616;
    wire N__8613;
    wire N__8612;
    wire N__8609;
    wire N__8604;
    wire N__8601;
    wire N__8600;
    wire N__8599;
    wire N__8596;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8528;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8520;
    wire N__8515;
    wire N__8512;
    wire N__8507;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8499;
    wire N__8494;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8449;
    wire N__8446;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8426;
    wire N__8423;
    wire N__8422;
    wire N__8421;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8381;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8343;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8322;
    wire N__8319;
    wire N__8312;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8291;
    wire N__8288;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8276;
    wire N__8271;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8252;
    wire N__8249;
    wire N__8244;
    wire N__8239;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8210;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8186;
    wire N__8181;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8167;
    wire N__8162;
    wire N__8161;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8142;
    wire N__8137;
    wire N__8136;
    wire N__8133;
    wire N__8130;
    wire N__8127;
    wire N__8124;
    wire N__8119;
    wire N__8116;
    wire N__8113;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8101;
    wire N__8100;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8092;
    wire N__8089;
    wire N__8088;
    wire N__8085;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7969;
    wire N__7966;
    wire N__7963;
    wire N__7962;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7948;
    wire N__7947;
    wire N__7942;
    wire N__7939;
    wire N__7938;
    wire N__7933;
    wire N__7930;
    wire N__7929;
    wire N__7924;
    wire N__7921;
    wire N__7920;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7876;
    wire TVP_VIDEO_c_3;
    wire VCCG0;
    wire TVP_VIDEO_c_5;
    wire TVP_VIDEO_c_4;
    wire GNDG0;
    wire TVP_VIDEO_c_7;
    wire TVP_VIDEO_c_6;
    wire TVP_VIDEO_c_8;
    wire TVP_VIDEO_c_9;
    wire TVP_VIDEO_c_2;
    wire \transmit_module.Y_DELTA_PATTERN_55 ;
    wire \transmit_module.Y_DELTA_PATTERN_54 ;
    wire \transmit_module.Y_DELTA_PATTERN_53 ;
    wire \transmit_module.Y_DELTA_PATTERN_52 ;
    wire \transmit_module.Y_DELTA_PATTERN_14 ;
    wire \transmit_module.Y_DELTA_PATTERN_15 ;
    wire \transmit_module.Y_DELTA_PATTERN_16 ;
    wire \transmit_module.Y_DELTA_PATTERN_17 ;
    wire \transmit_module.Y_DELTA_PATTERN_19 ;
    wire \transmit_module.Y_DELTA_PATTERN_18 ;
    wire \transmit_module.Y_DELTA_PATTERN_71 ;
    wire \transmit_module.Y_DELTA_PATTERN_70 ;
    wire \transmit_module.Y_DELTA_PATTERN_60 ;
    wire \transmit_module.Y_DELTA_PATTERN_59 ;
    wire \transmit_module.Y_DELTA_PATTERN_42 ;
    wire \transmit_module.Y_DELTA_PATTERN_41 ;
    wire \transmit_module.Y_DELTA_PATTERN_69 ;
    wire \transmit_module.Y_DELTA_PATTERN_56 ;
    wire \transmit_module.Y_DELTA_PATTERN_58 ;
    wire \transmit_module.Y_DELTA_PATTERN_57 ;
    wire \transmit_module.Y_DELTA_PATTERN_61 ;
    wire \line_buffer.n639 ;
    wire \line_buffer.n631 ;
    wire \transmit_module.X_DELTA_PATTERN_11 ;
    wire \transmit_module.X_DELTA_PATTERN_10 ;
    wire \transmit_module.Y_DELTA_PATTERN_24 ;
    wire \transmit_module.Y_DELTA_PATTERN_6 ;
    wire \transmit_module.Y_DELTA_PATTERN_20 ;
    wire \transmit_module.Y_DELTA_PATTERN_21 ;
    wire \transmit_module.Y_DELTA_PATTERN_23 ;
    wire \transmit_module.Y_DELTA_PATTERN_22 ;
    wire \transmit_module.Y_DELTA_PATTERN_5 ;
    wire \transmit_module.Y_DELTA_PATTERN_1 ;
    wire \transmit_module.Y_DELTA_PATTERN_4 ;
    wire \transmit_module.Y_DELTA_PATTERN_45 ;
    wire \transmit_module.Y_DELTA_PATTERN_77 ;
    wire \transmit_module.Y_DELTA_PATTERN_3 ;
    wire \transmit_module.Y_DELTA_PATTERN_2 ;
    wire \transmit_module.Y_DELTA_PATTERN_46 ;
    wire \transmit_module.Y_DELTA_PATTERN_78 ;
    wire \transmit_module.Y_DELTA_PATTERN_68 ;
    wire \transmit_module.Y_DELTA_PATTERN_79 ;
    wire \transmit_module.Y_DELTA_PATTERN_48 ;
    wire \transmit_module.Y_DELTA_PATTERN_47 ;
    wire \transmit_module.Y_DELTA_PATTERN_67 ;
    wire \transmit_module.Y_DELTA_PATTERN_82 ;
    wire \transmit_module.Y_DELTA_PATTERN_44 ;
    wire \transmit_module.Y_DELTA_PATTERN_43 ;
    wire \transmit_module.Y_DELTA_PATTERN_81 ;
    wire \transmit_module.Y_DELTA_PATTERN_80 ;
    wire \transmit_module.Y_DELTA_PATTERN_66 ;
    wire \transmit_module.Y_DELTA_PATTERN_76 ;
    wire \transmit_module.Y_DELTA_PATTERN_75 ;
    wire \transmit_module.Y_DELTA_PATTERN_51 ;
    wire \transmit_module.Y_DELTA_PATTERN_63 ;
    wire \transmit_module.Y_DELTA_PATTERN_62 ;
    wire \transmit_module.Y_DELTA_PATTERN_74 ;
    wire \transmit_module.Y_DELTA_PATTERN_50 ;
    wire \transmit_module.Y_DELTA_PATTERN_49 ;
    wire \transmit_module.Y_DELTA_PATTERN_65 ;
    wire \transmit_module.Y_DELTA_PATTERN_64 ;
    wire \transmit_module.X_DELTA_PATTERN_12 ;
    wire \transmit_module.X_DELTA_PATTERN_13 ;
    wire old_HS;
    wire bfn_11_9_0_;
    wire \receive_module.rx_counter.n3349 ;
    wire \receive_module.rx_counter.n3350 ;
    wire \receive_module.rx_counter.n3351 ;
    wire \receive_module.rx_counter.n3352 ;
    wire \receive_module.rx_counter.n3353 ;
    wire \receive_module.rx_counter.n3354 ;
    wire \receive_module.rx_counter.n3355 ;
    wire \receive_module.rx_counter.n3356 ;
    wire bfn_11_10_0_;
    wire n2057;
    wire \transmit_module.Y_DELTA_PATTERN_26 ;
    wire \transmit_module.Y_DELTA_PATTERN_25 ;
    wire \transmit_module.Y_DELTA_PATTERN_7 ;
    wire \transmit_module.Y_DELTA_PATTERN_27 ;
    wire \transmit_module.Y_DELTA_PATTERN_10 ;
    wire \transmit_module.Y_DELTA_PATTERN_13 ;
    wire \transmit_module.Y_DELTA_PATTERN_9 ;
    wire \transmit_module.Y_DELTA_PATTERN_8 ;
    wire \transmit_module.Y_DELTA_PATTERN_12 ;
    wire \transmit_module.Y_DELTA_PATTERN_11 ;
    wire \transmit_module.Y_DELTA_PATTERN_83 ;
    wire \transmit_module.Y_DELTA_PATTERN_84 ;
    wire \transmit_module.Y_DELTA_PATTERN_95 ;
    wire \transmit_module.Y_DELTA_PATTERN_94 ;
    wire \transmit_module.Y_DELTA_PATTERN_93 ;
    wire \transmit_module.Y_DELTA_PATTERN_85 ;
    wire \transmit_module.Y_DELTA_PATTERN_86 ;
    wire \transmit_module.Y_DELTA_PATTERN_92 ;
    wire \transmit_module.Y_DELTA_PATTERN_91 ;
    wire bfn_11_15_0_;
    wire \transmit_module.video_signal_controller.n3377 ;
    wire \transmit_module.video_signal_controller.n3378 ;
    wire \transmit_module.video_signal_controller.n3379 ;
    wire \transmit_module.video_signal_controller.n3380 ;
    wire \transmit_module.video_signal_controller.n3381 ;
    wire \transmit_module.video_signal_controller.n3382 ;
    wire \transmit_module.video_signal_controller.n3383 ;
    wire \transmit_module.video_signal_controller.n3384 ;
    wire bfn_11_16_0_;
    wire \transmit_module.video_signal_controller.n3385 ;
    wire \transmit_module.video_signal_controller.n3386 ;
    wire \transmit_module.Y_DELTA_PATTERN_28 ;
    wire \transmit_module.Y_DELTA_PATTERN_29 ;
    wire \transmit_module.Y_DELTA_PATTERN_30 ;
    wire \transmit_module.Y_DELTA_PATTERN_31 ;
    wire \transmit_module.Y_DELTA_PATTERN_73 ;
    wire \transmit_module.Y_DELTA_PATTERN_72 ;
    wire n22;
    wire \transmit_module.X_DELTA_PATTERN_15 ;
    wire \transmit_module.X_DELTA_PATTERN_14 ;
    wire \line_buffer.n630 ;
    wire \line_buffer.n638 ;
    wire \receive_module.rx_counter.Y_6 ;
    wire \receive_module.rx_counter.Y_5 ;
    wire \receive_module.rx_counter.n3619_cascade_ ;
    wire \line_buffer.n642 ;
    wire \line_buffer.n578 ;
    wire \receive_module.rx_counter.n14_cascade_ ;
    wire \receive_module.rx_counter.Y_8 ;
    wire \receive_module.rx_counter.Y_7 ;
    wire \receive_module.rx_counter.n15_cascade_ ;
    wire \receive_module.rx_counter.n3861 ;
    wire \receive_module.rx_counter.Y_0 ;
    wire \receive_module.rx_counter.n10_adj_570 ;
    wire \receive_module.rx_counter.Y_2 ;
    wire \line_buffer.n610 ;
    wire \line_buffer.n512 ;
    wire \transmit_module.Y_DELTA_PATTERN_99 ;
    wire \transmit_module.Y_DELTA_PATTERN_90 ;
    wire \transmit_module.Y_DELTA_PATTERN_87 ;
    wire \transmit_module.Y_DELTA_PATTERN_89 ;
    wire \transmit_module.Y_DELTA_PATTERN_88 ;
    wire \transmit_module.Y_DELTA_PATTERN_98 ;
    wire \transmit_module.Y_DELTA_PATTERN_97 ;
    wire \transmit_module.Y_DELTA_PATTERN_96 ;
    wire \transmit_module.video_signal_controller.VGA_X_1 ;
    wire \transmit_module.video_signal_controller.VGA_X_2 ;
    wire \transmit_module.video_signal_controller.VGA_X_0 ;
    wire \transmit_module.video_signal_controller.n8_adj_569_cascade_ ;
    wire \transmit_module.video_signal_controller.n3029_cascade_ ;
    wire \transmit_module.video_signal_controller.n3857_cascade_ ;
    wire \transmit_module.n2125 ;
    wire \transmit_module.n3859_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_7 ;
    wire \transmit_module.video_signal_controller.n4_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_6 ;
    wire \transmit_module.video_signal_controller.n23_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_10 ;
    wire \transmit_module.video_signal_controller.VGA_X_9 ;
    wire \transmit_module.n214 ;
    wire \transmit_module.n182 ;
    wire \transmit_module.n214_cascade_ ;
    wire n20;
    wire \transmit_module.n215_cascade_ ;
    wire n23;
    wire \transmit_module.n183 ;
    wire \transmit_module.n215 ;
    wire \transmit_module.n212 ;
    wire \transmit_module.n180 ;
    wire \transmit_module.n212_cascade_ ;
    wire \transmit_module.X_DELTA_PATTERN_9 ;
    wire \transmit_module.X_DELTA_PATTERN_8 ;
    wire \transmit_module.X_DELTA_PATTERN_7 ;
    wire \transmit_module.X_DELTA_PATTERN_6 ;
    wire \line_buffer.n574 ;
    wire \line_buffer.n3785 ;
    wire \line_buffer.n566 ;
    wire \line_buffer.n577 ;
    wire \line_buffer.n513 ;
    wire \receive_module.rx_counter.Y_4 ;
    wire \receive_module.rx_counter.n4 ;
    wire \receive_module.rx_counter.Y_3 ;
    wire \receive_module.rx_counter.Y_1 ;
    wire \receive_module.rx_counter.n3657 ;
    wire \receive_module.rx_counter.n3619 ;
    wire \receive_module.rx_counter.n3648_cascade_ ;
    wire DEBUG_c_5_cascade_;
    wire \line_buffer.n641 ;
    wire \line_buffer.n609 ;
    wire bfn_13_10_0_;
    wire \receive_module.rx_counter.n3387 ;
    wire \receive_module.rx_counter.n3388 ;
    wire \receive_module.rx_counter.n3389 ;
    wire \receive_module.rx_counter.n3390 ;
    wire \receive_module.rx_counter.n3391 ;
    wire DEBUG_c_5;
    wire \transmit_module.video_signal_controller.VGA_X_4 ;
    wire \transmit_module.video_signal_controller.VGA_X_3 ;
    wire \transmit_module.video_signal_controller.VGA_X_5 ;
    wire \transmit_module.video_signal_controller.n21 ;
    wire \transmit_module.video_signal_controller.n3023_cascade_ ;
    wire \transmit_module.video_signal_controller.n3697_cascade_ ;
    wire \transmit_module.video_signal_controller.n8 ;
    wire \transmit_module.video_signal_controller.n3577 ;
    wire \transmit_module.video_signal_controller.n6_adj_568_cascade_ ;
    wire \transmit_module.video_signal_controller.n3603 ;
    wire \transmit_module.video_signal_controller.n6_cascade_ ;
    wire \transmit_module.video_signal_controller.n3575 ;
    wire \transmit_module.video_signal_controller.n2015 ;
    wire \transmit_module.video_signal_controller.n3857 ;
    wire \transmit_module.video_signal_controller.VGA_X_8 ;
    wire \transmit_module.video_signal_controller.n3856 ;
    wire \transmit_module.n220_cascade_ ;
    wire n28;
    wire \transmit_module.BRAM_ADDR_13_N_256_13 ;
    wire \transmit_module.n219_cascade_ ;
    wire n27;
    wire n1850;
    wire n1849;
    wire n1848;
    wire n1847;
    wire n1846;
    wire n1845;
    wire n1844;
    wire ADV_B_c;
    wire INVADV_R__i1C_net;
    wire n2404;
    wire \transmit_module.n220 ;
    wire \transmit_module.n218_cascade_ ;
    wire n26;
    wire \transmit_module.n187 ;
    wire \transmit_module.n219 ;
    wire \transmit_module.n187_cascade_ ;
    wire \transmit_module.n218 ;
    wire \transmit_module.n186 ;
    wire \transmit_module.n204 ;
    wire bfn_13_18_0_;
    wire \transmit_module.n203 ;
    wire \transmit_module.n3336 ;
    wire \transmit_module.n202 ;
    wire \transmit_module.n3337 ;
    wire \transmit_module.n3338 ;
    wire \transmit_module.n3339 ;
    wire \transmit_module.n199 ;
    wire \transmit_module.n3340 ;
    wire \transmit_module.n198 ;
    wire \transmit_module.n3341 ;
    wire \transmit_module.n3342 ;
    wire \transmit_module.n3343 ;
    wire \transmit_module.n196 ;
    wire bfn_13_19_0_;
    wire \transmit_module.n3344 ;
    wire \transmit_module.n3345 ;
    wire \transmit_module.n193 ;
    wire \transmit_module.n3346 ;
    wire \transmit_module.n192 ;
    wire \transmit_module.n3347 ;
    wire \transmit_module.n3348 ;
    wire \transmit_module.n191 ;
    wire \transmit_module.TX_ADDR_8 ;
    wire \transmit_module.ADDR_Y_COMPONENT_8 ;
    wire \transmit_module.X_DELTA_PATTERN_0 ;
    wire \transmit_module.X_DELTA_PATTERN_1 ;
    wire \transmit_module.X_DELTA_PATTERN_2 ;
    wire \transmit_module.X_DELTA_PATTERN_5 ;
    wire \transmit_module.X_DELTA_PATTERN_4 ;
    wire \transmit_module.X_DELTA_PATTERN_3 ;
    wire \transmit_module.n2099 ;
    wire \line_buffer.n3788 ;
    wire TX_DATA_6;
    wire \receive_module.rx_counter.FRAME_COUNTER_4 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_2 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_5 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_1 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_0 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_3 ;
    wire \receive_module.rx_counter.n3693_cascade_ ;
    wire \receive_module.rx_counter.n7 ;
    wire \receive_module.rx_counter.n11_cascade_ ;
    wire \receive_module.rx_counter.PULSE_1HZ_N_94 ;
    wire \receive_module.rx_counter.n2562 ;
    wire RX_ADDR_0;
    wire \receive_module.n136 ;
    wire bfn_14_11_0_;
    wire RX_ADDR_1;
    wire \receive_module.n135 ;
    wire \receive_module.n3323 ;
    wire RX_ADDR_2;
    wire \receive_module.n134 ;
    wire \receive_module.n3324 ;
    wire RX_ADDR_3;
    wire \receive_module.n133 ;
    wire \receive_module.n3325 ;
    wire RX_ADDR_4;
    wire \receive_module.n132 ;
    wire \receive_module.n3326 ;
    wire RX_ADDR_5;
    wire \receive_module.n131 ;
    wire \receive_module.n3327 ;
    wire RX_ADDR_6;
    wire \receive_module.n130 ;
    wire \receive_module.n3328 ;
    wire RX_ADDR_7;
    wire \receive_module.n129 ;
    wire \receive_module.n3329 ;
    wire \receive_module.n3330 ;
    wire RX_ADDR_8;
    wire \receive_module.n128 ;
    wire bfn_14_12_0_;
    wire RX_ADDR_9;
    wire \receive_module.n127 ;
    wire \receive_module.n3331 ;
    wire RX_ADDR_10;
    wire \receive_module.n126 ;
    wire \receive_module.n3332 ;
    wire RX_ADDR_11;
    wire \receive_module.n3333 ;
    wire RX_ADDR_12;
    wire \receive_module.n3334 ;
    wire \receive_module.n3854 ;
    wire DEBUG_c_3;
    wire \receive_module.n3335 ;
    wire \receive_module.n123 ;
    wire \transmit_module.video_signal_controller.VGA_Y_0 ;
    wire bfn_14_13_0_;
    wire \transmit_module.video_signal_controller.VGA_Y_1 ;
    wire \transmit_module.video_signal_controller.n3366 ;
    wire \transmit_module.video_signal_controller.VGA_Y_2 ;
    wire \transmit_module.video_signal_controller.n3367 ;
    wire \transmit_module.video_signal_controller.VGA_Y_3 ;
    wire \transmit_module.video_signal_controller.n3368 ;
    wire \transmit_module.video_signal_controller.VGA_Y_4 ;
    wire \transmit_module.video_signal_controller.n3369 ;
    wire \transmit_module.video_signal_controller.VGA_Y_5 ;
    wire \transmit_module.video_signal_controller.n3370 ;
    wire \transmit_module.video_signal_controller.VGA_Y_6 ;
    wire \transmit_module.video_signal_controller.n3371 ;
    wire \transmit_module.video_signal_controller.VGA_Y_7 ;
    wire \transmit_module.video_signal_controller.n3372 ;
    wire \transmit_module.video_signal_controller.n3373 ;
    wire \transmit_module.video_signal_controller.VGA_Y_8 ;
    wire bfn_14_14_0_;
    wire \transmit_module.video_signal_controller.VGA_Y_9 ;
    wire \transmit_module.video_signal_controller.n3374 ;
    wire \transmit_module.video_signal_controller.n3375 ;
    wire \transmit_module.video_signal_controller.n3376 ;
    wire \transmit_module.old_VGA_HS ;
    wire ADV_HSYNC_c;
    wire \transmit_module.n188 ;
    wire \transmit_module.n3859 ;
    wire \transmit_module.TX_ADDR_1 ;
    wire \transmit_module.ADDR_Y_COMPONENT_1 ;
    wire \transmit_module.ADDR_Y_COMPONENT_11 ;
    wire \transmit_module.ADDR_Y_COMPONENT_12 ;
    wire \transmit_module.ADDR_Y_COMPONENT_13 ;
    wire \transmit_module.TX_ADDR_0 ;
    wire \transmit_module.ADDR_Y_COMPONENT_0 ;
    wire \transmit_module.TX_ADDR_5 ;
    wire \transmit_module.ADDR_Y_COMPONENT_5 ;
    wire \transmit_module.TX_ADDR_6 ;
    wire \transmit_module.ADDR_Y_COMPONENT_6 ;
    wire \transmit_module.TX_ADDR_2 ;
    wire \transmit_module.ADDR_Y_COMPONENT_2 ;
    wire \transmit_module.ADDR_Y_COMPONENT_7 ;
    wire \transmit_module.ADDR_Y_COMPONENT_4 ;
    wire \transmit_module.n184_cascade_ ;
    wire \transmit_module.n200 ;
    wire \transmit_module.TX_ADDR_4 ;
    wire \transmit_module.n197 ;
    wire \transmit_module.n213_cascade_ ;
    wire \transmit_module.TX_ADDR_7 ;
    wire \transmit_module.n184 ;
    wire \transmit_module.n216 ;
    wire n24;
    wire \transmit_module.ADDR_Y_COMPONENT_9 ;
    wire \transmit_module.n181 ;
    wire \transmit_module.n213 ;
    wire n21;
    wire \line_buffer.n509 ;
    wire \line_buffer.n501 ;
    wire \line_buffer.n3770 ;
    wire \line_buffer.n571 ;
    wire \line_buffer.n563 ;
    wire \receive_module.rx_counter.n11 ;
    wire LED_c;
    wire \receive_module.rx_counter.n3862 ;
    wire TVP_VSYNC_c;
    wire \receive_module.BRAM_ADDR_13__N_31 ;
    wire \transmit_module.video_signal_controller.n2030 ;
    wire \transmit_module.video_signal_controller.n2551 ;
    wire DEBUG_c_6;
    wire \transmit_module.video_signal_controller.SYNC_BUFF1 ;
    wire \transmit_module.video_signal_controller.SYNC_BUFF2 ;
    wire n3852;
    wire \transmit_module.n2039 ;
    wire \line_buffer.n603 ;
    wire \line_buffer.n595 ;
    wire \line_buffer.n569 ;
    wire \line_buffer.n561 ;
    wire \line_buffer.n3830_cascade_ ;
    wire TX_DATA_1;
    wire \transmit_module.video_signal_controller.VGA_Y_11 ;
    wire \transmit_module.video_signal_controller.VGA_Y_10 ;
    wire \transmit_module.video_signal_controller.n3858 ;
    wire \transmit_module.Y_DELTA_PATTERN_38 ;
    wire \transmit_module.Y_DELTA_PATTERN_35 ;
    wire \transmit_module.Y_DELTA_PATTERN_37 ;
    wire \transmit_module.Y_DELTA_PATTERN_36 ;
    wire \transmit_module.Y_DELTA_PATTERN_40 ;
    wire \transmit_module.Y_DELTA_PATTERN_39 ;
    wire \transmit_module.Y_DELTA_PATTERN_34 ;
    wire \transmit_module.n3865 ;
    wire \line_buffer.n570 ;
    wire \line_buffer.n562 ;
    wire \line_buffer.n3705 ;
    wire \line_buffer.n3715 ;
    wire \line_buffer.n3773_cascade_ ;
    wire TX_DATA_3;
    wire \line_buffer.n594 ;
    wire \line_buffer.n602 ;
    wire \line_buffer.n497 ;
    wire \line_buffer.n3803_cascade_ ;
    wire \line_buffer.n505 ;
    wire \line_buffer.n3806_cascade_ ;
    wire \line_buffer.n3782 ;
    wire TX_DATA_2;
    wire \line_buffer.n635 ;
    wire \line_buffer.n627 ;
    wire \line_buffer.n3706 ;
    wire \line_buffer.n626 ;
    wire \line_buffer.n634 ;
    wire \line_buffer.n3779 ;
    wire \line_buffer.n3703 ;
    wire \line_buffer.n3791_cascade_ ;
    wire TX_DATA_7;
    wire \line_buffer.n575 ;
    wire \line_buffer.n567 ;
    wire \line_buffer.n3702 ;
    wire \transmit_module.ADDR_Y_COMPONENT_3 ;
    wire \transmit_module.n2321 ;
    wire \line_buffer.n625 ;
    wire \line_buffer.n633 ;
    wire \line_buffer.n3827 ;
    wire \line_buffer.n598 ;
    wire \line_buffer.n606 ;
    wire \line_buffer.n3767 ;
    wire \line_buffer.n506 ;
    wire \line_buffer.n498 ;
    wire \line_buffer.n3714 ;
    wire \line_buffer.n510 ;
    wire \line_buffer.n502 ;
    wire \line_buffer.n3717 ;
    wire \receive_module.rx_counter.n3547_cascade_ ;
    wire \receive_module.rx_counter.n3547 ;
    wire \receive_module.rx_counter.n3646_cascade_ ;
    wire \receive_module.rx_counter.n3613 ;
    wire \receive_module.rx_counter.n28 ;
    wire \line_buffer.n629 ;
    wire \line_buffer.n637 ;
    wire \line_buffer.n565 ;
    wire \line_buffer.n3761_cascade_ ;
    wire \line_buffer.n573 ;
    wire \line_buffer.n3764 ;
    wire TX_DATA_5;
    wire \transmit_module.Y_DELTA_PATTERN_33 ;
    wire \transmit_module.Y_DELTA_PATTERN_32 ;
    wire \transmit_module.n3864 ;
    wire \line_buffer.n607 ;
    wire \line_buffer.n599 ;
    wire \line_buffer.n3718 ;
    wire \transmit_module.n194 ;
    wire \transmit_module.n210_cascade_ ;
    wire \transmit_module.n201 ;
    wire \transmit_module.n217_cascade_ ;
    wire \transmit_module.TX_ADDR_3 ;
    wire \transmit_module.n3855 ;
    wire \transmit_module.n195 ;
    wire \transmit_module.TX_ADDR_9 ;
    wire \transmit_module.n3549 ;
    wire \transmit_module.n217 ;
    wire \transmit_module.n185 ;
    wire n25;
    wire \transmit_module.Y_DELTA_PATTERN_0 ;
    wire \transmit_module.ADDR_Y_COMPONENT_10 ;
    wire \transmit_module.TX_ADDR_10 ;
    wire \transmit_module.n178 ;
    wire \transmit_module.n210 ;
    wire \transmit_module.n178_cascade_ ;
    wire n18;
    wire GB_BUFFER_TVP_CLK_c_THRU_CO;
    wire TVP_HSYNC_c;
    wire \receive_module.rx_counter.n10 ;
    wire bfn_17_9_0_;
    wire \receive_module.rx_counter.n9 ;
    wire \receive_module.rx_counter.n3357 ;
    wire \receive_module.rx_counter.n8 ;
    wire \receive_module.rx_counter.n3358 ;
    wire \receive_module.rx_counter.X_3 ;
    wire \receive_module.rx_counter.n3359 ;
    wire \receive_module.rx_counter.X_4 ;
    wire \receive_module.rx_counter.n3360 ;
    wire \receive_module.rx_counter.X_5 ;
    wire \receive_module.rx_counter.n3361 ;
    wire \receive_module.rx_counter.X_6 ;
    wire \receive_module.rx_counter.n3362 ;
    wire \receive_module.rx_counter.X_7 ;
    wire \receive_module.rx_counter.n3363 ;
    wire \receive_module.rx_counter.n3364 ;
    wire \receive_module.rx_counter.X_8 ;
    wire bfn_17_10_0_;
    wire \receive_module.rx_counter.n3365 ;
    wire \receive_module.rx_counter.X_9 ;
    wire TVP_CLK_c;
    wire n3860;
    wire \line_buffer.n597 ;
    wire \line_buffer.n605 ;
    wire \line_buffer.n604 ;
    wire \line_buffer.n596 ;
    wire \line_buffer.n508 ;
    wire \line_buffer.n3833 ;
    wire \line_buffer.n500 ;
    wire \line_buffer.n3836 ;
    wire \line_buffer.n3721 ;
    wire TX_DATA_4;
    wire \transmit_module.n179 ;
    wire \transmit_module.n211 ;
    wire ADV_VSYNC_c;
    wire \transmit_module.n3853 ;
    wire n19;
    wire \line_buffer.n507 ;
    wire \line_buffer.n499 ;
    wire \line_buffer.n3720 ;
    wire \line_buffer.n592 ;
    wire \line_buffer.n600 ;
    wire \line_buffer.n572 ;
    wire \line_buffer.n564 ;
    wire \line_buffer.n503 ;
    wire \line_buffer.n3815 ;
    wire \line_buffer.n495 ;
    wire \line_buffer.n568 ;
    wire \line_buffer.n560 ;
    wire \line_buffer.n3824_cascade_ ;
    wire \line_buffer.n3818 ;
    wire TX_DATA_0;
    wire ADV_CLK_c;
    wire \line_buffer.n3699 ;
    wire DEBUG_c_2;
    wire \line_buffer.n3797 ;
    wire \line_buffer.n636 ;
    wire \line_buffer.n628 ;
    wire \line_buffer.n3700 ;
    wire \line_buffer.n624 ;
    wire \line_buffer.n632 ;
    wire \line_buffer.n3821 ;
    wire \line_buffer.n593 ;
    wire \line_buffer.n601 ;
    wire TX_ADDR_11;
    wire TX_ADDR_12;
    wire \line_buffer.n496 ;
    wire \line_buffer.n3809_cascade_ ;
    wire \line_buffer.n504 ;
    wire \line_buffer.n3812 ;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \tx_pll.TX_PLL_inst .TEST_MODE=1'b0;
    defparam \tx_pll.TX_PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \tx_pll.TX_PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \tx_pll.TX_PLL_inst .FILTER_RANGE=3'b010;
    defparam \tx_pll.TX_PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \tx_pll.TX_PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \tx_pll.TX_PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \tx_pll.TX_PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \tx_pll.TX_PLL_inst .DIVR=4'b0000;
    defparam \tx_pll.TX_PLL_inst .DIVQ=3'b100;
    defparam \tx_pll.TX_PLL_inst .DIVF=7'b0100110;
    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \tx_pll.TX_PLL_inst  (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(ADV_CLK_c),
            .REFERENCECLK(N__18875),
            .RESETB(N__22507),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .PLLOUTGLOBAL());
    defparam \line_buffer.mem2_physical .WRITE_MODE=3;
    defparam \line_buffer.mem2_physical .READ_MODE=3;
    defparam \line_buffer.mem2_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem2_physical  (
            .RDATA({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,\line_buffer.n510 ,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,\line_buffer.n509 ,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .RADDR({N__18946,N__19984,N__10507,N__16900,N__9670,N__10279,N__17137,N__19336,N__12127,N__11581,N__11806}),
            .WADDR({N__16030,N__13693,N__13948,N__14203,N__14437,N__14698,N__14926,N__15193,N__15454,N__13090,N__13324}),
            .MASK({dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37}),
            .WDATA({dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,N__8493,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,N__8636,dangling_wire_49,dangling_wire_50,dangling_wire_51}),
            .RCLKE(),
            .RCLK(N__21957),
            .RE(N__22516),
            .WCLKE(),
            .WCLK(N__21039),
            .WE(N__10778));
    defparam \line_buffer.mem14_physical .WRITE_MODE=3;
    defparam \line_buffer.mem14_physical .READ_MODE=3;
    defparam \line_buffer.mem14_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem14_physical  (
            .RDATA({dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,\line_buffer.n597 ,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,\line_buffer.n596 ,dangling_wire_63,dangling_wire_64,dangling_wire_65}),
            .RADDR({N__19018,N__20056,N__10579,N__16972,N__9742,N__10351,N__17209,N__19408,N__12199,N__11653,N__11878}),
            .WADDR({N__16102,N__13765,N__14020,N__14275,N__14509,N__14770,N__14998,N__15265,N__15526,N__13162,N__13396}),
            .MASK({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .WDATA({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,N__8421,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,N__8291,dangling_wire_93,dangling_wire_94,dangling_wire_95}),
            .RCLKE(),
            .RCLK(N__22053),
            .RE(N__22621),
            .WCLKE(),
            .WCLK(N__21024),
            .WE(N__10970));
    defparam \line_buffer.mem5_physical .WRITE_MODE=3;
    defparam \line_buffer.mem5_physical .READ_MODE=3;
    defparam \line_buffer.mem5_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem5_physical  (
            .RDATA({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,\line_buffer.n607 ,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\line_buffer.n606 ,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .RADDR({N__18949,N__19999,N__10510,N__16909,N__9679,N__10288,N__17146,N__19345,N__12130,N__11596,N__11827}),
            .WADDR({N__16045,N__13708,N__13969,N__14212,N__14452,N__14695,N__14953,N__15208,N__15463,N__13099,N__13357}),
            .MASK({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .WDATA({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,N__8520,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,N__8637,dangling_wire_137,dangling_wire_138,dangling_wire_139}),
            .RCLKE(),
            .RCLK(N__21490),
            .RE(N__22607),
            .WCLKE(),
            .WCLK(N__21035),
            .WE(N__9917));
    defparam \line_buffer.mem11_physical .WRITE_MODE=3;
    defparam \line_buffer.mem11_physical .READ_MODE=3;
    defparam \line_buffer.mem11_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem11_physical  (
            .RDATA({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,\line_buffer.n565 ,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,\line_buffer.n564 ,dangling_wire_151,dangling_wire_152,dangling_wire_153}),
            .RADDR({N__19054,N__20092,N__10615,N__17008,N__9778,N__10387,N__17245,N__19444,N__12235,N__11689,N__11914}),
            .WADDR({N__16138,N__13801,N__14056,N__14311,N__14545,N__14806,N__15034,N__15301,N__15562,N__13198,N__13432}),
            .MASK({dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169}),
            .WDATA({dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,N__8381,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,N__8270,dangling_wire_181,dangling_wire_182,dangling_wire_183}),
            .RCLKE(),
            .RCLK(N__22150),
            .RE(N__22667),
            .WCLKE(),
            .WCLK(N__21016),
            .WE(N__10831));
    defparam \line_buffer.mem21_physical .WRITE_MODE=3;
    defparam \line_buffer.mem21_physical .READ_MODE=3;
    defparam \line_buffer.mem21_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem21_physical  (
            .RDATA({dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,\line_buffer.n627 ,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,\line_buffer.n626 ,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .RADDR({N__18922,N__19960,N__10483,N__16876,N__9646,N__10255,N__17113,N__19312,N__12103,N__11557,N__11782}),
            .WADDR({N__16006,N__13669,N__13924,N__14179,N__14413,N__14674,N__14902,N__15169,N__15430,N__13066,N__13300}),
            .MASK({dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213}),
            .WDATA({dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,N__8210,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,N__8108,dangling_wire_225,dangling_wire_226,dangling_wire_227}),
            .RCLKE(),
            .RCLK(N__21808),
            .RE(N__22471),
            .WCLKE(),
            .WCLK(N__21043),
            .WE(N__11033));
    defparam \line_buffer.mem12_physical .WRITE_MODE=3;
    defparam \line_buffer.mem12_physical .READ_MODE=3;
    defparam \line_buffer.mem12_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem12_physical  (
            .RDATA({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,\line_buffer.n563 ,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,\line_buffer.n562 ,dangling_wire_239,dangling_wire_240,dangling_wire_241}),
            .RADDR({N__19042,N__20080,N__10603,N__16996,N__9766,N__10375,N__17233,N__19432,N__12223,N__11677,N__11902}),
            .WADDR({N__16126,N__13789,N__14044,N__14299,N__14533,N__14794,N__15022,N__15289,N__15550,N__13186,N__13420}),
            .MASK({dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .WDATA({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,N__8167,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,N__8100,dangling_wire_269,dangling_wire_270,dangling_wire_271}),
            .RCLKE(),
            .RCLK(N__22124),
            .RE(N__22508),
            .WCLKE(),
            .WCLK(N__21020),
            .WE(N__10814));
    defparam \line_buffer.mem18_physical .WRITE_MODE=3;
    defparam \line_buffer.mem18_physical .READ_MODE=3;
    defparam \line_buffer.mem18_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem18_physical  (
            .RDATA({dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,\line_buffer.n506 ,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,\line_buffer.n505 ,dangling_wire_283,dangling_wire_284,dangling_wire_285}),
            .RADDR({N__18970,N__20008,N__10531,N__16924,N__9694,N__10303,N__17161,N__19360,N__12151,N__11605,N__11830}),
            .WADDR({N__16054,N__13717,N__13972,N__14227,N__14461,N__14722,N__14950,N__15217,N__15478,N__13114,N__13348}),
            .MASK({dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301}),
            .WDATA({dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,N__8199,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,N__8101,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .RCLKE(),
            .RCLK(N__21765),
            .RE(N__22557),
            .WCLKE(),
            .WCLK(N__21032),
            .WE(N__10774));
    defparam \line_buffer.mem24_physical .WRITE_MODE=3;
    defparam \line_buffer.mem24_physical .READ_MODE=3;
    defparam \line_buffer.mem24_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem24_physical  (
            .RDATA({dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,\line_buffer.n571 ,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,\line_buffer.n570 ,dangling_wire_327,dangling_wire_328,dangling_wire_329}),
            .RADDR({N__19069,N__20119,N__10630,N__17029,N__9799,N__10408,N__17266,N__19465,N__12250,N__11716,N__11947}),
            .WADDR({N__16165,N__13828,N__14089,N__14332,N__14572,N__14815,N__15071,N__15328,N__15583,N__13219,N__13472}),
            .MASK({dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345}),
            .WDATA({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,N__8136,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,N__8025,dangling_wire_357,dangling_wire_358,dangling_wire_359}),
            .RCLKE(),
            .RCLK(N__21682),
            .RE(N__22693),
            .WCLKE(),
            .WCLK(N__21007),
            .WE(N__9468));
    defparam \line_buffer.mem1_physical .WRITE_MODE=3;
    defparam \line_buffer.mem1_physical .READ_MODE=3;
    defparam \line_buffer.mem1_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem1_physical  (
            .RDATA({dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,\line_buffer.n599 ,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,\line_buffer.n598 ,dangling_wire_371,dangling_wire_372,dangling_wire_373}),
            .RADDR({N__19078,N__20116,N__10639,N__17032,N__9802,N__10411,N__17269,N__19468,N__12259,N__11713,N__11938}),
            .WADDR({N__16162,N__13825,N__14080,N__14335,N__14569,N__14828,N__15058,N__15325,N__15586,N__13222,N__13456}),
            .MASK({dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389}),
            .WDATA({dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,N__8474,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,N__8600,dangling_wire_401,dangling_wire_402,dangling_wire_403}),
            .RCLKE(),
            .RCLK(N__22159),
            .RE(N__22684),
            .WCLKE(),
            .WCLK(N__21004),
            .WE(N__10977));
    defparam \line_buffer.mem15_physical .WRITE_MODE=3;
    defparam \line_buffer.mem15_physical .READ_MODE=3;
    defparam \line_buffer.mem15_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem15_physical  (
            .RDATA({dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,\line_buffer.n595 ,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,\line_buffer.n594 ,dangling_wire_415,dangling_wire_416,dangling_wire_417}),
            .RADDR({N__19006,N__20044,N__10567,N__16960,N__9730,N__10339,N__17197,N__19396,N__12187,N__11641,N__11866}),
            .WADDR({N__16090,N__13753,N__14008,N__14263,N__14497,N__14758,N__14986,N__15253,N__15514,N__13150,N__13384}),
            .MASK({dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .WDATA({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,N__8180,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,N__8092,dangling_wire_445,dangling_wire_446,dangling_wire_447}),
            .RCLKE(),
            .RCLK(N__22052),
            .RE(N__22620),
            .WCLKE(),
            .WCLK(N__21026),
            .WE(N__10978));
    defparam \line_buffer.mem27_physical .WRITE_MODE=3;
    defparam \line_buffer.mem27_physical .READ_MODE=3;
    defparam \line_buffer.mem27_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem27_physical  (
            .RDATA({dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,\line_buffer.n603 ,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,\line_buffer.n602 ,dangling_wire_459,dangling_wire_460,dangling_wire_461}),
            .RADDR({N__19033,N__20083,N__10594,N__16993,N__9763,N__10372,N__17230,N__19429,N__12214,N__11680,N__11911}),
            .WADDR({N__16129,N__13792,N__14053,N__14296,N__14536,N__14779,N__15037,N__15292,N__15547,N__13183,N__13441}),
            .MASK({dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477}),
            .WDATA({dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,N__8161,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,N__8056,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .RCLKE(),
            .RCLK(N__21959),
            .RE(N__22672),
            .WCLKE(),
            .WCLK(N__21021),
            .WE(N__9896));
    defparam \line_buffer.mem4_physical .WRITE_MODE=3;
    defparam \line_buffer.mem4_physical .READ_MODE=3;
    defparam \line_buffer.mem4_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem4_physical  (
            .RDATA({dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,\line_buffer.n575 ,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,\line_buffer.n574 ,dangling_wire_503,dangling_wire_504,dangling_wire_505}),
            .RADDR({N__18961,N__20011,N__10522,N__16921,N__9691,N__10300,N__17158,N__19357,N__12142,N__11608,N__11839}),
            .WADDR({N__16057,N__13720,N__13981,N__14224,N__14464,N__14707,N__14965,N__15220,N__15475,N__13111,N__13369}),
            .MASK({dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521}),
            .WDATA({dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,N__8499,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,N__8626,dangling_wire_533,dangling_wire_534,dangling_wire_535}),
            .RCLKE(),
            .RCLK(N__21723),
            .RE(N__22608),
            .WCLKE(),
            .WCLK(N__21033),
            .WE(N__9476));
    defparam \line_buffer.mem16_physical .WRITE_MODE=3;
    defparam \line_buffer.mem16_physical .READ_MODE=3;
    defparam \line_buffer.mem16_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem16_physical  (
            .RDATA({dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,\line_buffer.n593 ,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,\line_buffer.n592 ,dangling_wire_547,dangling_wire_548,dangling_wire_549}),
            .RADDR({N__18994,N__20032,N__10555,N__16948,N__9718,N__10327,N__17185,N__19384,N__12175,N__11629,N__11854}),
            .WADDR({N__16078,N__13741,N__13996,N__14251,N__14485,N__14746,N__14974,N__15241,N__15502,N__13138,N__13372}),
            .MASK({dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565}),
            .WDATA({dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,N__7962,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,N__8758,dangling_wire_577,dangling_wire_578,dangling_wire_579}),
            .RCLKE(),
            .RCLK(N__21926),
            .RE(N__22592),
            .WCLKE(),
            .WCLK(N__21028),
            .WE(N__10979));
    defparam \line_buffer.mem30_physical .WRITE_MODE=3;
    defparam \line_buffer.mem30_physical .READ_MODE=3;
    defparam \line_buffer.mem30_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem30_physical  (
            .RDATA({dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,\line_buffer.n635 ,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,\line_buffer.n634 ,dangling_wire_591,dangling_wire_592,dangling_wire_593}),
            .RADDR({N__18985,N__20035,N__10546,N__16945,N__9715,N__10324,N__17182,N__19381,N__12166,N__11632,N__11863}),
            .WADDR({N__16081,N__13744,N__14005,N__14248,N__14488,N__14731,N__14989,N__15244,N__15499,N__13135,N__13393}),
            .MASK({dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609}),
            .WDATA({dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,N__8186,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,N__8088,dangling_wire_621,dangling_wire_622,dangling_wire_623}),
            .RCLKE(),
            .RCLK(N__22089),
            .RE(N__22590),
            .WCLKE(),
            .WCLK(N__21029),
            .WE(N__9507));
    defparam \line_buffer.mem7_physical .WRITE_MODE=3;
    defparam \line_buffer.mem7_physical .READ_MODE=3;
    defparam \line_buffer.mem7_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem7_physical  (
            .RDATA({dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,\line_buffer.n502 ,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,\line_buffer.n501 ,dangling_wire_635,dangling_wire_636,dangling_wire_637}),
            .RADDR({N__18925,N__19975,N__10486,N__16885,N__9655,N__10264,N__17122,N__19321,N__12106,N__11572,N__11803}),
            .WADDR({N__16021,N__13684,N__13945,N__14188,N__14428,N__14671,N__14929,N__15184,N__15439,N__13075,N__13333}),
            .MASK({dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653}),
            .WDATA({dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,N__8528,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,N__8642,dangling_wire_665,dangling_wire_666,dangling_wire_667}),
            .RCLKE(),
            .RCLK(N__21446),
            .RE(N__22574),
            .WCLKE(),
            .WCLK(N__21042),
            .WE(N__9861));
    defparam \line_buffer.mem20_physical .WRITE_MODE=3;
    defparam \line_buffer.mem20_physical .READ_MODE=3;
    defparam \line_buffer.mem20_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem20_physical  (
            .RDATA({dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,\line_buffer.n629 ,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,\line_buffer.n628 ,dangling_wire_679,dangling_wire_680,dangling_wire_681}),
            .RADDR({N__18934,N__19972,N__10495,N__16888,N__9658,N__10267,N__17125,N__19324,N__12115,N__11569,N__11794}),
            .WADDR({N__16018,N__13681,N__13936,N__14191,N__14425,N__14686,N__14914,N__15181,N__15442,N__13078,N__13312}),
            .MASK({dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697}),
            .WDATA({dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,N__8420,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,N__8312,dangling_wire_709,dangling_wire_710,dangling_wire_711}),
            .RCLKE(),
            .RCLK(N__21809),
            .RE(N__22515),
            .WCLKE(),
            .WCLK(N__21041),
            .WE(N__11028));
    defparam \line_buffer.mem13_physical .WRITE_MODE=3;
    defparam \line_buffer.mem13_physical .READ_MODE=3;
    defparam \line_buffer.mem13_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem13_physical  (
            .RDATA({dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,\line_buffer.n561 ,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,\line_buffer.n560 ,dangling_wire_723,dangling_wire_724,dangling_wire_725}),
            .RADDR({N__19030,N__20068,N__10591,N__16984,N__9754,N__10363,N__17221,N__19420,N__12211,N__11665,N__11890}),
            .WADDR({N__16114,N__13777,N__14032,N__14287,N__14521,N__14782,N__15010,N__15277,N__15538,N__13174,N__13408}),
            .MASK({dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741}),
            .WDATA({dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,N__7947,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,N__8751,dangling_wire_753,dangling_wire_754,dangling_wire_755}),
            .RCLKE(),
            .RCLK(N__22123),
            .RE(N__22645),
            .WCLKE(),
            .WCLK(N__21022),
            .WE(N__10824));
    defparam \line_buffer.mem19_physical .WRITE_MODE=3;
    defparam \line_buffer.mem19_physical .READ_MODE=3;
    defparam \line_buffer.mem19_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem19_physical  (
            .RDATA({dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,\line_buffer.n504 ,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,\line_buffer.n503 ,dangling_wire_767,dangling_wire_768,dangling_wire_769}),
            .RADDR({N__18958,N__19996,N__10519,N__16912,N__9682,N__10291,N__17149,N__19348,N__12139,N__11593,N__11818}),
            .WADDR({N__16042,N__13705,N__13960,N__14215,N__14449,N__14710,N__14938,N__15205,N__15466,N__13102,N__13336}),
            .MASK({dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785}),
            .WDATA({dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,N__7969,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,N__8770,dangling_wire_797,dangling_wire_798,dangling_wire_799}),
            .RCLKE(),
            .RCLK(N__21958),
            .RE(N__22556),
            .WCLKE(),
            .WCLK(N__21034),
            .WE(N__10773));
    defparam \line_buffer.mem23_physical .WRITE_MODE=3;
    defparam \line_buffer.mem23_physical .READ_MODE=3;
    defparam \line_buffer.mem23_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem23_physical  (
            .RDATA({dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,\line_buffer.n573 ,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,\line_buffer.n572 ,dangling_wire_811,dangling_wire_812,dangling_wire_813}),
            .RADDR({N__19081,N__20129,N__10642,N__17041,N__9811,N__10420,N__17278,N__19477,N__12262,N__11726,N__11954}),
            .WADDR({N__16175,N__13838,N__14096,N__14344,N__14582,N__14827,N__15077,N__15338,N__15595,N__13231,N__13478}),
            .MASK({dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829}),
            .WDATA({dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,N__8397,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,N__8238,dangling_wire_841,dangling_wire_842,dangling_wire_843}),
            .RCLKE(),
            .RCLK(N__22137),
            .RE(N__22694),
            .WCLKE(),
            .WCLK(N__21003),
            .WE(N__9475));
    defparam \line_buffer.mem0_physical .WRITE_MODE=3;
    defparam \line_buffer.mem0_physical .READ_MODE=3;
    defparam \line_buffer.mem0_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem0_physical  (
            .RDATA({dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,\line_buffer.n567 ,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,\line_buffer.n566 ,dangling_wire_855,dangling_wire_856,dangling_wire_857}),
            .RADDR({N__19085,N__20128,N__10646,N__17042,N__9812,N__10421,N__17279,N__19478,N__12266,N__11725,N__11950}),
            .WADDR({N__16174,N__13837,N__14092,N__14345,N__14581,N__14834,N__15070,N__15337,N__15596,N__13232,N__13468}),
            .MASK({dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873}),
            .WDATA({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,N__8449,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,N__8599,dangling_wire_885,dangling_wire_886,dangling_wire_887}),
            .RCLKE(),
            .RCLK(N__22160),
            .RE(N__22555),
            .WCLKE(),
            .WCLK(N__21001),
            .WE(N__10832));
    defparam \line_buffer.mem26_physical .WRITE_MODE=3;
    defparam \line_buffer.mem26_physical .READ_MODE=3;
    defparam \line_buffer.mem26_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem26_physical  (
            .RDATA({dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,\line_buffer.n605 ,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,\line_buffer.n604 ,dangling_wire_899,dangling_wire_900,dangling_wire_901}),
            .RADDR({N__19045,N__20095,N__10606,N__17005,N__9775,N__10384,N__17242,N__19441,N__12226,N__11692,N__11923}),
            .WADDR({N__16141,N__13804,N__14065,N__14308,N__14548,N__14791,N__15049,N__15304,N__15559,N__13195,N__13453}),
            .MASK({dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917}),
            .WDATA({dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,N__8380,dangling_wire_922,dangling_wire_923,dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,dangling_wire_928,N__8263,dangling_wire_929,dangling_wire_930,dangling_wire_931}),
            .RCLKE(),
            .RCLK(N__22158),
            .RE(N__22685),
            .WCLKE(),
            .WCLK(N__21019),
            .WE(N__9907));
    defparam \line_buffer.mem3_physical .WRITE_MODE=3;
    defparam \line_buffer.mem3_physical .READ_MODE=3;
    defparam \line_buffer.mem3_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem3_physical  (
            .RDATA({dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,\line_buffer.n631 ,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,\line_buffer.n630 ,dangling_wire_943,dangling_wire_944,dangling_wire_945}),
            .RADDR({N__18997,N__20047,N__10558,N__16957,N__9727,N__10336,N__17194,N__19393,N__12178,N__11644,N__11875}),
            .WADDR({N__16093,N__13756,N__14017,N__14260,N__14500,N__14743,N__15001,N__15256,N__15511,N__13147,N__13405}),
            .MASK({dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961}),
            .WDATA({dangling_wire_962,dangling_wire_963,dangling_wire_964,dangling_wire_965,N__8506,dangling_wire_966,dangling_wire_967,dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,dangling_wire_972,N__8612,dangling_wire_973,dangling_wire_974,dangling_wire_975}),
            .RCLKE(),
            .RCLK(N__21553),
            .RE(N__22652),
            .WCLKE(),
            .WCLK(N__21027),
            .WE(N__11027));
    defparam \line_buffer.mem17_physical .WRITE_MODE=3;
    defparam \line_buffer.mem17_physical .READ_MODE=3;
    defparam \line_buffer.mem17_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem17_physical  (
            .RDATA({dangling_wire_976,dangling_wire_977,dangling_wire_978,dangling_wire_979,\line_buffer.n508 ,dangling_wire_980,dangling_wire_981,dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,\line_buffer.n507 ,dangling_wire_987,dangling_wire_988,dangling_wire_989}),
            .RADDR({N__18982,N__20020,N__10543,N__16936,N__9706,N__10315,N__17173,N__19372,N__12163,N__11617,N__11842}),
            .WADDR({N__16066,N__13729,N__13984,N__14239,N__14473,N__14734,N__14962,N__15229,N__15490,N__13126,N__13360}),
            .MASK({dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997,dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005}),
            .WDATA({dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,dangling_wire_1009,N__8404,dangling_wire_1010,dangling_wire_1011,dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,dangling_wire_1016,N__8301,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019}),
            .RCLKE(),
            .RCLK(N__21925),
            .RE(N__22591),
            .WCLKE(),
            .WCLK(N__21030),
            .WE(N__10766));
    defparam \line_buffer.mem31_physical .WRITE_MODE=3;
    defparam \line_buffer.mem31_physical .READ_MODE=3;
    defparam \line_buffer.mem31_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem31_physical  (
            .RDATA({dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,dangling_wire_1023,\line_buffer.n633 ,dangling_wire_1024,dangling_wire_1025,dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,\line_buffer.n632 ,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033}),
            .RADDR({N__18973,N__20023,N__10534,N__16933,N__9703,N__10312,N__17170,N__19369,N__12154,N__11620,N__11851}),
            .WADDR({N__16069,N__13732,N__13993,N__14236,N__14476,N__14719,N__14977,N__15232,N__15487,N__13123,N__13381}),
            .MASK({dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041,dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049}),
            .WDATA({dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,dangling_wire_1053,N__7929,dangling_wire_1054,dangling_wire_1055,dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,dangling_wire_1060,N__8736,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063}),
            .RCLKE(),
            .RCLK(N__22119),
            .RE(N__22631),
            .WCLKE(),
            .WCLK(N__21031),
            .WE(N__9514));
    defparam \line_buffer.mem9_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .WRITE_MODE=3;
    defparam \line_buffer.mem9_physical .READ_MODE=3;
    defparam \line_buffer.mem9_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem9_physical  (
            .RDATA({dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,dangling_wire_1067,\line_buffer.n498 ,dangling_wire_1068,dangling_wire_1069,dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,\line_buffer.n497 ,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077}),
            .RADDR({N__18901,N__19951,N__10462,N__16861,N__9631,N__10240,N__17098,N__19297,N__12082,N__11548,N__11779}),
            .WADDR({N__15997,N__13660,N__13921,N__14164,N__14404,N__14647,N__14905,N__15160,N__15415,N__13051,N__13309}),
            .MASK({dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085,dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093}),
            .WDATA({dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,dangling_wire_1097,N__8209,dangling_wire_1098,dangling_wire_1099,dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,dangling_wire_1104,N__8099,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107}),
            .RCLKE(),
            .RCLK(N__21509),
            .RE(N__22533),
            .WCLKE(),
            .WCLK(N__21046),
            .WE(N__9869));
    defparam \line_buffer.mem29_physical .WRITE_MODE=3;
    defparam \line_buffer.mem29_physical .READ_MODE=3;
    defparam \line_buffer.mem29_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem29_physical  (
            .RDATA({dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,dangling_wire_1111,\line_buffer.n637 ,dangling_wire_1112,dangling_wire_1113,dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,\line_buffer.n636 ,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121}),
            .RADDR({N__19009,N__20059,N__10570,N__16969,N__9739,N__10348,N__17206,N__19405,N__12190,N__11656,N__11887}),
            .WADDR({N__16105,N__13768,N__14029,N__14272,N__14512,N__14755,N__15013,N__15268,N__15523,N__13159,N__13417}),
            .MASK({dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129,dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137}),
            .WDATA({dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,dangling_wire_1141,N__8422,dangling_wire_1142,dangling_wire_1143,dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,dangling_wire_1148,N__8276,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151}),
            .RCLKE(),
            .RCLK(N__21817),
            .RE(N__22653),
            .WCLKE(),
            .WCLK(N__21025),
            .WE(N__9498));
    defparam \line_buffer.mem6_physical .WRITE_MODE=3;
    defparam \line_buffer.mem6_physical .READ_MODE=3;
    defparam \line_buffer.mem6_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem6_physical  (
            .RDATA({dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,dangling_wire_1155,\line_buffer.n639 ,dangling_wire_1156,dangling_wire_1157,dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,\line_buffer.n638 ,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165}),
            .RADDR({N__18937,N__19987,N__10498,N__16897,N__9667,N__10276,N__17134,N__19333,N__12118,N__11584,N__11815}),
            .WADDR({N__16033,N__13696,N__13957,N__14200,N__14440,N__14683,N__14941,N__15196,N__15451,N__13087,N__13345}),
            .MASK({dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173,dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181}),
            .WDATA({dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,dangling_wire_1185,N__8527,dangling_wire_1186,dangling_wire_1187,dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,dangling_wire_1192,N__8638,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195}),
            .RCLKE(),
            .RCLK(N__21782),
            .RE(N__22575),
            .WCLKE(),
            .WCLK(N__21040),
            .WE(N__9518));
    defparam \line_buffer.mem10_physical .WRITE_MODE=3;
    defparam \line_buffer.mem10_physical .READ_MODE=3;
    defparam \line_buffer.mem10_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem10_physical  (
            .RDATA({dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,dangling_wire_1199,\line_buffer.n496 ,dangling_wire_1200,dangling_wire_1201,dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,\line_buffer.n495 ,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209}),
            .RADDR({N__19066,N__20104,N__10627,N__17020,N__9790,N__10399,N__17257,N__19456,N__12247,N__11701,N__11926}),
            .WADDR({N__16150,N__13813,N__14068,N__14323,N__14557,N__14818,N__15046,N__15313,N__15574,N__13210,N__13444}),
            .MASK({dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217,dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225}),
            .WDATA({dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,dangling_wire_1229,N__7938,dangling_wire_1230,dangling_wire_1231,dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,dangling_wire_1236,N__8737,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239}),
            .RCLKE(),
            .RCLK(N__22151),
            .RE(N__22554),
            .WCLKE(),
            .WCLK(N__21008),
            .WE(N__9852));
    defparam \line_buffer.mem22_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .WRITE_MODE=3;
    defparam \line_buffer.mem22_physical .READ_MODE=3;
    defparam \line_buffer.mem22_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem22_physical  (
            .RDATA({dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,dangling_wire_1243,\line_buffer.n625 ,dangling_wire_1244,dangling_wire_1245,dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,\line_buffer.n624 ,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253}),
            .RADDR({N__18910,N__19948,N__10471,N__16864,N__9634,N__10243,N__17101,N__19300,N__12091,N__11545,N__11770}),
            .WADDR({N__15994,N__13657,N__13912,N__14167,N__14401,N__14662,N__14890,N__15157,N__15418,N__13054,N__13288}),
            .MASK({dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261,dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269}),
            .WDATA({dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,dangling_wire_1273,N__7976,dangling_wire_1274,dangling_wire_1275,dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,dangling_wire_1280,N__8777,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283}),
            .RCLKE(),
            .RCLK(N__21804),
            .RE(N__22432),
            .WCLKE(),
            .WCLK(N__21045),
            .WE(N__11029));
    defparam \line_buffer.mem25_physical .WRITE_MODE=3;
    defparam \line_buffer.mem25_physical .READ_MODE=3;
    defparam \line_buffer.mem25_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem25_physical  (
            .RDATA({dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,dangling_wire_1287,\line_buffer.n569 ,dangling_wire_1288,dangling_wire_1289,dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,\line_buffer.n568 ,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297}),
            .RADDR({N__19057,N__20107,N__10618,N__17017,N__9787,N__10396,N__17254,N__19453,N__12238,N__11704,N__11935}),
            .WADDR({N__16153,N__13816,N__14077,N__14320,N__14560,N__14803,N__15061,N__15316,N__15571,N__13207,N__13465}),
            .MASK({dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305,dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313}),
            .WDATA({dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,dangling_wire_1317,N__7920,dangling_wire_1318,dangling_wire_1319,dangling_wire_1320,dangling_wire_1321,dangling_wire_1322,dangling_wire_1323,dangling_wire_1324,N__8705,dangling_wire_1325,dangling_wire_1326,dangling_wire_1327}),
            .RCLKE(),
            .RCLK(N__22073),
            .RE(N__22686),
            .WCLKE(),
            .WCLK(N__21011),
            .WE(N__9458));
    defparam \line_buffer.mem8_physical .WRITE_MODE=3;
    defparam \line_buffer.mem8_physical .READ_MODE=3;
    defparam \line_buffer.mem8_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem8_physical  (
            .RDATA({dangling_wire_1328,dangling_wire_1329,dangling_wire_1330,dangling_wire_1331,\line_buffer.n500 ,dangling_wire_1332,dangling_wire_1333,dangling_wire_1334,dangling_wire_1335,dangling_wire_1336,dangling_wire_1337,dangling_wire_1338,\line_buffer.n499 ,dangling_wire_1339,dangling_wire_1340,dangling_wire_1341}),
            .RADDR({N__18913,N__19963,N__10474,N__16873,N__9643,N__10252,N__17110,N__19309,N__12094,N__11560,N__11791}),
            .WADDR({N__16009,N__13672,N__13933,N__14176,N__14416,N__14659,N__14917,N__15172,N__15427,N__13063,N__13321}),
            .MASK({dangling_wire_1342,dangling_wire_1343,dangling_wire_1344,dangling_wire_1345,dangling_wire_1346,dangling_wire_1347,dangling_wire_1348,dangling_wire_1349,dangling_wire_1350,dangling_wire_1351,dangling_wire_1352,dangling_wire_1353,dangling_wire_1354,dangling_wire_1355,dangling_wire_1356,dangling_wire_1357}),
            .WDATA({dangling_wire_1358,dangling_wire_1359,dangling_wire_1360,dangling_wire_1361,N__8426,dangling_wire_1362,dangling_wire_1363,dangling_wire_1364,dangling_wire_1365,dangling_wire_1366,dangling_wire_1367,dangling_wire_1368,N__8311,dangling_wire_1369,dangling_wire_1370,dangling_wire_1371}),
            .RCLKE(),
            .RCLK(N__21628),
            .RE(N__22534),
            .WCLKE(),
            .WCLK(N__21044),
            .WE(N__9868));
    defparam \line_buffer.mem28_physical .WRITE_MODE=3;
    defparam \line_buffer.mem28_physical .READ_MODE=3;
    defparam \line_buffer.mem28_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem28_physical  (
            .RDATA({dangling_wire_1372,dangling_wire_1373,dangling_wire_1374,dangling_wire_1375,\line_buffer.n601 ,dangling_wire_1376,dangling_wire_1377,dangling_wire_1378,dangling_wire_1379,dangling_wire_1380,dangling_wire_1381,dangling_wire_1382,\line_buffer.n600 ,dangling_wire_1383,dangling_wire_1384,dangling_wire_1385}),
            .RADDR({N__19021,N__20071,N__10582,N__16981,N__9751,N__10360,N__17218,N__19417,N__12202,N__11668,N__11899}),
            .WADDR({N__16117,N__13780,N__14041,N__14284,N__14524,N__14767,N__15025,N__15280,N__15535,N__13171,N__13429}),
            .MASK({dangling_wire_1386,dangling_wire_1387,dangling_wire_1388,dangling_wire_1389,dangling_wire_1390,dangling_wire_1391,dangling_wire_1392,dangling_wire_1393,dangling_wire_1394,dangling_wire_1395,dangling_wire_1396,dangling_wire_1397,dangling_wire_1398,dangling_wire_1399,dangling_wire_1400,dangling_wire_1401}),
            .WDATA({dangling_wire_1402,dangling_wire_1403,dangling_wire_1404,dangling_wire_1405,N__7919,dangling_wire_1406,dangling_wire_1407,dangling_wire_1408,dangling_wire_1409,dangling_wire_1410,dangling_wire_1411,dangling_wire_1412,N__8718,dangling_wire_1413,dangling_wire_1414,dangling_wire_1415}),
            .RCLKE(),
            .RCLK(N__22144),
            .RE(N__22671),
            .WCLKE(),
            .WCLK(N__21023),
            .WE(N__9906));
    PRE_IO_GBUF TVP_CLK_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__23673),
            .GLOBALBUFFEROUTPUT(TVP_CLK_c));
    defparam TVP_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_CLK_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_CLK_pad_iopad (
            .OE(N__23675),
            .DIN(N__23674),
            .DOUT(N__23673),
            .PACKAGEPIN(TVP_CLK));
    defparam TVP_CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_CLK_pad_preio (
            .PADOEN(N__23675),
            .PADOUT(N__23674),
            .PADIN(N__23673),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_CLK_pad_iopad (
            .OE(N__23664),
            .DIN(N__23663),
            .DOUT(N__23662),
            .PACKAGEPIN(ADV_CLK));
    defparam ADV_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_CLK_pad_preio (
            .PADOEN(N__23664),
            .PADOUT(N__23663),
            .PADIN(N__23662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21956),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_3_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_3_iopad (
            .OE(N__23655),
            .DIN(N__23654),
            .DOUT(N__23653),
            .PACKAGEPIN(DEBUG[3]));
    defparam DEBUG_pad_3_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_3_preio (
            .PADOEN(N__23655),
            .PADOUT(N__23654),
            .PADIN(N__23653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15773),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_2_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_2_iopad (
            .OE(N__23646),
            .DIN(N__23645),
            .DOUT(N__23644),
            .PACKAGEPIN(TVP_VIDEO[2]));
    defparam TVP_VIDEO_pad_2_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_2_preio (
            .PADOEN(N__23646),
            .PADOUT(N__23645),
            .PADIN(N__23644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_5_iopad (
            .OE(N__23637),
            .DIN(N__23636),
            .DOUT(N__23635),
            .PACKAGEPIN(ADV_G[5]));
    defparam ADV_G_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_5_preio (
            .PADOEN(N__23637),
            .PADOUT(N__23636),
            .PADIN(N__23635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12470),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_3_iopad (
            .OE(N__23628),
            .DIN(N__23627),
            .DOUT(N__23626),
            .PACKAGEPIN(ADV_R[3]));
    defparam ADV_R_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_3_preio (
            .PADOEN(N__23628),
            .PADOUT(N__23627),
            .PADIN(N__23626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12579),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_5_iopad (
            .OE(N__23619),
            .DIN(N__23618),
            .DOUT(N__23617),
            .PACKAGEPIN(ADV_B[5]));
    defparam ADV_B_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_5_preio (
            .PADOEN(N__23619),
            .PADOUT(N__23618),
            .PADIN(N__23617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12469),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_7_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_7_iopad (
            .OE(N__23610),
            .DIN(N__23609),
            .DOUT(N__23608),
            .PACKAGEPIN(DEBUG[7]));
    defparam DEBUG_pad_7_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_7_preio (
            .PADOEN(N__23610),
            .PADOUT(N__23609),
            .PADIN(N__23608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_6_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_6_iopad (
            .OE(N__23601),
            .DIN(N__23600),
            .DOUT(N__23599),
            .PACKAGEPIN(TVP_VIDEO[6]));
    defparam TVP_VIDEO_pad_6_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_6_preio (
            .PADOEN(N__23601),
            .PADOUT(N__23600),
            .PADIN(N__23599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_1_iopad (
            .OE(N__23592),
            .DIN(N__23591),
            .DOUT(N__23590),
            .PACKAGEPIN(ADV_G[1]));
    defparam ADV_G_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_1_preio (
            .PADOEN(N__23592),
            .PADOUT(N__23591),
            .PADIN(N__23590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11453),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_0_iopad (
            .OE(N__23583),
            .DIN(N__23582),
            .DOUT(N__23581),
            .PACKAGEPIN(ADV_R[0]));
    defparam ADV_R_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_0_preio (
            .PADOEN(N__23583),
            .PADOUT(N__23582),
            .PADIN(N__23581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11506),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_2_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_2_iopad (
            .OE(N__23574),
            .DIN(N__23573),
            .DOUT(N__23572),
            .PACKAGEPIN(DEBUG[2]));
    defparam DEBUG_pad_2_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_2_preio (
            .PADOEN(N__23574),
            .PADOUT(N__23573),
            .PADIN(N__23572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21296),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_3_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_3_iopad (
            .OE(N__23565),
            .DIN(N__23564),
            .DOUT(N__23563),
            .PACKAGEPIN(TVP_VIDEO[3]));
    defparam TVP_VIDEO_pad_3_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_3_preio (
            .PADOEN(N__23565),
            .PADOUT(N__23564),
            .PADIN(N__23563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_4_iopad (
            .OE(N__23556),
            .DIN(N__23555),
            .DOUT(N__23554),
            .PACKAGEPIN(ADV_G[4]));
    defparam ADV_G_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_4_preio (
            .PADOEN(N__23556),
            .PADOUT(N__23555),
            .PADIN(N__23554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12516),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_5_iopad (
            .OE(N__23547),
            .DIN(N__23546),
            .DOUT(N__23545),
            .PACKAGEPIN(ADV_R[5]));
    defparam ADV_R_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_5_preio (
            .PADOEN(N__23547),
            .PADOUT(N__23546),
            .PADIN(N__23545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12468),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_9_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_9_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_9_iopad (
            .OE(N__23538),
            .DIN(N__23537),
            .DOUT(N__23536),
            .PACKAGEPIN(TVP_VIDEO[9]));
    defparam TVP_VIDEO_pad_9_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_9_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_9_preio (
            .PADOEN(N__23538),
            .PADOUT(N__23537),
            .PADIN(N__23536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_1_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_1_iopad (
            .OE(N__23529),
            .DIN(N__23528),
            .DOUT(N__23527),
            .PACKAGEPIN(DEBUG[1]));
    defparam DEBUG_pad_1_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_1_preio (
            .PADOEN(N__23529),
            .PADOUT(N__23528),
            .PADIN(N__23527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_1_iopad (
            .OE(N__23520),
            .DIN(N__23519),
            .DOUT(N__23518),
            .PACKAGEPIN(ADV_B[1]));
    defparam ADV_B_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_1_preio (
            .PADOEN(N__23520),
            .PADOUT(N__23519),
            .PADIN(N__23518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11448),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_SYNC_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_SYNC_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_SYNC_N_pad_iopad (
            .OE(N__23511),
            .DIN(N__23510),
            .DOUT(N__23509),
            .PACKAGEPIN(ADV_SYNC_N));
    defparam ADV_SYNC_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_SYNC_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_SYNC_N_pad_preio (
            .PADOEN(N__23511),
            .PADOUT(N__23510),
            .PADIN(N__23509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_6_iopad (
            .OE(N__23502),
            .DIN(N__23501),
            .DOUT(N__23500),
            .PACKAGEPIN(ADV_B[6]));
    defparam ADV_B_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_6_preio (
            .PADOEN(N__23502),
            .PADOUT(N__23501),
            .PADIN(N__23500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12416),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_6_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_6_iopad (
            .OE(N__23493),
            .DIN(N__23492),
            .DOUT(N__23491),
            .PACKAGEPIN(DEBUG[6]));
    defparam DEBUG_pad_6_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_6_preio (
            .PADOEN(N__23493),
            .PADOUT(N__23492),
            .PADIN(N__23491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17573),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_7_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_7_iopad (
            .OE(N__23484),
            .DIN(N__23483),
            .DOUT(N__23482),
            .PACKAGEPIN(TVP_VIDEO[7]));
    defparam TVP_VIDEO_pad_7_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_7_preio (
            .PADOEN(N__23484),
            .PADOUT(N__23483),
            .PADIN(N__23482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_0_iopad (
            .OE(N__23475),
            .DIN(N__23474),
            .DOUT(N__23473),
            .PACKAGEPIN(ADV_G[0]));
    defparam ADV_G_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_0_preio (
            .PADOEN(N__23475),
            .PADOUT(N__23474),
            .PADIN(N__23473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11507),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_1_iopad (
            .OE(N__23466),
            .DIN(N__23465),
            .DOUT(N__23464),
            .PACKAGEPIN(ADV_R[1]));
    defparam ADV_R_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_1_preio (
            .PADOEN(N__23466),
            .PADOUT(N__23465),
            .PADIN(N__23464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11449),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_5_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_5_iopad (
            .OE(N__23457),
            .DIN(N__23456),
            .DOUT(N__23455),
            .PACKAGEPIN(DEBUG[5]));
    defparam DEBUG_pad_5_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_5_preio (
            .PADOEN(N__23457),
            .PADOUT(N__23456),
            .PADIN(N__23455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11333),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_HSYNC_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_HSYNC_pad_iopad (
            .OE(N__23448),
            .DIN(N__23447),
            .DOUT(N__23446),
            .PACKAGEPIN(TVP_HSYNC));
    defparam TVP_HSYNC_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_HSYNC_pad_preio (
            .PADOEN(N__23448),
            .PADOUT(N__23447),
            .PADIN(N__23446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_HSYNC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_7_iopad (
            .OE(N__23439),
            .DIN(N__23438),
            .DOUT(N__23437),
            .PACKAGEPIN(ADV_G[7]));
    defparam ADV_G_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_7_preio (
            .PADOEN(N__23439),
            .PADOUT(N__23438),
            .PADIN(N__23437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12345),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_6_iopad (
            .OE(N__23430),
            .DIN(N__23429),
            .DOUT(N__23428),
            .PACKAGEPIN(ADV_R[6]));
    defparam ADV_R_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_6_preio (
            .PADOEN(N__23430),
            .PADOUT(N__23429),
            .PADIN(N__23428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12412),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VSYNC_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_VSYNC_pad_iopad (
            .OE(N__23421),
            .DIN(N__23420),
            .DOUT(N__23419),
            .PACKAGEPIN(TVP_VSYNC));
    defparam TVP_VSYNC_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VSYNC_pad_preio (
            .PADOEN(N__23421),
            .PADOUT(N__23420),
            .PADIN(N__23419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VSYNC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_BLANK_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_BLANK_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_BLANK_N_pad_iopad (
            .OE(N__23412),
            .DIN(N__23411),
            .DOUT(N__23410),
            .PACKAGEPIN(ADV_BLANK_N));
    defparam ADV_BLANK_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_BLANK_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_BLANK_N_pad_preio (
            .PADOEN(N__23412),
            .PADOUT(N__23411),
            .PADIN(N__23410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22506),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_0_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_0_iopad (
            .OE(N__23403),
            .DIN(N__23402),
            .DOUT(N__23401),
            .PACKAGEPIN(DEBUG[0]));
    defparam DEBUG_pad_0_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_0_preio (
            .PADOEN(N__23403),
            .PADOUT(N__23402),
            .PADIN(N__23401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_2_iopad (
            .OE(N__23394),
            .DIN(N__23393),
            .DOUT(N__23392),
            .PACKAGEPIN(ADV_B[2]));
    defparam ADV_B_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_2_preio (
            .PADOEN(N__23394),
            .PADOUT(N__23393),
            .PADIN(N__23392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12637),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_7_iopad (
            .OE(N__23385),
            .DIN(N__23384),
            .DOUT(N__23383),
            .PACKAGEPIN(ADV_B[7]));
    defparam ADV_B_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_7_preio (
            .PADOEN(N__23385),
            .PADOUT(N__23384),
            .PADIN(N__23383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12353),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__23376),
            .DIN(N__23375),
            .DOUT(N__23374),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__23376),
            .PADOUT(N__23375),
            .PADIN(N__23374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16748),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_4_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_4_iopad (
            .OE(N__23367),
            .DIN(N__23366),
            .DOUT(N__23365),
            .PACKAGEPIN(TVP_VIDEO[4]));
    defparam TVP_VIDEO_pad_4_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_4_preio (
            .PADOEN(N__23367),
            .PADOUT(N__23366),
            .PADIN(N__23365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_3_iopad (
            .OE(N__23358),
            .DIN(N__23357),
            .DOUT(N__23356),
            .PACKAGEPIN(ADV_G[3]));
    defparam ADV_G_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_3_preio (
            .PADOEN(N__23358),
            .PADOUT(N__23357),
            .PADIN(N__23356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12580),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_HSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_HSYNC_pad_iopad (
            .OE(N__23349),
            .DIN(N__23348),
            .DOUT(N__23347),
            .PACKAGEPIN(ADV_HSYNC));
    defparam ADV_HSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_HSYNC_pad_preio (
            .PADOEN(N__23349),
            .PADOUT(N__23348),
            .PADIN(N__23347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16235),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_2_iopad (
            .OE(N__23340),
            .DIN(N__23339),
            .DOUT(N__23338),
            .PACKAGEPIN(ADV_R[2]));
    defparam ADV_R_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_2_preio (
            .PADOEN(N__23340),
            .PADOUT(N__23339),
            .PADIN(N__23338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12636),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_4_iopad (
            .OE(N__23331),
            .DIN(N__23330),
            .DOUT(N__23329),
            .PACKAGEPIN(ADV_B[4]));
    defparam ADV_B_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_4_preio (
            .PADOEN(N__23331),
            .PADOUT(N__23330),
            .PADIN(N__23329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12524),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_4_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_4_iopad (
            .OE(N__23322),
            .DIN(N__23321),
            .DOUT(N__23320),
            .PACKAGEPIN(DEBUG[4]));
    defparam DEBUG_pad_4_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_4_preio (
            .PADOEN(N__23322),
            .PADOUT(N__23321),
            .PADIN(N__23320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17528),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_6_iopad (
            .OE(N__23313),
            .DIN(N__23312),
            .DOUT(N__23311),
            .PACKAGEPIN(ADV_G[6]));
    defparam ADV_G_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_6_preio (
            .PADOEN(N__23313),
            .PADOUT(N__23312),
            .PADIN(N__23311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12411),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_7_iopad (
            .OE(N__23304),
            .DIN(N__23303),
            .DOUT(N__23302),
            .PACKAGEPIN(ADV_R[7]));
    defparam ADV_R_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_7_preio (
            .PADOEN(N__23304),
            .PADOUT(N__23303),
            .PADIN(N__23302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12349),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_3_iopad (
            .OE(N__23295),
            .DIN(N__23294),
            .DOUT(N__23293),
            .PACKAGEPIN(ADV_B[3]));
    defparam ADV_B_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_3_preio (
            .PADOEN(N__23295),
            .PADOUT(N__23294),
            .PADIN(N__23293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12581),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_4_iopad (
            .OE(N__23286),
            .DIN(N__23285),
            .DOUT(N__23284),
            .PACKAGEPIN(ADV_R[4]));
    defparam ADV_R_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_4_preio (
            .PADOEN(N__23286),
            .PADOUT(N__23285),
            .PADIN(N__23284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12523),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_8_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_8_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_8_iopad (
            .OE(N__23277),
            .DIN(N__23276),
            .DOUT(N__23275),
            .PACKAGEPIN(TVP_VIDEO[8]));
    defparam TVP_VIDEO_pad_8_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_8_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_8_preio (
            .PADOEN(N__23277),
            .PADOUT(N__23276),
            .PADIN(N__23275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_0_iopad (
            .OE(N__23268),
            .DIN(N__23267),
            .DOUT(N__23266),
            .PACKAGEPIN(ADV_B[0]));
    defparam ADV_B_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_0_preio (
            .PADOEN(N__23268),
            .PADOUT(N__23267),
            .PADIN(N__23266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11496),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_5_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_5_iopad (
            .OE(N__23259),
            .DIN(N__23258),
            .DOUT(N__23257),
            .PACKAGEPIN(TVP_VIDEO[5]));
    defparam TVP_VIDEO_pad_5_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_5_preio (
            .PADOEN(N__23259),
            .PADOUT(N__23258),
            .PADIN(N__23257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_2_iopad (
            .OE(N__23250),
            .DIN(N__23249),
            .DOUT(N__23248),
            .PACKAGEPIN(ADV_G[2]));
    defparam ADV_G_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_2_preio (
            .PADOEN(N__23250),
            .PADOUT(N__23249),
            .PADIN(N__23248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12638),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_VSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_VSYNC_pad_iopad (
            .OE(N__23241),
            .DIN(N__23240),
            .DOUT(N__23239),
            .PACKAGEPIN(ADV_VSYNC));
    defparam ADV_VSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_VSYNC_pad_preio (
            .PADOEN(N__23241),
            .PADOUT(N__23240),
            .PADIN(N__23239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20699),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5604 (
            .O(N__23222),
            .I(N__23219));
    LocalMux I__5603 (
            .O(N__23219),
            .I(N__23216));
    Span4Mux_v I__5602 (
            .O(N__23216),
            .I(N__23213));
    Span4Mux_v I__5601 (
            .O(N__23213),
            .I(N__23210));
    Sp12to4 I__5600 (
            .O(N__23210),
            .I(N__23207));
    Span12Mux_h I__5599 (
            .O(N__23207),
            .I(N__23204));
    Odrv12 I__5598 (
            .O(N__23204),
            .I(\line_buffer.n624 ));
    CascadeMux I__5597 (
            .O(N__23201),
            .I(N__23198));
    InMux I__5596 (
            .O(N__23198),
            .I(N__23195));
    LocalMux I__5595 (
            .O(N__23195),
            .I(N__23192));
    Span4Mux_v I__5594 (
            .O(N__23192),
            .I(N__23189));
    Sp12to4 I__5593 (
            .O(N__23189),
            .I(N__23186));
    Odrv12 I__5592 (
            .O(N__23186),
            .I(\line_buffer.n632 ));
    InMux I__5591 (
            .O(N__23183),
            .I(N__23180));
    LocalMux I__5590 (
            .O(N__23180),
            .I(N__23177));
    Odrv4 I__5589 (
            .O(N__23177),
            .I(\line_buffer.n3821 ));
    InMux I__5588 (
            .O(N__23174),
            .I(N__23171));
    LocalMux I__5587 (
            .O(N__23171),
            .I(N__23168));
    Span4Mux_v I__5586 (
            .O(N__23168),
            .I(N__23165));
    Span4Mux_h I__5585 (
            .O(N__23165),
            .I(N__23162));
    Odrv4 I__5584 (
            .O(N__23162),
            .I(\line_buffer.n593 ));
    CascadeMux I__5583 (
            .O(N__23159),
            .I(N__23156));
    InMux I__5582 (
            .O(N__23156),
            .I(N__23153));
    LocalMux I__5581 (
            .O(N__23153),
            .I(N__23150));
    Span12Mux_v I__5580 (
            .O(N__23150),
            .I(N__23147));
    Odrv12 I__5579 (
            .O(N__23147),
            .I(\line_buffer.n601 ));
    InMux I__5578 (
            .O(N__23144),
            .I(N__23138));
    InMux I__5577 (
            .O(N__23143),
            .I(N__23126));
    InMux I__5576 (
            .O(N__23142),
            .I(N__23122));
    InMux I__5575 (
            .O(N__23141),
            .I(N__23119));
    LocalMux I__5574 (
            .O(N__23138),
            .I(N__23114));
    InMux I__5573 (
            .O(N__23137),
            .I(N__23109));
    InMux I__5572 (
            .O(N__23136),
            .I(N__23109));
    InMux I__5571 (
            .O(N__23135),
            .I(N__23101));
    InMux I__5570 (
            .O(N__23134),
            .I(N__23101));
    InMux I__5569 (
            .O(N__23133),
            .I(N__23098));
    InMux I__5568 (
            .O(N__23132),
            .I(N__23095));
    InMux I__5567 (
            .O(N__23131),
            .I(N__23087));
    InMux I__5566 (
            .O(N__23130),
            .I(N__23084));
    InMux I__5565 (
            .O(N__23129),
            .I(N__23081));
    LocalMux I__5564 (
            .O(N__23126),
            .I(N__23078));
    InMux I__5563 (
            .O(N__23125),
            .I(N__23075));
    LocalMux I__5562 (
            .O(N__23122),
            .I(N__23072));
    LocalMux I__5561 (
            .O(N__23119),
            .I(N__23069));
    InMux I__5560 (
            .O(N__23118),
            .I(N__23066));
    InMux I__5559 (
            .O(N__23117),
            .I(N__23063));
    Span4Mux_v I__5558 (
            .O(N__23114),
            .I(N__23060));
    LocalMux I__5557 (
            .O(N__23109),
            .I(N__23057));
    InMux I__5556 (
            .O(N__23108),
            .I(N__23054));
    InMux I__5555 (
            .O(N__23107),
            .I(N__23051));
    InMux I__5554 (
            .O(N__23106),
            .I(N__23048));
    LocalMux I__5553 (
            .O(N__23101),
            .I(N__23045));
    LocalMux I__5552 (
            .O(N__23098),
            .I(N__23042));
    LocalMux I__5551 (
            .O(N__23095),
            .I(N__23039));
    InMux I__5550 (
            .O(N__23094),
            .I(N__23036));
    InMux I__5549 (
            .O(N__23093),
            .I(N__23033));
    InMux I__5548 (
            .O(N__23092),
            .I(N__23030));
    InMux I__5547 (
            .O(N__23091),
            .I(N__23025));
    InMux I__5546 (
            .O(N__23090),
            .I(N__23025));
    LocalMux I__5545 (
            .O(N__23087),
            .I(N__23016));
    LocalMux I__5544 (
            .O(N__23084),
            .I(N__23016));
    LocalMux I__5543 (
            .O(N__23081),
            .I(N__23016));
    Span4Mux_v I__5542 (
            .O(N__23078),
            .I(N__23016));
    LocalMux I__5541 (
            .O(N__23075),
            .I(N__23013));
    Span4Mux_v I__5540 (
            .O(N__23072),
            .I(N__23008));
    Span4Mux_v I__5539 (
            .O(N__23069),
            .I(N__23008));
    LocalMux I__5538 (
            .O(N__23066),
            .I(N__23005));
    LocalMux I__5537 (
            .O(N__23063),
            .I(N__23002));
    Span4Mux_v I__5536 (
            .O(N__23060),
            .I(N__22997));
    Span4Mux_v I__5535 (
            .O(N__23057),
            .I(N__22997));
    LocalMux I__5534 (
            .O(N__23054),
            .I(N__22994));
    LocalMux I__5533 (
            .O(N__23051),
            .I(N__22991));
    LocalMux I__5532 (
            .O(N__23048),
            .I(N__22986));
    Span4Mux_v I__5531 (
            .O(N__23045),
            .I(N__22986));
    Span4Mux_h I__5530 (
            .O(N__23042),
            .I(N__22981));
    Span4Mux_v I__5529 (
            .O(N__23039),
            .I(N__22981));
    LocalMux I__5528 (
            .O(N__23036),
            .I(N__22970));
    LocalMux I__5527 (
            .O(N__23033),
            .I(N__22970));
    LocalMux I__5526 (
            .O(N__23030),
            .I(N__22970));
    LocalMux I__5525 (
            .O(N__23025),
            .I(N__22970));
    Span4Mux_v I__5524 (
            .O(N__23016),
            .I(N__22970));
    Span4Mux_v I__5523 (
            .O(N__23013),
            .I(N__22965));
    Span4Mux_h I__5522 (
            .O(N__23008),
            .I(N__22965));
    Span4Mux_v I__5521 (
            .O(N__23005),
            .I(N__22960));
    Span4Mux_v I__5520 (
            .O(N__23002),
            .I(N__22960));
    Span4Mux_h I__5519 (
            .O(N__22997),
            .I(N__22955));
    Span4Mux_v I__5518 (
            .O(N__22994),
            .I(N__22955));
    Span4Mux_v I__5517 (
            .O(N__22991),
            .I(N__22946));
    Span4Mux_h I__5516 (
            .O(N__22986),
            .I(N__22946));
    Span4Mux_v I__5515 (
            .O(N__22981),
            .I(N__22946));
    Span4Mux_v I__5514 (
            .O(N__22970),
            .I(N__22946));
    Span4Mux_h I__5513 (
            .O(N__22965),
            .I(N__22943));
    Odrv4 I__5512 (
            .O(N__22960),
            .I(TX_ADDR_11));
    Odrv4 I__5511 (
            .O(N__22955),
            .I(TX_ADDR_11));
    Odrv4 I__5510 (
            .O(N__22946),
            .I(TX_ADDR_11));
    Odrv4 I__5509 (
            .O(N__22943),
            .I(TX_ADDR_11));
    InMux I__5508 (
            .O(N__22934),
            .I(N__22922));
    InMux I__5507 (
            .O(N__22933),
            .I(N__22915));
    InMux I__5506 (
            .O(N__22932),
            .I(N__22912));
    InMux I__5505 (
            .O(N__22931),
            .I(N__22909));
    InMux I__5504 (
            .O(N__22930),
            .I(N__22904));
    InMux I__5503 (
            .O(N__22929),
            .I(N__22901));
    InMux I__5502 (
            .O(N__22928),
            .I(N__22898));
    InMux I__5501 (
            .O(N__22927),
            .I(N__22893));
    InMux I__5500 (
            .O(N__22926),
            .I(N__22888));
    InMux I__5499 (
            .O(N__22925),
            .I(N__22885));
    LocalMux I__5498 (
            .O(N__22922),
            .I(N__22882));
    InMux I__5497 (
            .O(N__22921),
            .I(N__22873));
    InMux I__5496 (
            .O(N__22920),
            .I(N__22873));
    InMux I__5495 (
            .O(N__22919),
            .I(N__22873));
    InMux I__5494 (
            .O(N__22918),
            .I(N__22873));
    LocalMux I__5493 (
            .O(N__22915),
            .I(N__22867));
    LocalMux I__5492 (
            .O(N__22912),
            .I(N__22867));
    LocalMux I__5491 (
            .O(N__22909),
            .I(N__22861));
    InMux I__5490 (
            .O(N__22908),
            .I(N__22858));
    InMux I__5489 (
            .O(N__22907),
            .I(N__22855));
    LocalMux I__5488 (
            .O(N__22904),
            .I(N__22850));
    LocalMux I__5487 (
            .O(N__22901),
            .I(N__22850));
    LocalMux I__5486 (
            .O(N__22898),
            .I(N__22847));
    InMux I__5485 (
            .O(N__22897),
            .I(N__22842));
    InMux I__5484 (
            .O(N__22896),
            .I(N__22842));
    LocalMux I__5483 (
            .O(N__22893),
            .I(N__22839));
    InMux I__5482 (
            .O(N__22892),
            .I(N__22836));
    InMux I__5481 (
            .O(N__22891),
            .I(N__22833));
    LocalMux I__5480 (
            .O(N__22888),
            .I(N__22827));
    LocalMux I__5479 (
            .O(N__22885),
            .I(N__22827));
    Span4Mux_h I__5478 (
            .O(N__22882),
            .I(N__22824));
    LocalMux I__5477 (
            .O(N__22873),
            .I(N__22821));
    InMux I__5476 (
            .O(N__22872),
            .I(N__22818));
    Span4Mux_v I__5475 (
            .O(N__22867),
            .I(N__22815));
    InMux I__5474 (
            .O(N__22866),
            .I(N__22812));
    InMux I__5473 (
            .O(N__22865),
            .I(N__22807));
    InMux I__5472 (
            .O(N__22864),
            .I(N__22807));
    Span4Mux_h I__5471 (
            .O(N__22861),
            .I(N__22802));
    LocalMux I__5470 (
            .O(N__22858),
            .I(N__22802));
    LocalMux I__5469 (
            .O(N__22855),
            .I(N__22795));
    Span4Mux_h I__5468 (
            .O(N__22850),
            .I(N__22795));
    Span4Mux_h I__5467 (
            .O(N__22847),
            .I(N__22795));
    LocalMux I__5466 (
            .O(N__22842),
            .I(N__22788));
    Span4Mux_v I__5465 (
            .O(N__22839),
            .I(N__22788));
    LocalMux I__5464 (
            .O(N__22836),
            .I(N__22788));
    LocalMux I__5463 (
            .O(N__22833),
            .I(N__22785));
    InMux I__5462 (
            .O(N__22832),
            .I(N__22782));
    Span4Mux_v I__5461 (
            .O(N__22827),
            .I(N__22779));
    Span4Mux_v I__5460 (
            .O(N__22824),
            .I(N__22774));
    Span4Mux_h I__5459 (
            .O(N__22821),
            .I(N__22774));
    LocalMux I__5458 (
            .O(N__22818),
            .I(N__22765));
    Sp12to4 I__5457 (
            .O(N__22815),
            .I(N__22765));
    LocalMux I__5456 (
            .O(N__22812),
            .I(N__22765));
    LocalMux I__5455 (
            .O(N__22807),
            .I(N__22765));
    Span4Mux_h I__5454 (
            .O(N__22802),
            .I(N__22758));
    Span4Mux_v I__5453 (
            .O(N__22795),
            .I(N__22758));
    Span4Mux_h I__5452 (
            .O(N__22788),
            .I(N__22758));
    Span12Mux_h I__5451 (
            .O(N__22785),
            .I(N__22753));
    LocalMux I__5450 (
            .O(N__22782),
            .I(N__22753));
    Odrv4 I__5449 (
            .O(N__22779),
            .I(TX_ADDR_12));
    Odrv4 I__5448 (
            .O(N__22774),
            .I(TX_ADDR_12));
    Odrv12 I__5447 (
            .O(N__22765),
            .I(TX_ADDR_12));
    Odrv4 I__5446 (
            .O(N__22758),
            .I(TX_ADDR_12));
    Odrv12 I__5445 (
            .O(N__22753),
            .I(TX_ADDR_12));
    InMux I__5444 (
            .O(N__22742),
            .I(N__22739));
    LocalMux I__5443 (
            .O(N__22739),
            .I(N__22736));
    Span4Mux_v I__5442 (
            .O(N__22736),
            .I(N__22733));
    Span4Mux_h I__5441 (
            .O(N__22733),
            .I(N__22730));
    Span4Mux_v I__5440 (
            .O(N__22730),
            .I(N__22727));
    Odrv4 I__5439 (
            .O(N__22727),
            .I(\line_buffer.n496 ));
    CascadeMux I__5438 (
            .O(N__22724),
            .I(\line_buffer.n3809_cascade_ ));
    InMux I__5437 (
            .O(N__22721),
            .I(N__22718));
    LocalMux I__5436 (
            .O(N__22718),
            .I(N__22715));
    Span4Mux_v I__5435 (
            .O(N__22715),
            .I(N__22712));
    Span4Mux_v I__5434 (
            .O(N__22712),
            .I(N__22709));
    Span4Mux_h I__5433 (
            .O(N__22709),
            .I(N__22706));
    Odrv4 I__5432 (
            .O(N__22706),
            .I(\line_buffer.n504 ));
    InMux I__5431 (
            .O(N__22703),
            .I(N__22700));
    LocalMux I__5430 (
            .O(N__22700),
            .I(N__22697));
    Odrv12 I__5429 (
            .O(N__22697),
            .I(\line_buffer.n3812 ));
    SRMux I__5428 (
            .O(N__22694),
            .I(N__22690));
    SRMux I__5427 (
            .O(N__22693),
            .I(N__22687));
    LocalMux I__5426 (
            .O(N__22690),
            .I(N__22679));
    LocalMux I__5425 (
            .O(N__22687),
            .I(N__22679));
    SRMux I__5424 (
            .O(N__22686),
            .I(N__22676));
    SRMux I__5423 (
            .O(N__22685),
            .I(N__22673));
    SRMux I__5422 (
            .O(N__22684),
            .I(N__22668));
    Span4Mux_s2_v I__5421 (
            .O(N__22679),
            .I(N__22660));
    LocalMux I__5420 (
            .O(N__22676),
            .I(N__22660));
    LocalMux I__5419 (
            .O(N__22673),
            .I(N__22660));
    SRMux I__5418 (
            .O(N__22672),
            .I(N__22657));
    SRMux I__5417 (
            .O(N__22671),
            .I(N__22654));
    LocalMux I__5416 (
            .O(N__22668),
            .I(N__22649));
    SRMux I__5415 (
            .O(N__22667),
            .I(N__22646));
    Span4Mux_v I__5414 (
            .O(N__22660),
            .I(N__22638));
    LocalMux I__5413 (
            .O(N__22657),
            .I(N__22638));
    LocalMux I__5412 (
            .O(N__22654),
            .I(N__22638));
    SRMux I__5411 (
            .O(N__22653),
            .I(N__22635));
    SRMux I__5410 (
            .O(N__22652),
            .I(N__22632));
    Span4Mux_h I__5409 (
            .O(N__22649),
            .I(N__22628));
    LocalMux I__5408 (
            .O(N__22646),
            .I(N__22625));
    SRMux I__5407 (
            .O(N__22645),
            .I(N__22622));
    Span4Mux_v I__5406 (
            .O(N__22638),
            .I(N__22615));
    LocalMux I__5405 (
            .O(N__22635),
            .I(N__22615));
    LocalMux I__5404 (
            .O(N__22632),
            .I(N__22612));
    SRMux I__5403 (
            .O(N__22631),
            .I(N__22609));
    Span4Mux_v I__5402 (
            .O(N__22628),
            .I(N__22602));
    Span4Mux_h I__5401 (
            .O(N__22625),
            .I(N__22602));
    LocalMux I__5400 (
            .O(N__22622),
            .I(N__22599));
    SRMux I__5399 (
            .O(N__22621),
            .I(N__22596));
    SRMux I__5398 (
            .O(N__22620),
            .I(N__22593));
    Span4Mux_v I__5397 (
            .O(N__22615),
            .I(N__22585));
    Span4Mux_h I__5396 (
            .O(N__22612),
            .I(N__22585));
    LocalMux I__5395 (
            .O(N__22609),
            .I(N__22582));
    SRMux I__5394 (
            .O(N__22608),
            .I(N__22579));
    SRMux I__5393 (
            .O(N__22607),
            .I(N__22576));
    Span4Mux_v I__5392 (
            .O(N__22602),
            .I(N__22567));
    Span4Mux_h I__5391 (
            .O(N__22599),
            .I(N__22567));
    LocalMux I__5390 (
            .O(N__22596),
            .I(N__22567));
    LocalMux I__5389 (
            .O(N__22593),
            .I(N__22564));
    SRMux I__5388 (
            .O(N__22592),
            .I(N__22561));
    SRMux I__5387 (
            .O(N__22591),
            .I(N__22558));
    SRMux I__5386 (
            .O(N__22590),
            .I(N__22551));
    Span4Mux_v I__5385 (
            .O(N__22585),
            .I(N__22546));
    Span4Mux_h I__5384 (
            .O(N__22582),
            .I(N__22546));
    LocalMux I__5383 (
            .O(N__22579),
            .I(N__22541));
    LocalMux I__5382 (
            .O(N__22576),
            .I(N__22541));
    SRMux I__5381 (
            .O(N__22575),
            .I(N__22538));
    SRMux I__5380 (
            .O(N__22574),
            .I(N__22535));
    Span4Mux_v I__5379 (
            .O(N__22567),
            .I(N__22526));
    Span4Mux_h I__5378 (
            .O(N__22564),
            .I(N__22526));
    LocalMux I__5377 (
            .O(N__22561),
            .I(N__22526));
    LocalMux I__5376 (
            .O(N__22558),
            .I(N__22523));
    SRMux I__5375 (
            .O(N__22557),
            .I(N__22520));
    SRMux I__5374 (
            .O(N__22556),
            .I(N__22517));
    SRMux I__5373 (
            .O(N__22555),
            .I(N__22512));
    SRMux I__5372 (
            .O(N__22554),
            .I(N__22509));
    LocalMux I__5371 (
            .O(N__22551),
            .I(N__22503));
    Span4Mux_v I__5370 (
            .O(N__22546),
            .I(N__22494));
    Span4Mux_v I__5369 (
            .O(N__22541),
            .I(N__22494));
    LocalMux I__5368 (
            .O(N__22538),
            .I(N__22494));
    LocalMux I__5367 (
            .O(N__22535),
            .I(N__22494));
    SRMux I__5366 (
            .O(N__22534),
            .I(N__22491));
    SRMux I__5365 (
            .O(N__22533),
            .I(N__22488));
    Span4Mux_v I__5364 (
            .O(N__22526),
            .I(N__22481));
    Span4Mux_h I__5363 (
            .O(N__22523),
            .I(N__22481));
    LocalMux I__5362 (
            .O(N__22520),
            .I(N__22481));
    LocalMux I__5361 (
            .O(N__22517),
            .I(N__22478));
    SRMux I__5360 (
            .O(N__22516),
            .I(N__22475));
    SRMux I__5359 (
            .O(N__22515),
            .I(N__22472));
    LocalMux I__5358 (
            .O(N__22512),
            .I(N__22466));
    LocalMux I__5357 (
            .O(N__22509),
            .I(N__22466));
    SRMux I__5356 (
            .O(N__22508),
            .I(N__22463));
    IoInMux I__5355 (
            .O(N__22507),
            .I(N__22460));
    IoInMux I__5354 (
            .O(N__22506),
            .I(N__22457));
    Sp12to4 I__5353 (
            .O(N__22503),
            .I(N__22454));
    Span4Mux_v I__5352 (
            .O(N__22494),
            .I(N__22449));
    LocalMux I__5351 (
            .O(N__22491),
            .I(N__22449));
    LocalMux I__5350 (
            .O(N__22488),
            .I(N__22446));
    Span4Mux_v I__5349 (
            .O(N__22481),
            .I(N__22439));
    Span4Mux_h I__5348 (
            .O(N__22478),
            .I(N__22439));
    LocalMux I__5347 (
            .O(N__22475),
            .I(N__22439));
    LocalMux I__5346 (
            .O(N__22472),
            .I(N__22436));
    SRMux I__5345 (
            .O(N__22471),
            .I(N__22433));
    Span12Mux_s6_v I__5344 (
            .O(N__22466),
            .I(N__22427));
    LocalMux I__5343 (
            .O(N__22463),
            .I(N__22427));
    LocalMux I__5342 (
            .O(N__22460),
            .I(N__22422));
    LocalMux I__5341 (
            .O(N__22457),
            .I(N__22422));
    Span12Mux_v I__5340 (
            .O(N__22454),
            .I(N__22419));
    Span4Mux_v I__5339 (
            .O(N__22449),
            .I(N__22414));
    Span4Mux_h I__5338 (
            .O(N__22446),
            .I(N__22414));
    Span4Mux_v I__5337 (
            .O(N__22439),
            .I(N__22407));
    Span4Mux_h I__5336 (
            .O(N__22436),
            .I(N__22407));
    LocalMux I__5335 (
            .O(N__22433),
            .I(N__22407));
    SRMux I__5334 (
            .O(N__22432),
            .I(N__22404));
    Span12Mux_v I__5333 (
            .O(N__22427),
            .I(N__22401));
    Span4Mux_s2_v I__5332 (
            .O(N__22422),
            .I(N__22398));
    Span12Mux_h I__5331 (
            .O(N__22419),
            .I(N__22395));
    Sp12to4 I__5330 (
            .O(N__22414),
            .I(N__22392));
    Span4Mux_v I__5329 (
            .O(N__22407),
            .I(N__22387));
    LocalMux I__5328 (
            .O(N__22404),
            .I(N__22387));
    Span12Mux_v I__5327 (
            .O(N__22401),
            .I(N__22384));
    Span4Mux_h I__5326 (
            .O(N__22398),
            .I(N__22381));
    Span12Mux_v I__5325 (
            .O(N__22395),
            .I(N__22374));
    Span12Mux_h I__5324 (
            .O(N__22392),
            .I(N__22374));
    Sp12to4 I__5323 (
            .O(N__22387),
            .I(N__22374));
    Odrv12 I__5322 (
            .O(N__22384),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5321 (
            .O(N__22381),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__5320 (
            .O(N__22374),
            .I(CONSTANT_ONE_NET));
    InMux I__5319 (
            .O(N__22367),
            .I(N__22364));
    LocalMux I__5318 (
            .O(N__22364),
            .I(N__22361));
    Odrv12 I__5317 (
            .O(N__22361),
            .I(\line_buffer.n507 ));
    InMux I__5316 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__5315 (
            .O(N__22355),
            .I(N__22352));
    Span4Mux_v I__5314 (
            .O(N__22352),
            .I(N__22349));
    Sp12to4 I__5313 (
            .O(N__22349),
            .I(N__22346));
    Span12Mux_h I__5312 (
            .O(N__22346),
            .I(N__22343));
    Odrv12 I__5311 (
            .O(N__22343),
            .I(\line_buffer.n499 ));
    CascadeMux I__5310 (
            .O(N__22340),
            .I(N__22337));
    InMux I__5309 (
            .O(N__22337),
            .I(N__22334));
    LocalMux I__5308 (
            .O(N__22334),
            .I(N__22331));
    Odrv4 I__5307 (
            .O(N__22331),
            .I(\line_buffer.n3720 ));
    InMux I__5306 (
            .O(N__22328),
            .I(N__22325));
    LocalMux I__5305 (
            .O(N__22325),
            .I(N__22322));
    Span4Mux_v I__5304 (
            .O(N__22322),
            .I(N__22319));
    Span4Mux_h I__5303 (
            .O(N__22319),
            .I(N__22316));
    Odrv4 I__5302 (
            .O(N__22316),
            .I(\line_buffer.n592 ));
    CascadeMux I__5301 (
            .O(N__22313),
            .I(N__22310));
    InMux I__5300 (
            .O(N__22310),
            .I(N__22307));
    LocalMux I__5299 (
            .O(N__22307),
            .I(N__22304));
    Span4Mux_v I__5298 (
            .O(N__22304),
            .I(N__22301));
    Span4Mux_h I__5297 (
            .O(N__22301),
            .I(N__22298));
    Span4Mux_h I__5296 (
            .O(N__22298),
            .I(N__22295));
    Odrv4 I__5295 (
            .O(N__22295),
            .I(\line_buffer.n600 ));
    InMux I__5294 (
            .O(N__22292),
            .I(N__22289));
    LocalMux I__5293 (
            .O(N__22289),
            .I(N__22286));
    Sp12to4 I__5292 (
            .O(N__22286),
            .I(N__22283));
    Span12Mux_v I__5291 (
            .O(N__22283),
            .I(N__22280));
    Odrv12 I__5290 (
            .O(N__22280),
            .I(\line_buffer.n572 ));
    InMux I__5289 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__5288 (
            .O(N__22274),
            .I(N__22271));
    Span4Mux_v I__5287 (
            .O(N__22271),
            .I(N__22268));
    Span4Mux_h I__5286 (
            .O(N__22268),
            .I(N__22265));
    Odrv4 I__5285 (
            .O(N__22265),
            .I(\line_buffer.n564 ));
    InMux I__5284 (
            .O(N__22262),
            .I(N__22259));
    LocalMux I__5283 (
            .O(N__22259),
            .I(N__22256));
    Span4Mux_h I__5282 (
            .O(N__22256),
            .I(N__22253));
    Span4Mux_v I__5281 (
            .O(N__22253),
            .I(N__22250));
    Span4Mux_v I__5280 (
            .O(N__22250),
            .I(N__22247));
    Span4Mux_h I__5279 (
            .O(N__22247),
            .I(N__22244));
    Odrv4 I__5278 (
            .O(N__22244),
            .I(\line_buffer.n503 ));
    InMux I__5277 (
            .O(N__22241),
            .I(N__22238));
    LocalMux I__5276 (
            .O(N__22238),
            .I(\line_buffer.n3815 ));
    CascadeMux I__5275 (
            .O(N__22235),
            .I(N__22232));
    InMux I__5274 (
            .O(N__22232),
            .I(N__22229));
    LocalMux I__5273 (
            .O(N__22229),
            .I(N__22226));
    Span4Mux_v I__5272 (
            .O(N__22226),
            .I(N__22223));
    Span4Mux_h I__5271 (
            .O(N__22223),
            .I(N__22220));
    Span4Mux_v I__5270 (
            .O(N__22220),
            .I(N__22217));
    Span4Mux_v I__5269 (
            .O(N__22217),
            .I(N__22214));
    Odrv4 I__5268 (
            .O(N__22214),
            .I(\line_buffer.n495 ));
    InMux I__5267 (
            .O(N__22211),
            .I(N__22208));
    LocalMux I__5266 (
            .O(N__22208),
            .I(N__22205));
    Sp12to4 I__5265 (
            .O(N__22205),
            .I(N__22202));
    Span12Mux_v I__5264 (
            .O(N__22202),
            .I(N__22199));
    Odrv12 I__5263 (
            .O(N__22199),
            .I(\line_buffer.n568 ));
    CascadeMux I__5262 (
            .O(N__22196),
            .I(N__22193));
    InMux I__5261 (
            .O(N__22193),
            .I(N__22190));
    LocalMux I__5260 (
            .O(N__22190),
            .I(N__22187));
    Span4Mux_h I__5259 (
            .O(N__22187),
            .I(N__22184));
    Span4Mux_v I__5258 (
            .O(N__22184),
            .I(N__22181));
    Odrv4 I__5257 (
            .O(N__22181),
            .I(\line_buffer.n560 ));
    CascadeMux I__5256 (
            .O(N__22178),
            .I(\line_buffer.n3824_cascade_ ));
    InMux I__5255 (
            .O(N__22175),
            .I(N__22172));
    LocalMux I__5254 (
            .O(N__22172),
            .I(\line_buffer.n3818 ));
    InMux I__5253 (
            .O(N__22169),
            .I(N__22166));
    LocalMux I__5252 (
            .O(N__22166),
            .I(N__22163));
    Odrv12 I__5251 (
            .O(N__22163),
            .I(TX_DATA_0));
    ClkMux I__5250 (
            .O(N__22160),
            .I(N__22155));
    ClkMux I__5249 (
            .O(N__22159),
            .I(N__22152));
    ClkMux I__5248 (
            .O(N__22158),
            .I(N__22146));
    LocalMux I__5247 (
            .O(N__22155),
            .I(N__22134));
    LocalMux I__5246 (
            .O(N__22152),
            .I(N__22131));
    ClkMux I__5245 (
            .O(N__22151),
            .I(N__22128));
    ClkMux I__5244 (
            .O(N__22150),
            .I(N__22125));
    ClkMux I__5243 (
            .O(N__22149),
            .I(N__22120));
    LocalMux I__5242 (
            .O(N__22146),
            .I(N__22114));
    ClkMux I__5241 (
            .O(N__22145),
            .I(N__22111));
    ClkMux I__5240 (
            .O(N__22144),
            .I(N__22108));
    ClkMux I__5239 (
            .O(N__22143),
            .I(N__22105));
    ClkMux I__5238 (
            .O(N__22142),
            .I(N__22100));
    ClkMux I__5237 (
            .O(N__22141),
            .I(N__22096));
    ClkMux I__5236 (
            .O(N__22140),
            .I(N__22092));
    ClkMux I__5235 (
            .O(N__22139),
            .I(N__22081));
    ClkMux I__5234 (
            .O(N__22138),
            .I(N__22078));
    ClkMux I__5233 (
            .O(N__22137),
            .I(N__22074));
    Span4Mux_s2_v I__5232 (
            .O(N__22134),
            .I(N__22063));
    Span4Mux_h I__5231 (
            .O(N__22131),
            .I(N__22063));
    LocalMux I__5230 (
            .O(N__22128),
            .I(N__22063));
    LocalMux I__5229 (
            .O(N__22125),
            .I(N__22060));
    ClkMux I__5228 (
            .O(N__22124),
            .I(N__22057));
    ClkMux I__5227 (
            .O(N__22123),
            .I(N__22054));
    LocalMux I__5226 (
            .O(N__22120),
            .I(N__22049));
    ClkMux I__5225 (
            .O(N__22119),
            .I(N__22046));
    ClkMux I__5224 (
            .O(N__22118),
            .I(N__22043));
    ClkMux I__5223 (
            .O(N__22117),
            .I(N__22038));
    Span4Mux_h I__5222 (
            .O(N__22114),
            .I(N__22032));
    LocalMux I__5221 (
            .O(N__22111),
            .I(N__22032));
    LocalMux I__5220 (
            .O(N__22108),
            .I(N__22027));
    LocalMux I__5219 (
            .O(N__22105),
            .I(N__22027));
    ClkMux I__5218 (
            .O(N__22104),
            .I(N__22024));
    ClkMux I__5217 (
            .O(N__22103),
            .I(N__22021));
    LocalMux I__5216 (
            .O(N__22100),
            .I(N__22018));
    ClkMux I__5215 (
            .O(N__22099),
            .I(N__22015));
    LocalMux I__5214 (
            .O(N__22096),
            .I(N__22011));
    ClkMux I__5213 (
            .O(N__22095),
            .I(N__22008));
    LocalMux I__5212 (
            .O(N__22092),
            .I(N__22004));
    ClkMux I__5211 (
            .O(N__22091),
            .I(N__22001));
    ClkMux I__5210 (
            .O(N__22090),
            .I(N__21998));
    ClkMux I__5209 (
            .O(N__22089),
            .I(N__21994));
    ClkMux I__5208 (
            .O(N__22088),
            .I(N__21991));
    ClkMux I__5207 (
            .O(N__22087),
            .I(N__21988));
    ClkMux I__5206 (
            .O(N__22086),
            .I(N__21984));
    ClkMux I__5205 (
            .O(N__22085),
            .I(N__21980));
    ClkMux I__5204 (
            .O(N__22084),
            .I(N__21977));
    LocalMux I__5203 (
            .O(N__22081),
            .I(N__21973));
    LocalMux I__5202 (
            .O(N__22078),
            .I(N__21970));
    ClkMux I__5201 (
            .O(N__22077),
            .I(N__21967));
    LocalMux I__5200 (
            .O(N__22074),
            .I(N__21963));
    ClkMux I__5199 (
            .O(N__22073),
            .I(N__21960));
    ClkMux I__5198 (
            .O(N__22072),
            .I(N__21953));
    ClkMux I__5197 (
            .O(N__22071),
            .I(N__21950));
    ClkMux I__5196 (
            .O(N__22070),
            .I(N__21943));
    Span4Mux_v I__5195 (
            .O(N__22063),
            .I(N__21936));
    Span4Mux_h I__5194 (
            .O(N__22060),
            .I(N__21936));
    LocalMux I__5193 (
            .O(N__22057),
            .I(N__21936));
    LocalMux I__5192 (
            .O(N__22054),
            .I(N__21933));
    ClkMux I__5191 (
            .O(N__22053),
            .I(N__21930));
    ClkMux I__5190 (
            .O(N__22052),
            .I(N__21927));
    Span4Mux_v I__5189 (
            .O(N__22049),
            .I(N__21921));
    LocalMux I__5188 (
            .O(N__22046),
            .I(N__21918));
    LocalMux I__5187 (
            .O(N__22043),
            .I(N__21915));
    ClkMux I__5186 (
            .O(N__22042),
            .I(N__21912));
    ClkMux I__5185 (
            .O(N__22041),
            .I(N__21909));
    LocalMux I__5184 (
            .O(N__22038),
            .I(N__21905));
    ClkMux I__5183 (
            .O(N__22037),
            .I(N__21902));
    Span4Mux_v I__5182 (
            .O(N__22032),
            .I(N__21893));
    Span4Mux_h I__5181 (
            .O(N__22027),
            .I(N__21893));
    LocalMux I__5180 (
            .O(N__22024),
            .I(N__21893));
    LocalMux I__5179 (
            .O(N__22021),
            .I(N__21893));
    Span4Mux_v I__5178 (
            .O(N__22018),
            .I(N__21888));
    LocalMux I__5177 (
            .O(N__22015),
            .I(N__21888));
    ClkMux I__5176 (
            .O(N__22014),
            .I(N__21885));
    Span4Mux_v I__5175 (
            .O(N__22011),
            .I(N__21880));
    LocalMux I__5174 (
            .O(N__22008),
            .I(N__21880));
    ClkMux I__5173 (
            .O(N__22007),
            .I(N__21877));
    Span4Mux_v I__5172 (
            .O(N__22004),
            .I(N__21870));
    LocalMux I__5171 (
            .O(N__22001),
            .I(N__21870));
    LocalMux I__5170 (
            .O(N__21998),
            .I(N__21867));
    ClkMux I__5169 (
            .O(N__21997),
            .I(N__21864));
    LocalMux I__5168 (
            .O(N__21994),
            .I(N__21859));
    LocalMux I__5167 (
            .O(N__21991),
            .I(N__21859));
    LocalMux I__5166 (
            .O(N__21988),
            .I(N__21856));
    ClkMux I__5165 (
            .O(N__21987),
            .I(N__21853));
    LocalMux I__5164 (
            .O(N__21984),
            .I(N__21850));
    ClkMux I__5163 (
            .O(N__21983),
            .I(N__21847));
    LocalMux I__5162 (
            .O(N__21980),
            .I(N__21842));
    LocalMux I__5161 (
            .O(N__21977),
            .I(N__21842));
    ClkMux I__5160 (
            .O(N__21976),
            .I(N__21839));
    Span4Mux_h I__5159 (
            .O(N__21973),
            .I(N__21832));
    Span4Mux_h I__5158 (
            .O(N__21970),
            .I(N__21832));
    LocalMux I__5157 (
            .O(N__21967),
            .I(N__21832));
    ClkMux I__5156 (
            .O(N__21966),
            .I(N__21829));
    Span4Mux_h I__5155 (
            .O(N__21963),
            .I(N__21824));
    LocalMux I__5154 (
            .O(N__21960),
            .I(N__21821));
    ClkMux I__5153 (
            .O(N__21959),
            .I(N__21818));
    ClkMux I__5152 (
            .O(N__21958),
            .I(N__21813));
    ClkMux I__5151 (
            .O(N__21957),
            .I(N__21810));
    IoInMux I__5150 (
            .O(N__21956),
            .I(N__21805));
    LocalMux I__5149 (
            .O(N__21953),
            .I(N__21799));
    LocalMux I__5148 (
            .O(N__21950),
            .I(N__21799));
    ClkMux I__5147 (
            .O(N__21949),
            .I(N__21796));
    ClkMux I__5146 (
            .O(N__21948),
            .I(N__21793));
    ClkMux I__5145 (
            .O(N__21947),
            .I(N__21790));
    ClkMux I__5144 (
            .O(N__21946),
            .I(N__21787));
    LocalMux I__5143 (
            .O(N__21943),
            .I(N__21783));
    Span4Mux_v I__5142 (
            .O(N__21936),
            .I(N__21775));
    Span4Mux_h I__5141 (
            .O(N__21933),
            .I(N__21775));
    LocalMux I__5140 (
            .O(N__21930),
            .I(N__21775));
    LocalMux I__5139 (
            .O(N__21927),
            .I(N__21772));
    ClkMux I__5138 (
            .O(N__21926),
            .I(N__21769));
    ClkMux I__5137 (
            .O(N__21925),
            .I(N__21766));
    ClkMux I__5136 (
            .O(N__21924),
            .I(N__21762));
    Span4Mux_h I__5135 (
            .O(N__21921),
            .I(N__21753));
    Span4Mux_h I__5134 (
            .O(N__21918),
            .I(N__21753));
    Span4Mux_v I__5133 (
            .O(N__21915),
            .I(N__21753));
    LocalMux I__5132 (
            .O(N__21912),
            .I(N__21753));
    LocalMux I__5131 (
            .O(N__21909),
            .I(N__21750));
    ClkMux I__5130 (
            .O(N__21908),
            .I(N__21747));
    Span4Mux_h I__5129 (
            .O(N__21905),
            .I(N__21742));
    LocalMux I__5128 (
            .O(N__21902),
            .I(N__21742));
    Span4Mux_v I__5127 (
            .O(N__21893),
            .I(N__21735));
    Span4Mux_v I__5126 (
            .O(N__21888),
            .I(N__21735));
    LocalMux I__5125 (
            .O(N__21885),
            .I(N__21735));
    Span4Mux_h I__5124 (
            .O(N__21880),
            .I(N__21730));
    LocalMux I__5123 (
            .O(N__21877),
            .I(N__21730));
    ClkMux I__5122 (
            .O(N__21876),
            .I(N__21727));
    ClkMux I__5121 (
            .O(N__21875),
            .I(N__21724));
    Span4Mux_v I__5120 (
            .O(N__21870),
            .I(N__21720));
    Span4Mux_v I__5119 (
            .O(N__21867),
            .I(N__21715));
    LocalMux I__5118 (
            .O(N__21864),
            .I(N__21715));
    Span4Mux_v I__5117 (
            .O(N__21859),
            .I(N__21708));
    Span4Mux_h I__5116 (
            .O(N__21856),
            .I(N__21708));
    LocalMux I__5115 (
            .O(N__21853),
            .I(N__21708));
    Span4Mux_v I__5114 (
            .O(N__21850),
            .I(N__21703));
    LocalMux I__5113 (
            .O(N__21847),
            .I(N__21703));
    Span4Mux_v I__5112 (
            .O(N__21842),
            .I(N__21698));
    LocalMux I__5111 (
            .O(N__21839),
            .I(N__21698));
    Span4Mux_h I__5110 (
            .O(N__21832),
            .I(N__21693));
    LocalMux I__5109 (
            .O(N__21829),
            .I(N__21693));
    ClkMux I__5108 (
            .O(N__21828),
            .I(N__21690));
    ClkMux I__5107 (
            .O(N__21827),
            .I(N__21687));
    Span4Mux_v I__5106 (
            .O(N__21824),
            .I(N__21677));
    Span4Mux_h I__5105 (
            .O(N__21821),
            .I(N__21677));
    LocalMux I__5104 (
            .O(N__21818),
            .I(N__21674));
    ClkMux I__5103 (
            .O(N__21817),
            .I(N__21671));
    ClkMux I__5102 (
            .O(N__21816),
            .I(N__21668));
    LocalMux I__5101 (
            .O(N__21813),
            .I(N__21662));
    LocalMux I__5100 (
            .O(N__21810),
            .I(N__21662));
    ClkMux I__5099 (
            .O(N__21809),
            .I(N__21659));
    ClkMux I__5098 (
            .O(N__21808),
            .I(N__21656));
    LocalMux I__5097 (
            .O(N__21805),
            .I(N__21653));
    ClkMux I__5096 (
            .O(N__21804),
            .I(N__21650));
    Span4Mux_v I__5095 (
            .O(N__21799),
            .I(N__21641));
    LocalMux I__5094 (
            .O(N__21796),
            .I(N__21641));
    LocalMux I__5093 (
            .O(N__21793),
            .I(N__21641));
    LocalMux I__5092 (
            .O(N__21790),
            .I(N__21641));
    LocalMux I__5091 (
            .O(N__21787),
            .I(N__21638));
    ClkMux I__5090 (
            .O(N__21786),
            .I(N__21635));
    Span4Mux_v I__5089 (
            .O(N__21783),
            .I(N__21632));
    ClkMux I__5088 (
            .O(N__21782),
            .I(N__21629));
    Span4Mux_v I__5087 (
            .O(N__21775),
            .I(N__21621));
    Span4Mux_h I__5086 (
            .O(N__21772),
            .I(N__21621));
    LocalMux I__5085 (
            .O(N__21769),
            .I(N__21621));
    LocalMux I__5084 (
            .O(N__21766),
            .I(N__21618));
    ClkMux I__5083 (
            .O(N__21765),
            .I(N__21615));
    LocalMux I__5082 (
            .O(N__21762),
            .I(N__21612));
    Span4Mux_v I__5081 (
            .O(N__21753),
            .I(N__21609));
    Span4Mux_v I__5080 (
            .O(N__21750),
            .I(N__21604));
    LocalMux I__5079 (
            .O(N__21747),
            .I(N__21604));
    Span4Mux_v I__5078 (
            .O(N__21742),
            .I(N__21593));
    Span4Mux_h I__5077 (
            .O(N__21735),
            .I(N__21593));
    Span4Mux_h I__5076 (
            .O(N__21730),
            .I(N__21593));
    LocalMux I__5075 (
            .O(N__21727),
            .I(N__21593));
    LocalMux I__5074 (
            .O(N__21724),
            .I(N__21593));
    ClkMux I__5073 (
            .O(N__21723),
            .I(N__21590));
    Span4Mux_v I__5072 (
            .O(N__21720),
            .I(N__21585));
    Span4Mux_v I__5071 (
            .O(N__21715),
            .I(N__21585));
    Span4Mux_h I__5070 (
            .O(N__21708),
            .I(N__21572));
    Span4Mux_h I__5069 (
            .O(N__21703),
            .I(N__21572));
    Span4Mux_v I__5068 (
            .O(N__21698),
            .I(N__21572));
    Span4Mux_v I__5067 (
            .O(N__21693),
            .I(N__21572));
    LocalMux I__5066 (
            .O(N__21690),
            .I(N__21572));
    LocalMux I__5065 (
            .O(N__21687),
            .I(N__21572));
    ClkMux I__5064 (
            .O(N__21686),
            .I(N__21569));
    ClkMux I__5063 (
            .O(N__21685),
            .I(N__21566));
    ClkMux I__5062 (
            .O(N__21684),
            .I(N__21563));
    ClkMux I__5061 (
            .O(N__21683),
            .I(N__21560));
    ClkMux I__5060 (
            .O(N__21682),
            .I(N__21554));
    Span4Mux_v I__5059 (
            .O(N__21677),
            .I(N__21548));
    Span4Mux_h I__5058 (
            .O(N__21674),
            .I(N__21548));
    LocalMux I__5057 (
            .O(N__21671),
            .I(N__21545));
    LocalMux I__5056 (
            .O(N__21668),
            .I(N__21542));
    ClkMux I__5055 (
            .O(N__21667),
            .I(N__21539));
    Span4Mux_v I__5054 (
            .O(N__21662),
            .I(N__21532));
    LocalMux I__5053 (
            .O(N__21659),
            .I(N__21532));
    LocalMux I__5052 (
            .O(N__21656),
            .I(N__21532));
    Span4Mux_s2_v I__5051 (
            .O(N__21653),
            .I(N__21529));
    LocalMux I__5050 (
            .O(N__21650),
            .I(N__21526));
    Span4Mux_v I__5049 (
            .O(N__21641),
            .I(N__21523));
    Span4Mux_v I__5048 (
            .O(N__21638),
            .I(N__21518));
    LocalMux I__5047 (
            .O(N__21635),
            .I(N__21518));
    Span4Mux_v I__5046 (
            .O(N__21632),
            .I(N__21513));
    LocalMux I__5045 (
            .O(N__21629),
            .I(N__21513));
    ClkMux I__5044 (
            .O(N__21628),
            .I(N__21510));
    Span4Mux_v I__5043 (
            .O(N__21621),
            .I(N__21502));
    Span4Mux_h I__5042 (
            .O(N__21618),
            .I(N__21502));
    LocalMux I__5041 (
            .O(N__21615),
            .I(N__21502));
    Span4Mux_v I__5040 (
            .O(N__21612),
            .I(N__21499));
    Span4Mux_v I__5039 (
            .O(N__21609),
            .I(N__21496));
    Span4Mux_v I__5038 (
            .O(N__21604),
            .I(N__21491));
    Span4Mux_v I__5037 (
            .O(N__21593),
            .I(N__21491));
    LocalMux I__5036 (
            .O(N__21590),
            .I(N__21487));
    Span4Mux_v I__5035 (
            .O(N__21585),
            .I(N__21480));
    Span4Mux_h I__5034 (
            .O(N__21572),
            .I(N__21480));
    LocalMux I__5033 (
            .O(N__21569),
            .I(N__21480));
    LocalMux I__5032 (
            .O(N__21566),
            .I(N__21476));
    LocalMux I__5031 (
            .O(N__21563),
            .I(N__21471));
    LocalMux I__5030 (
            .O(N__21560),
            .I(N__21471));
    ClkMux I__5029 (
            .O(N__21559),
            .I(N__21468));
    ClkMux I__5028 (
            .O(N__21558),
            .I(N__21465));
    ClkMux I__5027 (
            .O(N__21557),
            .I(N__21462));
    LocalMux I__5026 (
            .O(N__21554),
            .I(N__21459));
    ClkMux I__5025 (
            .O(N__21553),
            .I(N__21456));
    Span4Mux_v I__5024 (
            .O(N__21548),
            .I(N__21447));
    Span4Mux_h I__5023 (
            .O(N__21545),
            .I(N__21447));
    Span4Mux_h I__5022 (
            .O(N__21542),
            .I(N__21447));
    LocalMux I__5021 (
            .O(N__21539),
            .I(N__21447));
    Span4Mux_v I__5020 (
            .O(N__21532),
            .I(N__21439));
    Span4Mux_h I__5019 (
            .O(N__21529),
            .I(N__21439));
    Span4Mux_s2_v I__5018 (
            .O(N__21526),
            .I(N__21439));
    Span4Mux_v I__5017 (
            .O(N__21523),
            .I(N__21434));
    Span4Mux_v I__5016 (
            .O(N__21518),
            .I(N__21434));
    Span4Mux_v I__5015 (
            .O(N__21513),
            .I(N__21429));
    LocalMux I__5014 (
            .O(N__21510),
            .I(N__21429));
    ClkMux I__5013 (
            .O(N__21509),
            .I(N__21426));
    Span4Mux_v I__5012 (
            .O(N__21502),
            .I(N__21423));
    Span4Mux_v I__5011 (
            .O(N__21499),
            .I(N__21416));
    Span4Mux_h I__5010 (
            .O(N__21496),
            .I(N__21416));
    Span4Mux_v I__5009 (
            .O(N__21491),
            .I(N__21416));
    ClkMux I__5008 (
            .O(N__21490),
            .I(N__21413));
    Span4Mux_v I__5007 (
            .O(N__21487),
            .I(N__21408));
    Span4Mux_v I__5006 (
            .O(N__21480),
            .I(N__21408));
    ClkMux I__5005 (
            .O(N__21479),
            .I(N__21405));
    Span4Mux_v I__5004 (
            .O(N__21476),
            .I(N__21394));
    Span4Mux_v I__5003 (
            .O(N__21471),
            .I(N__21394));
    LocalMux I__5002 (
            .O(N__21468),
            .I(N__21394));
    LocalMux I__5001 (
            .O(N__21465),
            .I(N__21394));
    LocalMux I__5000 (
            .O(N__21462),
            .I(N__21394));
    Span12Mux_h I__4999 (
            .O(N__21459),
            .I(N__21391));
    LocalMux I__4998 (
            .O(N__21456),
            .I(N__21388));
    Span4Mux_h I__4997 (
            .O(N__21447),
            .I(N__21385));
    ClkMux I__4996 (
            .O(N__21446),
            .I(N__21382));
    Span4Mux_h I__4995 (
            .O(N__21439),
            .I(N__21379));
    Span4Mux_v I__4994 (
            .O(N__21434),
            .I(N__21376));
    Span4Mux_v I__4993 (
            .O(N__21429),
            .I(N__21371));
    LocalMux I__4992 (
            .O(N__21426),
            .I(N__21371));
    Sp12to4 I__4991 (
            .O(N__21423),
            .I(N__21366));
    Sp12to4 I__4990 (
            .O(N__21416),
            .I(N__21366));
    LocalMux I__4989 (
            .O(N__21413),
            .I(N__21361));
    Sp12to4 I__4988 (
            .O(N__21408),
            .I(N__21361));
    LocalMux I__4987 (
            .O(N__21405),
            .I(N__21356));
    Sp12to4 I__4986 (
            .O(N__21394),
            .I(N__21356));
    Span12Mux_v I__4985 (
            .O(N__21391),
            .I(N__21349));
    Span12Mux_h I__4984 (
            .O(N__21388),
            .I(N__21349));
    Sp12to4 I__4983 (
            .O(N__21385),
            .I(N__21349));
    LocalMux I__4982 (
            .O(N__21382),
            .I(N__21346));
    IoSpan4Mux I__4981 (
            .O(N__21379),
            .I(N__21343));
    Span4Mux_v I__4980 (
            .O(N__21376),
            .I(N__21340));
    Span4Mux_h I__4979 (
            .O(N__21371),
            .I(N__21337));
    Span12Mux_h I__4978 (
            .O(N__21366),
            .I(N__21330));
    Span12Mux_h I__4977 (
            .O(N__21361),
            .I(N__21330));
    Span12Mux_v I__4976 (
            .O(N__21356),
            .I(N__21330));
    Span12Mux_v I__4975 (
            .O(N__21349),
            .I(N__21325));
    Span12Mux_h I__4974 (
            .O(N__21346),
            .I(N__21325));
    IoSpan4Mux I__4973 (
            .O(N__21343),
            .I(N__21322));
    Span4Mux_h I__4972 (
            .O(N__21340),
            .I(N__21317));
    Span4Mux_h I__4971 (
            .O(N__21337),
            .I(N__21317));
    Odrv12 I__4970 (
            .O(N__21330),
            .I(ADV_CLK_c));
    Odrv12 I__4969 (
            .O(N__21325),
            .I(ADV_CLK_c));
    Odrv4 I__4968 (
            .O(N__21322),
            .I(ADV_CLK_c));
    Odrv4 I__4967 (
            .O(N__21317),
            .I(ADV_CLK_c));
    InMux I__4966 (
            .O(N__21308),
            .I(N__21305));
    LocalMux I__4965 (
            .O(N__21305),
            .I(N__21302));
    Span12Mux_v I__4964 (
            .O(N__21302),
            .I(N__21299));
    Odrv12 I__4963 (
            .O(N__21299),
            .I(\line_buffer.n3699 ));
    IoInMux I__4962 (
            .O(N__21296),
            .I(N__21292));
    CascadeMux I__4961 (
            .O(N__21295),
            .I(N__21285));
    LocalMux I__4960 (
            .O(N__21292),
            .I(N__21281));
    InMux I__4959 (
            .O(N__21291),
            .I(N__21278));
    CascadeMux I__4958 (
            .O(N__21290),
            .I(N__21273));
    CascadeMux I__4957 (
            .O(N__21289),
            .I(N__21268));
    InMux I__4956 (
            .O(N__21288),
            .I(N__21265));
    InMux I__4955 (
            .O(N__21285),
            .I(N__21262));
    InMux I__4954 (
            .O(N__21284),
            .I(N__21258));
    Span4Mux_s3_h I__4953 (
            .O(N__21281),
            .I(N__21254));
    LocalMux I__4952 (
            .O(N__21278),
            .I(N__21250));
    InMux I__4951 (
            .O(N__21277),
            .I(N__21247));
    InMux I__4950 (
            .O(N__21276),
            .I(N__21242));
    InMux I__4949 (
            .O(N__21273),
            .I(N__21242));
    InMux I__4948 (
            .O(N__21272),
            .I(N__21235));
    InMux I__4947 (
            .O(N__21271),
            .I(N__21235));
    InMux I__4946 (
            .O(N__21268),
            .I(N__21235));
    LocalMux I__4945 (
            .O(N__21265),
            .I(N__21230));
    LocalMux I__4944 (
            .O(N__21262),
            .I(N__21230));
    InMux I__4943 (
            .O(N__21261),
            .I(N__21227));
    LocalMux I__4942 (
            .O(N__21258),
            .I(N__21224));
    InMux I__4941 (
            .O(N__21257),
            .I(N__21221));
    Span4Mux_v I__4940 (
            .O(N__21254),
            .I(N__21218));
    InMux I__4939 (
            .O(N__21253),
            .I(N__21215));
    Span4Mux_v I__4938 (
            .O(N__21250),
            .I(N__21211));
    LocalMux I__4937 (
            .O(N__21247),
            .I(N__21208));
    LocalMux I__4936 (
            .O(N__21242),
            .I(N__21203));
    LocalMux I__4935 (
            .O(N__21235),
            .I(N__21203));
    Span4Mux_h I__4934 (
            .O(N__21230),
            .I(N__21200));
    LocalMux I__4933 (
            .O(N__21227),
            .I(N__21197));
    Span4Mux_v I__4932 (
            .O(N__21224),
            .I(N__21192));
    LocalMux I__4931 (
            .O(N__21221),
            .I(N__21192));
    Sp12to4 I__4930 (
            .O(N__21218),
            .I(N__21189));
    LocalMux I__4929 (
            .O(N__21215),
            .I(N__21186));
    InMux I__4928 (
            .O(N__21214),
            .I(N__21183));
    Span4Mux_h I__4927 (
            .O(N__21211),
            .I(N__21176));
    Span4Mux_v I__4926 (
            .O(N__21208),
            .I(N__21176));
    Span4Mux_v I__4925 (
            .O(N__21203),
            .I(N__21176));
    Span4Mux_h I__4924 (
            .O(N__21200),
            .I(N__21173));
    Span4Mux_v I__4923 (
            .O(N__21197),
            .I(N__21168));
    Span4Mux_v I__4922 (
            .O(N__21192),
            .I(N__21168));
    Odrv12 I__4921 (
            .O(N__21189),
            .I(DEBUG_c_2));
    Odrv4 I__4920 (
            .O(N__21186),
            .I(DEBUG_c_2));
    LocalMux I__4919 (
            .O(N__21183),
            .I(DEBUG_c_2));
    Odrv4 I__4918 (
            .O(N__21176),
            .I(DEBUG_c_2));
    Odrv4 I__4917 (
            .O(N__21173),
            .I(DEBUG_c_2));
    Odrv4 I__4916 (
            .O(N__21168),
            .I(DEBUG_c_2));
    InMux I__4915 (
            .O(N__21155),
            .I(N__21152));
    LocalMux I__4914 (
            .O(N__21152),
            .I(N__21149));
    Odrv4 I__4913 (
            .O(N__21149),
            .I(\line_buffer.n3797 ));
    InMux I__4912 (
            .O(N__21146),
            .I(N__21143));
    LocalMux I__4911 (
            .O(N__21143),
            .I(N__21140));
    Span4Mux_v I__4910 (
            .O(N__21140),
            .I(N__21137));
    Span4Mux_v I__4909 (
            .O(N__21137),
            .I(N__21134));
    Sp12to4 I__4908 (
            .O(N__21134),
            .I(N__21131));
    Odrv12 I__4907 (
            .O(N__21131),
            .I(\line_buffer.n636 ));
    InMux I__4906 (
            .O(N__21128),
            .I(N__21125));
    LocalMux I__4905 (
            .O(N__21125),
            .I(N__21122));
    Span4Mux_h I__4904 (
            .O(N__21122),
            .I(N__21119));
    Span4Mux_v I__4903 (
            .O(N__21119),
            .I(N__21116));
    Span4Mux_v I__4902 (
            .O(N__21116),
            .I(N__21113));
    Span4Mux_h I__4901 (
            .O(N__21113),
            .I(N__21110));
    Odrv4 I__4900 (
            .O(N__21110),
            .I(\line_buffer.n628 ));
    InMux I__4899 (
            .O(N__21107),
            .I(N__21104));
    LocalMux I__4898 (
            .O(N__21104),
            .I(N__21101));
    Odrv4 I__4897 (
            .O(N__21101),
            .I(\line_buffer.n3700 ));
    InMux I__4896 (
            .O(N__21098),
            .I(N__21093));
    InMux I__4895 (
            .O(N__21097),
            .I(N__21088));
    InMux I__4894 (
            .O(N__21096),
            .I(N__21088));
    LocalMux I__4893 (
            .O(N__21093),
            .I(\receive_module.rx_counter.X_7 ));
    LocalMux I__4892 (
            .O(N__21088),
            .I(\receive_module.rx_counter.X_7 ));
    InMux I__4891 (
            .O(N__21083),
            .I(\receive_module.rx_counter.n3363 ));
    InMux I__4890 (
            .O(N__21080),
            .I(N__21076));
    InMux I__4889 (
            .O(N__21079),
            .I(N__21073));
    LocalMux I__4888 (
            .O(N__21076),
            .I(\receive_module.rx_counter.X_8 ));
    LocalMux I__4887 (
            .O(N__21073),
            .I(\receive_module.rx_counter.X_8 ));
    InMux I__4886 (
            .O(N__21068),
            .I(bfn_17_10_0_));
    InMux I__4885 (
            .O(N__21065),
            .I(\receive_module.rx_counter.n3365 ));
    InMux I__4884 (
            .O(N__21062),
            .I(N__21058));
    InMux I__4883 (
            .O(N__21061),
            .I(N__21055));
    LocalMux I__4882 (
            .O(N__21058),
            .I(\receive_module.rx_counter.X_9 ));
    LocalMux I__4881 (
            .O(N__21055),
            .I(\receive_module.rx_counter.X_9 ));
    InMux I__4880 (
            .O(N__21050),
            .I(N__21047));
    LocalMux I__4879 (
            .O(N__21047),
            .I(N__21036));
    ClkMux I__4878 (
            .O(N__21046),
            .I(N__20909));
    ClkMux I__4877 (
            .O(N__21045),
            .I(N__20909));
    ClkMux I__4876 (
            .O(N__21044),
            .I(N__20909));
    ClkMux I__4875 (
            .O(N__21043),
            .I(N__20909));
    ClkMux I__4874 (
            .O(N__21042),
            .I(N__20909));
    ClkMux I__4873 (
            .O(N__21041),
            .I(N__20909));
    ClkMux I__4872 (
            .O(N__21040),
            .I(N__20909));
    ClkMux I__4871 (
            .O(N__21039),
            .I(N__20909));
    Glb2LocalMux I__4870 (
            .O(N__21036),
            .I(N__20909));
    ClkMux I__4869 (
            .O(N__21035),
            .I(N__20909));
    ClkMux I__4868 (
            .O(N__21034),
            .I(N__20909));
    ClkMux I__4867 (
            .O(N__21033),
            .I(N__20909));
    ClkMux I__4866 (
            .O(N__21032),
            .I(N__20909));
    ClkMux I__4865 (
            .O(N__21031),
            .I(N__20909));
    ClkMux I__4864 (
            .O(N__21030),
            .I(N__20909));
    ClkMux I__4863 (
            .O(N__21029),
            .I(N__20909));
    ClkMux I__4862 (
            .O(N__21028),
            .I(N__20909));
    ClkMux I__4861 (
            .O(N__21027),
            .I(N__20909));
    ClkMux I__4860 (
            .O(N__21026),
            .I(N__20909));
    ClkMux I__4859 (
            .O(N__21025),
            .I(N__20909));
    ClkMux I__4858 (
            .O(N__21024),
            .I(N__20909));
    ClkMux I__4857 (
            .O(N__21023),
            .I(N__20909));
    ClkMux I__4856 (
            .O(N__21022),
            .I(N__20909));
    ClkMux I__4855 (
            .O(N__21021),
            .I(N__20909));
    ClkMux I__4854 (
            .O(N__21020),
            .I(N__20909));
    ClkMux I__4853 (
            .O(N__21019),
            .I(N__20909));
    ClkMux I__4852 (
            .O(N__21018),
            .I(N__20909));
    ClkMux I__4851 (
            .O(N__21017),
            .I(N__20909));
    ClkMux I__4850 (
            .O(N__21016),
            .I(N__20909));
    ClkMux I__4849 (
            .O(N__21015),
            .I(N__20909));
    ClkMux I__4848 (
            .O(N__21014),
            .I(N__20909));
    ClkMux I__4847 (
            .O(N__21013),
            .I(N__20909));
    ClkMux I__4846 (
            .O(N__21012),
            .I(N__20909));
    ClkMux I__4845 (
            .O(N__21011),
            .I(N__20909));
    ClkMux I__4844 (
            .O(N__21010),
            .I(N__20909));
    ClkMux I__4843 (
            .O(N__21009),
            .I(N__20909));
    ClkMux I__4842 (
            .O(N__21008),
            .I(N__20909));
    ClkMux I__4841 (
            .O(N__21007),
            .I(N__20909));
    ClkMux I__4840 (
            .O(N__21006),
            .I(N__20909));
    ClkMux I__4839 (
            .O(N__21005),
            .I(N__20909));
    ClkMux I__4838 (
            .O(N__21004),
            .I(N__20909));
    ClkMux I__4837 (
            .O(N__21003),
            .I(N__20909));
    ClkMux I__4836 (
            .O(N__21002),
            .I(N__20909));
    ClkMux I__4835 (
            .O(N__21001),
            .I(N__20909));
    ClkMux I__4834 (
            .O(N__21000),
            .I(N__20909));
    GlobalMux I__4833 (
            .O(N__20909),
            .I(N__20906));
    gio2CtrlBuf I__4832 (
            .O(N__20906),
            .I(TVP_CLK_c));
    SRMux I__4831 (
            .O(N__20903),
            .I(N__20900));
    LocalMux I__4830 (
            .O(N__20900),
            .I(N__20896));
    SRMux I__4829 (
            .O(N__20899),
            .I(N__20893));
    Span4Mux_v I__4828 (
            .O(N__20896),
            .I(N__20890));
    LocalMux I__4827 (
            .O(N__20893),
            .I(N__20887));
    Odrv4 I__4826 (
            .O(N__20890),
            .I(n3860));
    Odrv12 I__4825 (
            .O(N__20887),
            .I(n3860));
    InMux I__4824 (
            .O(N__20882),
            .I(N__20879));
    LocalMux I__4823 (
            .O(N__20879),
            .I(N__20876));
    Odrv12 I__4822 (
            .O(N__20876),
            .I(\line_buffer.n597 ));
    CascadeMux I__4821 (
            .O(N__20873),
            .I(N__20870));
    InMux I__4820 (
            .O(N__20870),
            .I(N__20867));
    LocalMux I__4819 (
            .O(N__20867),
            .I(N__20864));
    Span4Mux_v I__4818 (
            .O(N__20864),
            .I(N__20861));
    Span4Mux_h I__4817 (
            .O(N__20861),
            .I(N__20858));
    Span4Mux_h I__4816 (
            .O(N__20858),
            .I(N__20855));
    Odrv4 I__4815 (
            .O(N__20855),
            .I(\line_buffer.n605 ));
    InMux I__4814 (
            .O(N__20852),
            .I(N__20849));
    LocalMux I__4813 (
            .O(N__20849),
            .I(N__20846));
    Span4Mux_v I__4812 (
            .O(N__20846),
            .I(N__20843));
    Span4Mux_h I__4811 (
            .O(N__20843),
            .I(N__20840));
    Span4Mux_h I__4810 (
            .O(N__20840),
            .I(N__20837));
    Odrv4 I__4809 (
            .O(N__20837),
            .I(\line_buffer.n604 ));
    InMux I__4808 (
            .O(N__20834),
            .I(N__20831));
    LocalMux I__4807 (
            .O(N__20831),
            .I(N__20828));
    Span12Mux_v I__4806 (
            .O(N__20828),
            .I(N__20825));
    Odrv12 I__4805 (
            .O(N__20825),
            .I(\line_buffer.n596 ));
    InMux I__4804 (
            .O(N__20822),
            .I(N__20819));
    LocalMux I__4803 (
            .O(N__20819),
            .I(N__20816));
    Span4Mux_h I__4802 (
            .O(N__20816),
            .I(N__20813));
    Span4Mux_v I__4801 (
            .O(N__20813),
            .I(N__20810));
    Span4Mux_h I__4800 (
            .O(N__20810),
            .I(N__20807));
    Odrv4 I__4799 (
            .O(N__20807),
            .I(\line_buffer.n508 ));
    InMux I__4798 (
            .O(N__20804),
            .I(N__20801));
    LocalMux I__4797 (
            .O(N__20801),
            .I(\line_buffer.n3833 ));
    CascadeMux I__4796 (
            .O(N__20798),
            .I(N__20795));
    InMux I__4795 (
            .O(N__20795),
            .I(N__20792));
    LocalMux I__4794 (
            .O(N__20792),
            .I(N__20789));
    Span4Mux_v I__4793 (
            .O(N__20789),
            .I(N__20786));
    Span4Mux_v I__4792 (
            .O(N__20786),
            .I(N__20783));
    Sp12to4 I__4791 (
            .O(N__20783),
            .I(N__20780));
    Span12Mux_h I__4790 (
            .O(N__20780),
            .I(N__20777));
    Odrv12 I__4789 (
            .O(N__20777),
            .I(\line_buffer.n500 ));
    InMux I__4788 (
            .O(N__20774),
            .I(N__20771));
    LocalMux I__4787 (
            .O(N__20771),
            .I(\line_buffer.n3836 ));
    InMux I__4786 (
            .O(N__20768),
            .I(N__20765));
    LocalMux I__4785 (
            .O(N__20765),
            .I(N__20762));
    Odrv12 I__4784 (
            .O(N__20762),
            .I(\line_buffer.n3721 ));
    InMux I__4783 (
            .O(N__20759),
            .I(N__20756));
    LocalMux I__4782 (
            .O(N__20756),
            .I(N__20753));
    Span4Mux_h I__4781 (
            .O(N__20753),
            .I(N__20750));
    Odrv4 I__4780 (
            .O(N__20750),
            .I(TX_DATA_4));
    InMux I__4779 (
            .O(N__20747),
            .I(N__20743));
    InMux I__4778 (
            .O(N__20746),
            .I(N__20740));
    LocalMux I__4777 (
            .O(N__20743),
            .I(N__20737));
    LocalMux I__4776 (
            .O(N__20740),
            .I(\transmit_module.n179 ));
    Odrv4 I__4775 (
            .O(N__20737),
            .I(\transmit_module.n179 ));
    InMux I__4774 (
            .O(N__20732),
            .I(N__20729));
    LocalMux I__4773 (
            .O(N__20729),
            .I(N__20725));
    InMux I__4772 (
            .O(N__20728),
            .I(N__20722));
    Odrv4 I__4771 (
            .O(N__20725),
            .I(\transmit_module.n211 ));
    LocalMux I__4770 (
            .O(N__20722),
            .I(\transmit_module.n211 ));
    SRMux I__4769 (
            .O(N__20717),
            .I(N__20714));
    LocalMux I__4768 (
            .O(N__20714),
            .I(N__20708));
    SRMux I__4767 (
            .O(N__20713),
            .I(N__20705));
    CascadeMux I__4766 (
            .O(N__20712),
            .I(N__20702));
    SRMux I__4765 (
            .O(N__20711),
            .I(N__20687));
    Span4Mux_v I__4764 (
            .O(N__20708),
            .I(N__20676));
    LocalMux I__4763 (
            .O(N__20705),
            .I(N__20676));
    InMux I__4762 (
            .O(N__20702),
            .I(N__20673));
    CascadeMux I__4761 (
            .O(N__20701),
            .I(N__20670));
    CascadeMux I__4760 (
            .O(N__20700),
            .I(N__20667));
    IoInMux I__4759 (
            .O(N__20699),
            .I(N__20662));
    SRMux I__4758 (
            .O(N__20698),
            .I(N__20657));
    SRMux I__4757 (
            .O(N__20697),
            .I(N__20653));
    SRMux I__4756 (
            .O(N__20696),
            .I(N__20650));
    SRMux I__4755 (
            .O(N__20695),
            .I(N__20646));
    SRMux I__4754 (
            .O(N__20694),
            .I(N__20643));
    SRMux I__4753 (
            .O(N__20693),
            .I(N__20640));
    SRMux I__4752 (
            .O(N__20692),
            .I(N__20637));
    SRMux I__4751 (
            .O(N__20691),
            .I(N__20634));
    SRMux I__4750 (
            .O(N__20690),
            .I(N__20631));
    LocalMux I__4749 (
            .O(N__20687),
            .I(N__20627));
    SRMux I__4748 (
            .O(N__20686),
            .I(N__20624));
    CascadeMux I__4747 (
            .O(N__20685),
            .I(N__20621));
    CascadeMux I__4746 (
            .O(N__20684),
            .I(N__20614));
    SRMux I__4745 (
            .O(N__20683),
            .I(N__20610));
    CascadeMux I__4744 (
            .O(N__20682),
            .I(N__20606));
    CascadeMux I__4743 (
            .O(N__20681),
            .I(N__20602));
    Span4Mux_v I__4742 (
            .O(N__20676),
            .I(N__20593));
    LocalMux I__4741 (
            .O(N__20673),
            .I(N__20593));
    InMux I__4740 (
            .O(N__20670),
            .I(N__20588));
    InMux I__4739 (
            .O(N__20667),
            .I(N__20588));
    CascadeMux I__4738 (
            .O(N__20666),
            .I(N__20584));
    CascadeMux I__4737 (
            .O(N__20665),
            .I(N__20581));
    LocalMux I__4736 (
            .O(N__20662),
            .I(N__20578));
    SRMux I__4735 (
            .O(N__20661),
            .I(N__20574));
    SRMux I__4734 (
            .O(N__20660),
            .I(N__20569));
    LocalMux I__4733 (
            .O(N__20657),
            .I(N__20565));
    SRMux I__4732 (
            .O(N__20656),
            .I(N__20562));
    LocalMux I__4731 (
            .O(N__20653),
            .I(N__20557));
    LocalMux I__4730 (
            .O(N__20650),
            .I(N__20557));
    SRMux I__4729 (
            .O(N__20649),
            .I(N__20554));
    LocalMux I__4728 (
            .O(N__20646),
            .I(N__20545));
    LocalMux I__4727 (
            .O(N__20643),
            .I(N__20545));
    LocalMux I__4726 (
            .O(N__20640),
            .I(N__20545));
    LocalMux I__4725 (
            .O(N__20637),
            .I(N__20545));
    LocalMux I__4724 (
            .O(N__20634),
            .I(N__20540));
    LocalMux I__4723 (
            .O(N__20631),
            .I(N__20540));
    SRMux I__4722 (
            .O(N__20630),
            .I(N__20537));
    Span4Mux_h I__4721 (
            .O(N__20627),
            .I(N__20532));
    LocalMux I__4720 (
            .O(N__20624),
            .I(N__20532));
    InMux I__4719 (
            .O(N__20621),
            .I(N__20525));
    InMux I__4718 (
            .O(N__20620),
            .I(N__20525));
    InMux I__4717 (
            .O(N__20619),
            .I(N__20525));
    SRMux I__4716 (
            .O(N__20618),
            .I(N__20522));
    CascadeMux I__4715 (
            .O(N__20617),
            .I(N__20519));
    InMux I__4714 (
            .O(N__20614),
            .I(N__20513));
    SRMux I__4713 (
            .O(N__20613),
            .I(N__20509));
    LocalMux I__4712 (
            .O(N__20610),
            .I(N__20505));
    SRMux I__4711 (
            .O(N__20609),
            .I(N__20502));
    InMux I__4710 (
            .O(N__20606),
            .I(N__20495));
    InMux I__4709 (
            .O(N__20605),
            .I(N__20495));
    InMux I__4708 (
            .O(N__20602),
            .I(N__20495));
    CascadeMux I__4707 (
            .O(N__20601),
            .I(N__20492));
    CascadeMux I__4706 (
            .O(N__20600),
            .I(N__20486));
    InMux I__4705 (
            .O(N__20599),
            .I(N__20481));
    InMux I__4704 (
            .O(N__20598),
            .I(N__20481));
    Span4Mux_h I__4703 (
            .O(N__20593),
            .I(N__20476));
    LocalMux I__4702 (
            .O(N__20588),
            .I(N__20476));
    InMux I__4701 (
            .O(N__20587),
            .I(N__20471));
    InMux I__4700 (
            .O(N__20584),
            .I(N__20471));
    InMux I__4699 (
            .O(N__20581),
            .I(N__20468));
    Span4Mux_s3_h I__4698 (
            .O(N__20578),
            .I(N__20465));
    SRMux I__4697 (
            .O(N__20577),
            .I(N__20462));
    LocalMux I__4696 (
            .O(N__20574),
            .I(N__20459));
    InMux I__4695 (
            .O(N__20573),
            .I(N__20456));
    CascadeMux I__4694 (
            .O(N__20572),
            .I(N__20453));
    LocalMux I__4693 (
            .O(N__20569),
            .I(N__20449));
    SRMux I__4692 (
            .O(N__20568),
            .I(N__20446));
    Span4Mux_v I__4691 (
            .O(N__20565),
            .I(N__20431));
    LocalMux I__4690 (
            .O(N__20562),
            .I(N__20431));
    Span4Mux_v I__4689 (
            .O(N__20557),
            .I(N__20431));
    LocalMux I__4688 (
            .O(N__20554),
            .I(N__20431));
    Span4Mux_v I__4687 (
            .O(N__20545),
            .I(N__20431));
    Span4Mux_h I__4686 (
            .O(N__20540),
            .I(N__20431));
    LocalMux I__4685 (
            .O(N__20537),
            .I(N__20431));
    Span4Mux_v I__4684 (
            .O(N__20532),
            .I(N__20424));
    LocalMux I__4683 (
            .O(N__20525),
            .I(N__20424));
    LocalMux I__4682 (
            .O(N__20522),
            .I(N__20424));
    InMux I__4681 (
            .O(N__20519),
            .I(N__20421));
    SRMux I__4680 (
            .O(N__20518),
            .I(N__20418));
    SRMux I__4679 (
            .O(N__20517),
            .I(N__20415));
    SRMux I__4678 (
            .O(N__20516),
            .I(N__20412));
    LocalMux I__4677 (
            .O(N__20513),
            .I(N__20409));
    InMux I__4676 (
            .O(N__20512),
            .I(N__20406));
    LocalMux I__4675 (
            .O(N__20509),
            .I(N__20403));
    InMux I__4674 (
            .O(N__20508),
            .I(N__20400));
    Span4Mux_h I__4673 (
            .O(N__20505),
            .I(N__20395));
    LocalMux I__4672 (
            .O(N__20502),
            .I(N__20395));
    LocalMux I__4671 (
            .O(N__20495),
            .I(N__20392));
    InMux I__4670 (
            .O(N__20492),
            .I(N__20385));
    InMux I__4669 (
            .O(N__20491),
            .I(N__20385));
    InMux I__4668 (
            .O(N__20490),
            .I(N__20385));
    InMux I__4667 (
            .O(N__20489),
            .I(N__20378));
    InMux I__4666 (
            .O(N__20486),
            .I(N__20378));
    LocalMux I__4665 (
            .O(N__20481),
            .I(N__20369));
    Span4Mux_h I__4664 (
            .O(N__20476),
            .I(N__20369));
    LocalMux I__4663 (
            .O(N__20471),
            .I(N__20369));
    LocalMux I__4662 (
            .O(N__20468),
            .I(N__20369));
    Sp12to4 I__4661 (
            .O(N__20465),
            .I(N__20363));
    LocalMux I__4660 (
            .O(N__20462),
            .I(N__20360));
    Span4Mux_v I__4659 (
            .O(N__20459),
            .I(N__20357));
    LocalMux I__4658 (
            .O(N__20456),
            .I(N__20354));
    InMux I__4657 (
            .O(N__20453),
            .I(N__20349));
    InMux I__4656 (
            .O(N__20452),
            .I(N__20349));
    Span4Mux_v I__4655 (
            .O(N__20449),
            .I(N__20342));
    LocalMux I__4654 (
            .O(N__20446),
            .I(N__20342));
    Span4Mux_v I__4653 (
            .O(N__20431),
            .I(N__20342));
    Span4Mux_v I__4652 (
            .O(N__20424),
            .I(N__20337));
    LocalMux I__4651 (
            .O(N__20421),
            .I(N__20337));
    LocalMux I__4650 (
            .O(N__20418),
            .I(N__20328));
    LocalMux I__4649 (
            .O(N__20415),
            .I(N__20328));
    LocalMux I__4648 (
            .O(N__20412),
            .I(N__20328));
    Span4Mux_v I__4647 (
            .O(N__20409),
            .I(N__20328));
    LocalMux I__4646 (
            .O(N__20406),
            .I(N__20315));
    Span4Mux_v I__4645 (
            .O(N__20403),
            .I(N__20315));
    LocalMux I__4644 (
            .O(N__20400),
            .I(N__20315));
    Span4Mux_h I__4643 (
            .O(N__20395),
            .I(N__20315));
    Span4Mux_h I__4642 (
            .O(N__20392),
            .I(N__20315));
    LocalMux I__4641 (
            .O(N__20385),
            .I(N__20315));
    InMux I__4640 (
            .O(N__20384),
            .I(N__20310));
    InMux I__4639 (
            .O(N__20383),
            .I(N__20310));
    LocalMux I__4638 (
            .O(N__20378),
            .I(N__20305));
    Span4Mux_v I__4637 (
            .O(N__20369),
            .I(N__20305));
    SRMux I__4636 (
            .O(N__20368),
            .I(N__20302));
    SRMux I__4635 (
            .O(N__20367),
            .I(N__20299));
    SRMux I__4634 (
            .O(N__20366),
            .I(N__20296));
    Span12Mux_v I__4633 (
            .O(N__20363),
            .I(N__20291));
    Span12Mux_v I__4632 (
            .O(N__20360),
            .I(N__20291));
    Span4Mux_h I__4631 (
            .O(N__20357),
            .I(N__20284));
    Span4Mux_v I__4630 (
            .O(N__20354),
            .I(N__20284));
    LocalMux I__4629 (
            .O(N__20349),
            .I(N__20284));
    Span4Mux_h I__4628 (
            .O(N__20342),
            .I(N__20277));
    Span4Mux_v I__4627 (
            .O(N__20337),
            .I(N__20277));
    Span4Mux_v I__4626 (
            .O(N__20328),
            .I(N__20277));
    Span4Mux_v I__4625 (
            .O(N__20315),
            .I(N__20270));
    LocalMux I__4624 (
            .O(N__20310),
            .I(N__20270));
    Span4Mux_h I__4623 (
            .O(N__20305),
            .I(N__20270));
    LocalMux I__4622 (
            .O(N__20302),
            .I(ADV_VSYNC_c));
    LocalMux I__4621 (
            .O(N__20299),
            .I(ADV_VSYNC_c));
    LocalMux I__4620 (
            .O(N__20296),
            .I(ADV_VSYNC_c));
    Odrv12 I__4619 (
            .O(N__20291),
            .I(ADV_VSYNC_c));
    Odrv4 I__4618 (
            .O(N__20284),
            .I(ADV_VSYNC_c));
    Odrv4 I__4617 (
            .O(N__20277),
            .I(ADV_VSYNC_c));
    Odrv4 I__4616 (
            .O(N__20270),
            .I(ADV_VSYNC_c));
    InMux I__4615 (
            .O(N__20255),
            .I(N__20246));
    InMux I__4614 (
            .O(N__20254),
            .I(N__20241));
    InMux I__4613 (
            .O(N__20253),
            .I(N__20241));
    InMux I__4612 (
            .O(N__20252),
            .I(N__20229));
    InMux I__4611 (
            .O(N__20251),
            .I(N__20222));
    InMux I__4610 (
            .O(N__20250),
            .I(N__20222));
    InMux I__4609 (
            .O(N__20249),
            .I(N__20222));
    LocalMux I__4608 (
            .O(N__20246),
            .I(N__20217));
    LocalMux I__4607 (
            .O(N__20241),
            .I(N__20217));
    InMux I__4606 (
            .O(N__20240),
            .I(N__20212));
    InMux I__4605 (
            .O(N__20239),
            .I(N__20212));
    InMux I__4604 (
            .O(N__20238),
            .I(N__20207));
    InMux I__4603 (
            .O(N__20237),
            .I(N__20207));
    InMux I__4602 (
            .O(N__20236),
            .I(N__20197));
    InMux I__4601 (
            .O(N__20235),
            .I(N__20197));
    InMux I__4600 (
            .O(N__20234),
            .I(N__20197));
    InMux I__4599 (
            .O(N__20233),
            .I(N__20197));
    InMux I__4598 (
            .O(N__20232),
            .I(N__20190));
    LocalMux I__4597 (
            .O(N__20229),
            .I(N__20187));
    LocalMux I__4596 (
            .O(N__20222),
            .I(N__20180));
    Span4Mux_h I__4595 (
            .O(N__20217),
            .I(N__20180));
    LocalMux I__4594 (
            .O(N__20212),
            .I(N__20180));
    LocalMux I__4593 (
            .O(N__20207),
            .I(N__20175));
    InMux I__4592 (
            .O(N__20206),
            .I(N__20172));
    LocalMux I__4591 (
            .O(N__20197),
            .I(N__20169));
    InMux I__4590 (
            .O(N__20196),
            .I(N__20160));
    InMux I__4589 (
            .O(N__20195),
            .I(N__20160));
    InMux I__4588 (
            .O(N__20194),
            .I(N__20160));
    InMux I__4587 (
            .O(N__20193),
            .I(N__20160));
    LocalMux I__4586 (
            .O(N__20190),
            .I(N__20157));
    Span4Mux_v I__4585 (
            .O(N__20187),
            .I(N__20152));
    Span4Mux_v I__4584 (
            .O(N__20180),
            .I(N__20152));
    InMux I__4583 (
            .O(N__20179),
            .I(N__20147));
    InMux I__4582 (
            .O(N__20178),
            .I(N__20147));
    Span4Mux_h I__4581 (
            .O(N__20175),
            .I(N__20136));
    LocalMux I__4580 (
            .O(N__20172),
            .I(N__20136));
    Span4Mux_v I__4579 (
            .O(N__20169),
            .I(N__20136));
    LocalMux I__4578 (
            .O(N__20160),
            .I(N__20136));
    Span4Mux_h I__4577 (
            .O(N__20157),
            .I(N__20136));
    Odrv4 I__4576 (
            .O(N__20152),
            .I(\transmit_module.n3853 ));
    LocalMux I__4575 (
            .O(N__20147),
            .I(\transmit_module.n3853 ));
    Odrv4 I__4574 (
            .O(N__20136),
            .I(\transmit_module.n3853 ));
    CascadeMux I__4573 (
            .O(N__20129),
            .I(N__20125));
    CascadeMux I__4572 (
            .O(N__20128),
            .I(N__20122));
    CascadeBuf I__4571 (
            .O(N__20125),
            .I(N__20119));
    CascadeBuf I__4570 (
            .O(N__20122),
            .I(N__20116));
    CascadeMux I__4569 (
            .O(N__20119),
            .I(N__20113));
    CascadeMux I__4568 (
            .O(N__20116),
            .I(N__20110));
    CascadeBuf I__4567 (
            .O(N__20113),
            .I(N__20107));
    CascadeBuf I__4566 (
            .O(N__20110),
            .I(N__20104));
    CascadeMux I__4565 (
            .O(N__20107),
            .I(N__20101));
    CascadeMux I__4564 (
            .O(N__20104),
            .I(N__20098));
    CascadeBuf I__4563 (
            .O(N__20101),
            .I(N__20095));
    CascadeBuf I__4562 (
            .O(N__20098),
            .I(N__20092));
    CascadeMux I__4561 (
            .O(N__20095),
            .I(N__20089));
    CascadeMux I__4560 (
            .O(N__20092),
            .I(N__20086));
    CascadeBuf I__4559 (
            .O(N__20089),
            .I(N__20083));
    CascadeBuf I__4558 (
            .O(N__20086),
            .I(N__20080));
    CascadeMux I__4557 (
            .O(N__20083),
            .I(N__20077));
    CascadeMux I__4556 (
            .O(N__20080),
            .I(N__20074));
    CascadeBuf I__4555 (
            .O(N__20077),
            .I(N__20071));
    CascadeBuf I__4554 (
            .O(N__20074),
            .I(N__20068));
    CascadeMux I__4553 (
            .O(N__20071),
            .I(N__20065));
    CascadeMux I__4552 (
            .O(N__20068),
            .I(N__20062));
    CascadeBuf I__4551 (
            .O(N__20065),
            .I(N__20059));
    CascadeBuf I__4550 (
            .O(N__20062),
            .I(N__20056));
    CascadeMux I__4549 (
            .O(N__20059),
            .I(N__20053));
    CascadeMux I__4548 (
            .O(N__20056),
            .I(N__20050));
    CascadeBuf I__4547 (
            .O(N__20053),
            .I(N__20047));
    CascadeBuf I__4546 (
            .O(N__20050),
            .I(N__20044));
    CascadeMux I__4545 (
            .O(N__20047),
            .I(N__20041));
    CascadeMux I__4544 (
            .O(N__20044),
            .I(N__20038));
    CascadeBuf I__4543 (
            .O(N__20041),
            .I(N__20035));
    CascadeBuf I__4542 (
            .O(N__20038),
            .I(N__20032));
    CascadeMux I__4541 (
            .O(N__20035),
            .I(N__20029));
    CascadeMux I__4540 (
            .O(N__20032),
            .I(N__20026));
    CascadeBuf I__4539 (
            .O(N__20029),
            .I(N__20023));
    CascadeBuf I__4538 (
            .O(N__20026),
            .I(N__20020));
    CascadeMux I__4537 (
            .O(N__20023),
            .I(N__20017));
    CascadeMux I__4536 (
            .O(N__20020),
            .I(N__20014));
    CascadeBuf I__4535 (
            .O(N__20017),
            .I(N__20011));
    CascadeBuf I__4534 (
            .O(N__20014),
            .I(N__20008));
    CascadeMux I__4533 (
            .O(N__20011),
            .I(N__20005));
    CascadeMux I__4532 (
            .O(N__20008),
            .I(N__20002));
    CascadeBuf I__4531 (
            .O(N__20005),
            .I(N__19999));
    CascadeBuf I__4530 (
            .O(N__20002),
            .I(N__19996));
    CascadeMux I__4529 (
            .O(N__19999),
            .I(N__19993));
    CascadeMux I__4528 (
            .O(N__19996),
            .I(N__19990));
    CascadeBuf I__4527 (
            .O(N__19993),
            .I(N__19987));
    CascadeBuf I__4526 (
            .O(N__19990),
            .I(N__19984));
    CascadeMux I__4525 (
            .O(N__19987),
            .I(N__19981));
    CascadeMux I__4524 (
            .O(N__19984),
            .I(N__19978));
    CascadeBuf I__4523 (
            .O(N__19981),
            .I(N__19975));
    CascadeBuf I__4522 (
            .O(N__19978),
            .I(N__19972));
    CascadeMux I__4521 (
            .O(N__19975),
            .I(N__19969));
    CascadeMux I__4520 (
            .O(N__19972),
            .I(N__19966));
    CascadeBuf I__4519 (
            .O(N__19969),
            .I(N__19963));
    CascadeBuf I__4518 (
            .O(N__19966),
            .I(N__19960));
    CascadeMux I__4517 (
            .O(N__19963),
            .I(N__19957));
    CascadeMux I__4516 (
            .O(N__19960),
            .I(N__19954));
    CascadeBuf I__4515 (
            .O(N__19957),
            .I(N__19951));
    CascadeBuf I__4514 (
            .O(N__19954),
            .I(N__19948));
    CascadeMux I__4513 (
            .O(N__19951),
            .I(N__19945));
    CascadeMux I__4512 (
            .O(N__19948),
            .I(N__19942));
    InMux I__4511 (
            .O(N__19945),
            .I(N__19939));
    InMux I__4510 (
            .O(N__19942),
            .I(N__19936));
    LocalMux I__4509 (
            .O(N__19939),
            .I(N__19933));
    LocalMux I__4508 (
            .O(N__19936),
            .I(N__19930));
    Span12Mux_h I__4507 (
            .O(N__19933),
            .I(N__19927));
    Span12Mux_s11_h I__4506 (
            .O(N__19930),
            .I(N__19924));
    Span12Mux_v I__4505 (
            .O(N__19927),
            .I(N__19921));
    Span12Mux_v I__4504 (
            .O(N__19924),
            .I(N__19918));
    Odrv12 I__4503 (
            .O(N__19921),
            .I(n19));
    Odrv12 I__4502 (
            .O(N__19918),
            .I(n19));
    InMux I__4501 (
            .O(N__19913),
            .I(N__19907));
    InMux I__4500 (
            .O(N__19912),
            .I(N__19907));
    LocalMux I__4499 (
            .O(N__19907),
            .I(N__19903));
    InMux I__4498 (
            .O(N__19906),
            .I(N__19900));
    Span4Mux_v I__4497 (
            .O(N__19903),
            .I(N__19897));
    LocalMux I__4496 (
            .O(N__19900),
            .I(N__19894));
    Span4Mux_h I__4495 (
            .O(N__19897),
            .I(N__19891));
    Span4Mux_h I__4494 (
            .O(N__19894),
            .I(N__19888));
    Span4Mux_h I__4493 (
            .O(N__19891),
            .I(N__19883));
    Span4Mux_v I__4492 (
            .O(N__19888),
            .I(N__19883));
    Odrv4 I__4491 (
            .O(N__19883),
            .I(TVP_HSYNC_c));
    InMux I__4490 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__4489 (
            .O(N__19877),
            .I(\receive_module.rx_counter.n10 ));
    InMux I__4488 (
            .O(N__19874),
            .I(bfn_17_9_0_));
    InMux I__4487 (
            .O(N__19871),
            .I(N__19868));
    LocalMux I__4486 (
            .O(N__19868),
            .I(\receive_module.rx_counter.n9 ));
    InMux I__4485 (
            .O(N__19865),
            .I(\receive_module.rx_counter.n3357 ));
    InMux I__4484 (
            .O(N__19862),
            .I(N__19859));
    LocalMux I__4483 (
            .O(N__19859),
            .I(\receive_module.rx_counter.n8 ));
    InMux I__4482 (
            .O(N__19856),
            .I(\receive_module.rx_counter.n3358 ));
    InMux I__4481 (
            .O(N__19853),
            .I(N__19849));
    InMux I__4480 (
            .O(N__19852),
            .I(N__19846));
    LocalMux I__4479 (
            .O(N__19849),
            .I(\receive_module.rx_counter.X_3 ));
    LocalMux I__4478 (
            .O(N__19846),
            .I(\receive_module.rx_counter.X_3 ));
    InMux I__4477 (
            .O(N__19841),
            .I(\receive_module.rx_counter.n3359 ));
    InMux I__4476 (
            .O(N__19838),
            .I(N__19834));
    InMux I__4475 (
            .O(N__19837),
            .I(N__19831));
    LocalMux I__4474 (
            .O(N__19834),
            .I(\receive_module.rx_counter.X_4 ));
    LocalMux I__4473 (
            .O(N__19831),
            .I(\receive_module.rx_counter.X_4 ));
    InMux I__4472 (
            .O(N__19826),
            .I(\receive_module.rx_counter.n3360 ));
    InMux I__4471 (
            .O(N__19823),
            .I(N__19819));
    InMux I__4470 (
            .O(N__19822),
            .I(N__19816));
    LocalMux I__4469 (
            .O(N__19819),
            .I(\receive_module.rx_counter.X_5 ));
    LocalMux I__4468 (
            .O(N__19816),
            .I(\receive_module.rx_counter.X_5 ));
    InMux I__4467 (
            .O(N__19811),
            .I(\receive_module.rx_counter.n3361 ));
    InMux I__4466 (
            .O(N__19808),
            .I(N__19803));
    InMux I__4465 (
            .O(N__19807),
            .I(N__19798));
    InMux I__4464 (
            .O(N__19806),
            .I(N__19798));
    LocalMux I__4463 (
            .O(N__19803),
            .I(\receive_module.rx_counter.X_6 ));
    LocalMux I__4462 (
            .O(N__19798),
            .I(\receive_module.rx_counter.X_6 ));
    InMux I__4461 (
            .O(N__19793),
            .I(\receive_module.rx_counter.n3362 ));
    CascadeMux I__4460 (
            .O(N__19790),
            .I(\transmit_module.n210_cascade_ ));
    CascadeMux I__4459 (
            .O(N__19787),
            .I(N__19784));
    InMux I__4458 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__4457 (
            .O(N__19781),
            .I(N__19778));
    Odrv4 I__4456 (
            .O(N__19778),
            .I(\transmit_module.n201 ));
    CascadeMux I__4455 (
            .O(N__19775),
            .I(\transmit_module.n217_cascade_ ));
    InMux I__4454 (
            .O(N__19772),
            .I(N__19769));
    LocalMux I__4453 (
            .O(N__19769),
            .I(N__19765));
    InMux I__4452 (
            .O(N__19768),
            .I(N__19760));
    Span4Mux_h I__4451 (
            .O(N__19765),
            .I(N__19757));
    InMux I__4450 (
            .O(N__19764),
            .I(N__19754));
    InMux I__4449 (
            .O(N__19763),
            .I(N__19751));
    LocalMux I__4448 (
            .O(N__19760),
            .I(N__19748));
    Odrv4 I__4447 (
            .O(N__19757),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__4446 (
            .O(N__19754),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__4445 (
            .O(N__19751),
            .I(\transmit_module.TX_ADDR_3 ));
    Odrv4 I__4444 (
            .O(N__19748),
            .I(\transmit_module.TX_ADDR_3 ));
    CascadeMux I__4443 (
            .O(N__19739),
            .I(N__19734));
    CascadeMux I__4442 (
            .O(N__19738),
            .I(N__19731));
    CascadeMux I__4441 (
            .O(N__19737),
            .I(N__19724));
    InMux I__4440 (
            .O(N__19734),
            .I(N__19716));
    InMux I__4439 (
            .O(N__19731),
            .I(N__19716));
    InMux I__4438 (
            .O(N__19730),
            .I(N__19709));
    InMux I__4437 (
            .O(N__19729),
            .I(N__19709));
    InMux I__4436 (
            .O(N__19728),
            .I(N__19709));
    CascadeMux I__4435 (
            .O(N__19727),
            .I(N__19704));
    InMux I__4434 (
            .O(N__19724),
            .I(N__19701));
    InMux I__4433 (
            .O(N__19723),
            .I(N__19698));
    InMux I__4432 (
            .O(N__19722),
            .I(N__19693));
    InMux I__4431 (
            .O(N__19721),
            .I(N__19693));
    LocalMux I__4430 (
            .O(N__19716),
            .I(N__19688));
    LocalMux I__4429 (
            .O(N__19709),
            .I(N__19688));
    InMux I__4428 (
            .O(N__19708),
            .I(N__19685));
    InMux I__4427 (
            .O(N__19707),
            .I(N__19682));
    InMux I__4426 (
            .O(N__19704),
            .I(N__19679));
    LocalMux I__4425 (
            .O(N__19701),
            .I(N__19674));
    LocalMux I__4424 (
            .O(N__19698),
            .I(N__19674));
    LocalMux I__4423 (
            .O(N__19693),
            .I(N__19669));
    Span4Mux_h I__4422 (
            .O(N__19688),
            .I(N__19669));
    LocalMux I__4421 (
            .O(N__19685),
            .I(\transmit_module.n3855 ));
    LocalMux I__4420 (
            .O(N__19682),
            .I(\transmit_module.n3855 ));
    LocalMux I__4419 (
            .O(N__19679),
            .I(\transmit_module.n3855 ));
    Odrv4 I__4418 (
            .O(N__19674),
            .I(\transmit_module.n3855 ));
    Odrv4 I__4417 (
            .O(N__19669),
            .I(\transmit_module.n3855 ));
    InMux I__4416 (
            .O(N__19658),
            .I(N__19655));
    LocalMux I__4415 (
            .O(N__19655),
            .I(N__19652));
    Span4Mux_v I__4414 (
            .O(N__19652),
            .I(N__19649));
    Odrv4 I__4413 (
            .O(N__19649),
            .I(\transmit_module.n195 ));
    CascadeMux I__4412 (
            .O(N__19646),
            .I(N__19643));
    InMux I__4411 (
            .O(N__19643),
            .I(N__19640));
    LocalMux I__4410 (
            .O(N__19640),
            .I(N__19637));
    Span4Mux_h I__4409 (
            .O(N__19637),
            .I(N__19631));
    InMux I__4408 (
            .O(N__19636),
            .I(N__19628));
    InMux I__4407 (
            .O(N__19635),
            .I(N__19623));
    InMux I__4406 (
            .O(N__19634),
            .I(N__19623));
    Odrv4 I__4405 (
            .O(N__19631),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__4404 (
            .O(N__19628),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__4403 (
            .O(N__19623),
            .I(\transmit_module.TX_ADDR_9 ));
    InMux I__4402 (
            .O(N__19616),
            .I(N__19610));
    InMux I__4401 (
            .O(N__19615),
            .I(N__19610));
    LocalMux I__4400 (
            .O(N__19610),
            .I(N__19602));
    InMux I__4399 (
            .O(N__19609),
            .I(N__19597));
    InMux I__4398 (
            .O(N__19608),
            .I(N__19597));
    InMux I__4397 (
            .O(N__19607),
            .I(N__19594));
    InMux I__4396 (
            .O(N__19606),
            .I(N__19586));
    InMux I__4395 (
            .O(N__19605),
            .I(N__19583));
    Span4Mux_v I__4394 (
            .O(N__19602),
            .I(N__19576));
    LocalMux I__4393 (
            .O(N__19597),
            .I(N__19576));
    LocalMux I__4392 (
            .O(N__19594),
            .I(N__19576));
    InMux I__4391 (
            .O(N__19593),
            .I(N__19569));
    InMux I__4390 (
            .O(N__19592),
            .I(N__19569));
    InMux I__4389 (
            .O(N__19591),
            .I(N__19569));
    InMux I__4388 (
            .O(N__19590),
            .I(N__19564));
    InMux I__4387 (
            .O(N__19589),
            .I(N__19561));
    LocalMux I__4386 (
            .O(N__19586),
            .I(N__19558));
    LocalMux I__4385 (
            .O(N__19583),
            .I(N__19555));
    Span4Mux_h I__4384 (
            .O(N__19576),
            .I(N__19550));
    LocalMux I__4383 (
            .O(N__19569),
            .I(N__19550));
    InMux I__4382 (
            .O(N__19568),
            .I(N__19537));
    InMux I__4381 (
            .O(N__19567),
            .I(N__19537));
    LocalMux I__4380 (
            .O(N__19564),
            .I(N__19530));
    LocalMux I__4379 (
            .O(N__19561),
            .I(N__19530));
    Span4Mux_h I__4378 (
            .O(N__19558),
            .I(N__19530));
    Span4Mux_v I__4377 (
            .O(N__19555),
            .I(N__19525));
    Span4Mux_v I__4376 (
            .O(N__19550),
            .I(N__19525));
    InMux I__4375 (
            .O(N__19549),
            .I(N__19516));
    InMux I__4374 (
            .O(N__19548),
            .I(N__19516));
    InMux I__4373 (
            .O(N__19547),
            .I(N__19516));
    InMux I__4372 (
            .O(N__19546),
            .I(N__19516));
    InMux I__4371 (
            .O(N__19545),
            .I(N__19507));
    InMux I__4370 (
            .O(N__19544),
            .I(N__19507));
    InMux I__4369 (
            .O(N__19543),
            .I(N__19507));
    InMux I__4368 (
            .O(N__19542),
            .I(N__19507));
    LocalMux I__4367 (
            .O(N__19537),
            .I(\transmit_module.n3549 ));
    Odrv4 I__4366 (
            .O(N__19530),
            .I(\transmit_module.n3549 ));
    Odrv4 I__4365 (
            .O(N__19525),
            .I(\transmit_module.n3549 ));
    LocalMux I__4364 (
            .O(N__19516),
            .I(\transmit_module.n3549 ));
    LocalMux I__4363 (
            .O(N__19507),
            .I(\transmit_module.n3549 ));
    InMux I__4362 (
            .O(N__19496),
            .I(N__19493));
    LocalMux I__4361 (
            .O(N__19493),
            .I(\transmit_module.n217 ));
    InMux I__4360 (
            .O(N__19490),
            .I(N__19486));
    InMux I__4359 (
            .O(N__19489),
            .I(N__19483));
    LocalMux I__4358 (
            .O(N__19486),
            .I(\transmit_module.n185 ));
    LocalMux I__4357 (
            .O(N__19483),
            .I(\transmit_module.n185 ));
    CascadeMux I__4356 (
            .O(N__19478),
            .I(N__19474));
    CascadeMux I__4355 (
            .O(N__19477),
            .I(N__19471));
    CascadeBuf I__4354 (
            .O(N__19474),
            .I(N__19468));
    CascadeBuf I__4353 (
            .O(N__19471),
            .I(N__19465));
    CascadeMux I__4352 (
            .O(N__19468),
            .I(N__19462));
    CascadeMux I__4351 (
            .O(N__19465),
            .I(N__19459));
    CascadeBuf I__4350 (
            .O(N__19462),
            .I(N__19456));
    CascadeBuf I__4349 (
            .O(N__19459),
            .I(N__19453));
    CascadeMux I__4348 (
            .O(N__19456),
            .I(N__19450));
    CascadeMux I__4347 (
            .O(N__19453),
            .I(N__19447));
    CascadeBuf I__4346 (
            .O(N__19450),
            .I(N__19444));
    CascadeBuf I__4345 (
            .O(N__19447),
            .I(N__19441));
    CascadeMux I__4344 (
            .O(N__19444),
            .I(N__19438));
    CascadeMux I__4343 (
            .O(N__19441),
            .I(N__19435));
    CascadeBuf I__4342 (
            .O(N__19438),
            .I(N__19432));
    CascadeBuf I__4341 (
            .O(N__19435),
            .I(N__19429));
    CascadeMux I__4340 (
            .O(N__19432),
            .I(N__19426));
    CascadeMux I__4339 (
            .O(N__19429),
            .I(N__19423));
    CascadeBuf I__4338 (
            .O(N__19426),
            .I(N__19420));
    CascadeBuf I__4337 (
            .O(N__19423),
            .I(N__19417));
    CascadeMux I__4336 (
            .O(N__19420),
            .I(N__19414));
    CascadeMux I__4335 (
            .O(N__19417),
            .I(N__19411));
    CascadeBuf I__4334 (
            .O(N__19414),
            .I(N__19408));
    CascadeBuf I__4333 (
            .O(N__19411),
            .I(N__19405));
    CascadeMux I__4332 (
            .O(N__19408),
            .I(N__19402));
    CascadeMux I__4331 (
            .O(N__19405),
            .I(N__19399));
    CascadeBuf I__4330 (
            .O(N__19402),
            .I(N__19396));
    CascadeBuf I__4329 (
            .O(N__19399),
            .I(N__19393));
    CascadeMux I__4328 (
            .O(N__19396),
            .I(N__19390));
    CascadeMux I__4327 (
            .O(N__19393),
            .I(N__19387));
    CascadeBuf I__4326 (
            .O(N__19390),
            .I(N__19384));
    CascadeBuf I__4325 (
            .O(N__19387),
            .I(N__19381));
    CascadeMux I__4324 (
            .O(N__19384),
            .I(N__19378));
    CascadeMux I__4323 (
            .O(N__19381),
            .I(N__19375));
    CascadeBuf I__4322 (
            .O(N__19378),
            .I(N__19372));
    CascadeBuf I__4321 (
            .O(N__19375),
            .I(N__19369));
    CascadeMux I__4320 (
            .O(N__19372),
            .I(N__19366));
    CascadeMux I__4319 (
            .O(N__19369),
            .I(N__19363));
    CascadeBuf I__4318 (
            .O(N__19366),
            .I(N__19360));
    CascadeBuf I__4317 (
            .O(N__19363),
            .I(N__19357));
    CascadeMux I__4316 (
            .O(N__19360),
            .I(N__19354));
    CascadeMux I__4315 (
            .O(N__19357),
            .I(N__19351));
    CascadeBuf I__4314 (
            .O(N__19354),
            .I(N__19348));
    CascadeBuf I__4313 (
            .O(N__19351),
            .I(N__19345));
    CascadeMux I__4312 (
            .O(N__19348),
            .I(N__19342));
    CascadeMux I__4311 (
            .O(N__19345),
            .I(N__19339));
    CascadeBuf I__4310 (
            .O(N__19342),
            .I(N__19336));
    CascadeBuf I__4309 (
            .O(N__19339),
            .I(N__19333));
    CascadeMux I__4308 (
            .O(N__19336),
            .I(N__19330));
    CascadeMux I__4307 (
            .O(N__19333),
            .I(N__19327));
    CascadeBuf I__4306 (
            .O(N__19330),
            .I(N__19324));
    CascadeBuf I__4305 (
            .O(N__19327),
            .I(N__19321));
    CascadeMux I__4304 (
            .O(N__19324),
            .I(N__19318));
    CascadeMux I__4303 (
            .O(N__19321),
            .I(N__19315));
    CascadeBuf I__4302 (
            .O(N__19318),
            .I(N__19312));
    CascadeBuf I__4301 (
            .O(N__19315),
            .I(N__19309));
    CascadeMux I__4300 (
            .O(N__19312),
            .I(N__19306));
    CascadeMux I__4299 (
            .O(N__19309),
            .I(N__19303));
    CascadeBuf I__4298 (
            .O(N__19306),
            .I(N__19300));
    CascadeBuf I__4297 (
            .O(N__19303),
            .I(N__19297));
    CascadeMux I__4296 (
            .O(N__19300),
            .I(N__19294));
    CascadeMux I__4295 (
            .O(N__19297),
            .I(N__19291));
    InMux I__4294 (
            .O(N__19294),
            .I(N__19288));
    InMux I__4293 (
            .O(N__19291),
            .I(N__19285));
    LocalMux I__4292 (
            .O(N__19288),
            .I(N__19282));
    LocalMux I__4291 (
            .O(N__19285),
            .I(N__19279));
    Span4Mux_h I__4290 (
            .O(N__19282),
            .I(N__19276));
    Span4Mux_h I__4289 (
            .O(N__19279),
            .I(N__19273));
    Sp12to4 I__4288 (
            .O(N__19276),
            .I(N__19270));
    Sp12to4 I__4287 (
            .O(N__19273),
            .I(N__19267));
    Span12Mux_v I__4286 (
            .O(N__19270),
            .I(N__19262));
    Span12Mux_v I__4285 (
            .O(N__19267),
            .I(N__19262));
    Odrv12 I__4284 (
            .O(N__19262),
            .I(n25));
    InMux I__4283 (
            .O(N__19259),
            .I(N__19254));
    InMux I__4282 (
            .O(N__19258),
            .I(N__19246));
    InMux I__4281 (
            .O(N__19257),
            .I(N__19242));
    LocalMux I__4280 (
            .O(N__19254),
            .I(N__19239));
    InMux I__4279 (
            .O(N__19253),
            .I(N__19236));
    InMux I__4278 (
            .O(N__19252),
            .I(N__19233));
    InMux I__4277 (
            .O(N__19251),
            .I(N__19228));
    InMux I__4276 (
            .O(N__19250),
            .I(N__19228));
    InMux I__4275 (
            .O(N__19249),
            .I(N__19223));
    LocalMux I__4274 (
            .O(N__19246),
            .I(N__19218));
    InMux I__4273 (
            .O(N__19245),
            .I(N__19215));
    LocalMux I__4272 (
            .O(N__19242),
            .I(N__19212));
    Span4Mux_h I__4271 (
            .O(N__19239),
            .I(N__19207));
    LocalMux I__4270 (
            .O(N__19236),
            .I(N__19207));
    LocalMux I__4269 (
            .O(N__19233),
            .I(N__19202));
    LocalMux I__4268 (
            .O(N__19228),
            .I(N__19202));
    InMux I__4267 (
            .O(N__19227),
            .I(N__19197));
    InMux I__4266 (
            .O(N__19226),
            .I(N__19197));
    LocalMux I__4265 (
            .O(N__19223),
            .I(N__19194));
    InMux I__4264 (
            .O(N__19222),
            .I(N__19189));
    InMux I__4263 (
            .O(N__19221),
            .I(N__19189));
    Sp12to4 I__4262 (
            .O(N__19218),
            .I(N__19183));
    LocalMux I__4261 (
            .O(N__19215),
            .I(N__19183));
    Span4Mux_v I__4260 (
            .O(N__19212),
            .I(N__19180));
    Span4Mux_h I__4259 (
            .O(N__19207),
            .I(N__19177));
    Span4Mux_v I__4258 (
            .O(N__19202),
            .I(N__19172));
    LocalMux I__4257 (
            .O(N__19197),
            .I(N__19172));
    Span4Mux_h I__4256 (
            .O(N__19194),
            .I(N__19167));
    LocalMux I__4255 (
            .O(N__19189),
            .I(N__19167));
    InMux I__4254 (
            .O(N__19188),
            .I(N__19164));
    Span12Mux_v I__4253 (
            .O(N__19183),
            .I(N__19161));
    Span4Mux_v I__4252 (
            .O(N__19180),
            .I(N__19158));
    Span4Mux_v I__4251 (
            .O(N__19177),
            .I(N__19155));
    Span4Mux_v I__4250 (
            .O(N__19172),
            .I(N__19150));
    Span4Mux_v I__4249 (
            .O(N__19167),
            .I(N__19150));
    LocalMux I__4248 (
            .O(N__19164),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv12 I__4247 (
            .O(N__19161),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4246 (
            .O(N__19158),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4245 (
            .O(N__19155),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4244 (
            .O(N__19150),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    InMux I__4243 (
            .O(N__19139),
            .I(N__19136));
    LocalMux I__4242 (
            .O(N__19136),
            .I(\transmit_module.ADDR_Y_COMPONENT_10 ));
    InMux I__4241 (
            .O(N__19133),
            .I(N__19129));
    CascadeMux I__4240 (
            .O(N__19132),
            .I(N__19124));
    LocalMux I__4239 (
            .O(N__19129),
            .I(N__19121));
    InMux I__4238 (
            .O(N__19128),
            .I(N__19118));
    InMux I__4237 (
            .O(N__19127),
            .I(N__19115));
    InMux I__4236 (
            .O(N__19124),
            .I(N__19112));
    Span4Mux_v I__4235 (
            .O(N__19121),
            .I(N__19109));
    LocalMux I__4234 (
            .O(N__19118),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__4233 (
            .O(N__19115),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__4232 (
            .O(N__19112),
            .I(\transmit_module.TX_ADDR_10 ));
    Odrv4 I__4231 (
            .O(N__19109),
            .I(\transmit_module.TX_ADDR_10 ));
    InMux I__4230 (
            .O(N__19100),
            .I(N__19097));
    LocalMux I__4229 (
            .O(N__19097),
            .I(\transmit_module.n178 ));
    InMux I__4228 (
            .O(N__19094),
            .I(N__19091));
    LocalMux I__4227 (
            .O(N__19091),
            .I(\transmit_module.n210 ));
    CascadeMux I__4226 (
            .O(N__19088),
            .I(\transmit_module.n178_cascade_ ));
    CascadeMux I__4225 (
            .O(N__19085),
            .I(N__19082));
    CascadeBuf I__4224 (
            .O(N__19082),
            .I(N__19078));
    CascadeMux I__4223 (
            .O(N__19081),
            .I(N__19075));
    CascadeMux I__4222 (
            .O(N__19078),
            .I(N__19072));
    CascadeBuf I__4221 (
            .O(N__19075),
            .I(N__19069));
    CascadeBuf I__4220 (
            .O(N__19072),
            .I(N__19066));
    CascadeMux I__4219 (
            .O(N__19069),
            .I(N__19063));
    CascadeMux I__4218 (
            .O(N__19066),
            .I(N__19060));
    CascadeBuf I__4217 (
            .O(N__19063),
            .I(N__19057));
    CascadeBuf I__4216 (
            .O(N__19060),
            .I(N__19054));
    CascadeMux I__4215 (
            .O(N__19057),
            .I(N__19051));
    CascadeMux I__4214 (
            .O(N__19054),
            .I(N__19048));
    CascadeBuf I__4213 (
            .O(N__19051),
            .I(N__19045));
    CascadeBuf I__4212 (
            .O(N__19048),
            .I(N__19042));
    CascadeMux I__4211 (
            .O(N__19045),
            .I(N__19039));
    CascadeMux I__4210 (
            .O(N__19042),
            .I(N__19036));
    CascadeBuf I__4209 (
            .O(N__19039),
            .I(N__19033));
    CascadeBuf I__4208 (
            .O(N__19036),
            .I(N__19030));
    CascadeMux I__4207 (
            .O(N__19033),
            .I(N__19027));
    CascadeMux I__4206 (
            .O(N__19030),
            .I(N__19024));
    CascadeBuf I__4205 (
            .O(N__19027),
            .I(N__19021));
    CascadeBuf I__4204 (
            .O(N__19024),
            .I(N__19018));
    CascadeMux I__4203 (
            .O(N__19021),
            .I(N__19015));
    CascadeMux I__4202 (
            .O(N__19018),
            .I(N__19012));
    CascadeBuf I__4201 (
            .O(N__19015),
            .I(N__19009));
    CascadeBuf I__4200 (
            .O(N__19012),
            .I(N__19006));
    CascadeMux I__4199 (
            .O(N__19009),
            .I(N__19003));
    CascadeMux I__4198 (
            .O(N__19006),
            .I(N__19000));
    CascadeBuf I__4197 (
            .O(N__19003),
            .I(N__18997));
    CascadeBuf I__4196 (
            .O(N__19000),
            .I(N__18994));
    CascadeMux I__4195 (
            .O(N__18997),
            .I(N__18991));
    CascadeMux I__4194 (
            .O(N__18994),
            .I(N__18988));
    CascadeBuf I__4193 (
            .O(N__18991),
            .I(N__18985));
    CascadeBuf I__4192 (
            .O(N__18988),
            .I(N__18982));
    CascadeMux I__4191 (
            .O(N__18985),
            .I(N__18979));
    CascadeMux I__4190 (
            .O(N__18982),
            .I(N__18976));
    CascadeBuf I__4189 (
            .O(N__18979),
            .I(N__18973));
    CascadeBuf I__4188 (
            .O(N__18976),
            .I(N__18970));
    CascadeMux I__4187 (
            .O(N__18973),
            .I(N__18967));
    CascadeMux I__4186 (
            .O(N__18970),
            .I(N__18964));
    CascadeBuf I__4185 (
            .O(N__18967),
            .I(N__18961));
    CascadeBuf I__4184 (
            .O(N__18964),
            .I(N__18958));
    CascadeMux I__4183 (
            .O(N__18961),
            .I(N__18955));
    CascadeMux I__4182 (
            .O(N__18958),
            .I(N__18952));
    CascadeBuf I__4181 (
            .O(N__18955),
            .I(N__18949));
    CascadeBuf I__4180 (
            .O(N__18952),
            .I(N__18946));
    CascadeMux I__4179 (
            .O(N__18949),
            .I(N__18943));
    CascadeMux I__4178 (
            .O(N__18946),
            .I(N__18940));
    CascadeBuf I__4177 (
            .O(N__18943),
            .I(N__18937));
    CascadeBuf I__4176 (
            .O(N__18940),
            .I(N__18934));
    CascadeMux I__4175 (
            .O(N__18937),
            .I(N__18931));
    CascadeMux I__4174 (
            .O(N__18934),
            .I(N__18928));
    CascadeBuf I__4173 (
            .O(N__18931),
            .I(N__18925));
    CascadeBuf I__4172 (
            .O(N__18928),
            .I(N__18922));
    CascadeMux I__4171 (
            .O(N__18925),
            .I(N__18919));
    CascadeMux I__4170 (
            .O(N__18922),
            .I(N__18916));
    CascadeBuf I__4169 (
            .O(N__18919),
            .I(N__18913));
    CascadeBuf I__4168 (
            .O(N__18916),
            .I(N__18910));
    CascadeMux I__4167 (
            .O(N__18913),
            .I(N__18907));
    CascadeMux I__4166 (
            .O(N__18910),
            .I(N__18904));
    CascadeBuf I__4165 (
            .O(N__18907),
            .I(N__18901));
    InMux I__4164 (
            .O(N__18904),
            .I(N__18898));
    CascadeMux I__4163 (
            .O(N__18901),
            .I(N__18895));
    LocalMux I__4162 (
            .O(N__18898),
            .I(N__18892));
    InMux I__4161 (
            .O(N__18895),
            .I(N__18889));
    Span12Mux_h I__4160 (
            .O(N__18892),
            .I(N__18886));
    LocalMux I__4159 (
            .O(N__18889),
            .I(N__18883));
    Span12Mux_v I__4158 (
            .O(N__18886),
            .I(N__18878));
    Span12Mux_v I__4157 (
            .O(N__18883),
            .I(N__18878));
    Odrv12 I__4156 (
            .O(N__18878),
            .I(n18));
    IoInMux I__4155 (
            .O(N__18875),
            .I(N__18872));
    LocalMux I__4154 (
            .O(N__18872),
            .I(N__18869));
    Span4Mux_s0_v I__4153 (
            .O(N__18869),
            .I(N__18866));
    Odrv4 I__4152 (
            .O(N__18866),
            .I(GB_BUFFER_TVP_CLK_c_THRU_CO));
    CascadeMux I__4151 (
            .O(N__18863),
            .I(\receive_module.rx_counter.n3547_cascade_ ));
    InMux I__4150 (
            .O(N__18860),
            .I(N__18857));
    LocalMux I__4149 (
            .O(N__18857),
            .I(\receive_module.rx_counter.n3547 ));
    CascadeMux I__4148 (
            .O(N__18854),
            .I(\receive_module.rx_counter.n3646_cascade_ ));
    InMux I__4147 (
            .O(N__18851),
            .I(N__18848));
    LocalMux I__4146 (
            .O(N__18848),
            .I(\receive_module.rx_counter.n3613 ));
    InMux I__4145 (
            .O(N__18845),
            .I(N__18842));
    LocalMux I__4144 (
            .O(N__18842),
            .I(N__18839));
    Odrv4 I__4143 (
            .O(N__18839),
            .I(\receive_module.rx_counter.n28 ));
    InMux I__4142 (
            .O(N__18836),
            .I(N__18833));
    LocalMux I__4141 (
            .O(N__18833),
            .I(N__18830));
    Span4Mux_h I__4140 (
            .O(N__18830),
            .I(N__18827));
    Sp12to4 I__4139 (
            .O(N__18827),
            .I(N__18824));
    Span12Mux_v I__4138 (
            .O(N__18824),
            .I(N__18821));
    Odrv12 I__4137 (
            .O(N__18821),
            .I(\line_buffer.n629 ));
    CascadeMux I__4136 (
            .O(N__18818),
            .I(N__18815));
    InMux I__4135 (
            .O(N__18815),
            .I(N__18812));
    LocalMux I__4134 (
            .O(N__18812),
            .I(N__18809));
    Odrv12 I__4133 (
            .O(N__18809),
            .I(\line_buffer.n637 ));
    InMux I__4132 (
            .O(N__18806),
            .I(N__18803));
    LocalMux I__4131 (
            .O(N__18803),
            .I(N__18800));
    Span4Mux_v I__4130 (
            .O(N__18800),
            .I(N__18797));
    Span4Mux_h I__4129 (
            .O(N__18797),
            .I(N__18794));
    Span4Mux_h I__4128 (
            .O(N__18794),
            .I(N__18791));
    Odrv4 I__4127 (
            .O(N__18791),
            .I(\line_buffer.n565 ));
    CascadeMux I__4126 (
            .O(N__18788),
            .I(\line_buffer.n3761_cascade_ ));
    InMux I__4125 (
            .O(N__18785),
            .I(N__18782));
    LocalMux I__4124 (
            .O(N__18782),
            .I(N__18779));
    Span4Mux_h I__4123 (
            .O(N__18779),
            .I(N__18776));
    Sp12to4 I__4122 (
            .O(N__18776),
            .I(N__18773));
    Span12Mux_v I__4121 (
            .O(N__18773),
            .I(N__18770));
    Odrv12 I__4120 (
            .O(N__18770),
            .I(\line_buffer.n573 ));
    InMux I__4119 (
            .O(N__18767),
            .I(N__18764));
    LocalMux I__4118 (
            .O(N__18764),
            .I(\line_buffer.n3764 ));
    InMux I__4117 (
            .O(N__18761),
            .I(N__18758));
    LocalMux I__4116 (
            .O(N__18758),
            .I(N__18755));
    Span4Mux_h I__4115 (
            .O(N__18755),
            .I(N__18752));
    Odrv4 I__4114 (
            .O(N__18752),
            .I(TX_DATA_5));
    InMux I__4113 (
            .O(N__18749),
            .I(N__18746));
    LocalMux I__4112 (
            .O(N__18746),
            .I(\transmit_module.Y_DELTA_PATTERN_33 ));
    InMux I__4111 (
            .O(N__18743),
            .I(N__18740));
    LocalMux I__4110 (
            .O(N__18740),
            .I(N__18737));
    Span12Mux_v I__4109 (
            .O(N__18737),
            .I(N__18734));
    Odrv12 I__4108 (
            .O(N__18734),
            .I(\transmit_module.Y_DELTA_PATTERN_32 ));
    CEMux I__4107 (
            .O(N__18731),
            .I(N__18727));
    CEMux I__4106 (
            .O(N__18730),
            .I(N__18721));
    LocalMux I__4105 (
            .O(N__18727),
            .I(N__18717));
    CEMux I__4104 (
            .O(N__18726),
            .I(N__18714));
    CEMux I__4103 (
            .O(N__18725),
            .I(N__18709));
    SRMux I__4102 (
            .O(N__18724),
            .I(N__18704));
    LocalMux I__4101 (
            .O(N__18721),
            .I(N__18698));
    CEMux I__4100 (
            .O(N__18720),
            .I(N__18695));
    Span4Mux_h I__4099 (
            .O(N__18717),
            .I(N__18688));
    LocalMux I__4098 (
            .O(N__18714),
            .I(N__18688));
    CEMux I__4097 (
            .O(N__18713),
            .I(N__18685));
    CEMux I__4096 (
            .O(N__18712),
            .I(N__18682));
    LocalMux I__4095 (
            .O(N__18709),
            .I(N__18679));
    CEMux I__4094 (
            .O(N__18708),
            .I(N__18676));
    CEMux I__4093 (
            .O(N__18707),
            .I(N__18673));
    LocalMux I__4092 (
            .O(N__18704),
            .I(N__18670));
    SRMux I__4091 (
            .O(N__18703),
            .I(N__18667));
    SRMux I__4090 (
            .O(N__18702),
            .I(N__18664));
    SRMux I__4089 (
            .O(N__18701),
            .I(N__18661));
    Span4Mux_h I__4088 (
            .O(N__18698),
            .I(N__18656));
    LocalMux I__4087 (
            .O(N__18695),
            .I(N__18656));
    SRMux I__4086 (
            .O(N__18694),
            .I(N__18653));
    SRMux I__4085 (
            .O(N__18693),
            .I(N__18650));
    Span4Mux_v I__4084 (
            .O(N__18688),
            .I(N__18647));
    LocalMux I__4083 (
            .O(N__18685),
            .I(N__18644));
    LocalMux I__4082 (
            .O(N__18682),
            .I(N__18641));
    Span4Mux_h I__4081 (
            .O(N__18679),
            .I(N__18638));
    LocalMux I__4080 (
            .O(N__18676),
            .I(N__18635));
    LocalMux I__4079 (
            .O(N__18673),
            .I(N__18632));
    Span4Mux_h I__4078 (
            .O(N__18670),
            .I(N__18627));
    LocalMux I__4077 (
            .O(N__18667),
            .I(N__18627));
    LocalMux I__4076 (
            .O(N__18664),
            .I(N__18624));
    LocalMux I__4075 (
            .O(N__18661),
            .I(N__18621));
    Span4Mux_v I__4074 (
            .O(N__18656),
            .I(N__18618));
    LocalMux I__4073 (
            .O(N__18653),
            .I(N__18613));
    LocalMux I__4072 (
            .O(N__18650),
            .I(N__18613));
    Span4Mux_h I__4071 (
            .O(N__18647),
            .I(N__18610));
    Span4Mux_h I__4070 (
            .O(N__18644),
            .I(N__18603));
    Span4Mux_v I__4069 (
            .O(N__18641),
            .I(N__18603));
    Span4Mux_h I__4068 (
            .O(N__18638),
            .I(N__18603));
    Span4Mux_h I__4067 (
            .O(N__18635),
            .I(N__18598));
    Span4Mux_v I__4066 (
            .O(N__18632),
            .I(N__18598));
    Span4Mux_v I__4065 (
            .O(N__18627),
            .I(N__18595));
    Span4Mux_v I__4064 (
            .O(N__18624),
            .I(N__18592));
    Span12Mux_s11_h I__4063 (
            .O(N__18621),
            .I(N__18589));
    Span4Mux_h I__4062 (
            .O(N__18618),
            .I(N__18584));
    Span4Mux_v I__4061 (
            .O(N__18613),
            .I(N__18584));
    Odrv4 I__4060 (
            .O(N__18610),
            .I(\transmit_module.n3864 ));
    Odrv4 I__4059 (
            .O(N__18603),
            .I(\transmit_module.n3864 ));
    Odrv4 I__4058 (
            .O(N__18598),
            .I(\transmit_module.n3864 ));
    Odrv4 I__4057 (
            .O(N__18595),
            .I(\transmit_module.n3864 ));
    Odrv4 I__4056 (
            .O(N__18592),
            .I(\transmit_module.n3864 ));
    Odrv12 I__4055 (
            .O(N__18589),
            .I(\transmit_module.n3864 ));
    Odrv4 I__4054 (
            .O(N__18584),
            .I(\transmit_module.n3864 ));
    InMux I__4053 (
            .O(N__18569),
            .I(N__18566));
    LocalMux I__4052 (
            .O(N__18566),
            .I(N__18563));
    Span4Mux_h I__4051 (
            .O(N__18563),
            .I(N__18560));
    Span4Mux_v I__4050 (
            .O(N__18560),
            .I(N__18557));
    Span4Mux_h I__4049 (
            .O(N__18557),
            .I(N__18554));
    Odrv4 I__4048 (
            .O(N__18554),
            .I(\line_buffer.n607 ));
    InMux I__4047 (
            .O(N__18551),
            .I(N__18548));
    LocalMux I__4046 (
            .O(N__18548),
            .I(N__18545));
    Span4Mux_v I__4045 (
            .O(N__18545),
            .I(N__18542));
    Sp12to4 I__4044 (
            .O(N__18542),
            .I(N__18539));
    Span12Mux_v I__4043 (
            .O(N__18539),
            .I(N__18536));
    Odrv12 I__4042 (
            .O(N__18536),
            .I(\line_buffer.n599 ));
    InMux I__4041 (
            .O(N__18533),
            .I(N__18530));
    LocalMux I__4040 (
            .O(N__18530),
            .I(\line_buffer.n3718 ));
    InMux I__4039 (
            .O(N__18527),
            .I(N__18524));
    LocalMux I__4038 (
            .O(N__18524),
            .I(N__18521));
    Span4Mux_h I__4037 (
            .O(N__18521),
            .I(N__18518));
    Odrv4 I__4036 (
            .O(N__18518),
            .I(\transmit_module.n194 ));
    InMux I__4035 (
            .O(N__18515),
            .I(N__18512));
    LocalMux I__4034 (
            .O(N__18512),
            .I(N__18509));
    Span4Mux_v I__4033 (
            .O(N__18509),
            .I(N__18506));
    Span4Mux_h I__4032 (
            .O(N__18506),
            .I(N__18503));
    Odrv4 I__4031 (
            .O(N__18503),
            .I(\line_buffer.n575 ));
    InMux I__4030 (
            .O(N__18500),
            .I(N__18497));
    LocalMux I__4029 (
            .O(N__18497),
            .I(N__18494));
    Span4Mux_v I__4028 (
            .O(N__18494),
            .I(N__18491));
    Sp12to4 I__4027 (
            .O(N__18491),
            .I(N__18488));
    Span12Mux_h I__4026 (
            .O(N__18488),
            .I(N__18485));
    Span12Mux_v I__4025 (
            .O(N__18485),
            .I(N__18482));
    Odrv12 I__4024 (
            .O(N__18482),
            .I(\line_buffer.n567 ));
    InMux I__4023 (
            .O(N__18479),
            .I(N__18476));
    LocalMux I__4022 (
            .O(N__18476),
            .I(\line_buffer.n3702 ));
    InMux I__4021 (
            .O(N__18473),
            .I(N__18470));
    LocalMux I__4020 (
            .O(N__18470),
            .I(\transmit_module.ADDR_Y_COMPONENT_3 ));
    CEMux I__4019 (
            .O(N__18467),
            .I(N__18463));
    CEMux I__4018 (
            .O(N__18466),
            .I(N__18460));
    LocalMux I__4017 (
            .O(N__18463),
            .I(N__18455));
    LocalMux I__4016 (
            .O(N__18460),
            .I(N__18452));
    CEMux I__4015 (
            .O(N__18459),
            .I(N__18449));
    CEMux I__4014 (
            .O(N__18458),
            .I(N__18446));
    Span4Mux_v I__4013 (
            .O(N__18455),
            .I(N__18443));
    Sp12to4 I__4012 (
            .O(N__18452),
            .I(N__18438));
    LocalMux I__4011 (
            .O(N__18449),
            .I(N__18438));
    LocalMux I__4010 (
            .O(N__18446),
            .I(N__18435));
    Odrv4 I__4009 (
            .O(N__18443),
            .I(\transmit_module.n2321 ));
    Odrv12 I__4008 (
            .O(N__18438),
            .I(\transmit_module.n2321 ));
    Odrv4 I__4007 (
            .O(N__18435),
            .I(\transmit_module.n2321 ));
    InMux I__4006 (
            .O(N__18428),
            .I(N__18425));
    LocalMux I__4005 (
            .O(N__18425),
            .I(N__18422));
    Span4Mux_v I__4004 (
            .O(N__18422),
            .I(N__18419));
    Span4Mux_v I__4003 (
            .O(N__18419),
            .I(N__18416));
    Span4Mux_v I__4002 (
            .O(N__18416),
            .I(N__18413));
    Sp12to4 I__4001 (
            .O(N__18413),
            .I(N__18410));
    Odrv12 I__4000 (
            .O(N__18410),
            .I(\line_buffer.n625 ));
    CascadeMux I__3999 (
            .O(N__18407),
            .I(N__18404));
    InMux I__3998 (
            .O(N__18404),
            .I(N__18401));
    LocalMux I__3997 (
            .O(N__18401),
            .I(N__18398));
    Span4Mux_v I__3996 (
            .O(N__18398),
            .I(N__18395));
    Span4Mux_h I__3995 (
            .O(N__18395),
            .I(N__18392));
    Odrv4 I__3994 (
            .O(N__18392),
            .I(\line_buffer.n633 ));
    InMux I__3993 (
            .O(N__18389),
            .I(N__18386));
    LocalMux I__3992 (
            .O(N__18386),
            .I(N__18383));
    Span4Mux_v I__3991 (
            .O(N__18383),
            .I(N__18380));
    Odrv4 I__3990 (
            .O(N__18380),
            .I(\line_buffer.n3827 ));
    InMux I__3989 (
            .O(N__18377),
            .I(N__18374));
    LocalMux I__3988 (
            .O(N__18374),
            .I(N__18371));
    Span4Mux_v I__3987 (
            .O(N__18371),
            .I(N__18368));
    Sp12to4 I__3986 (
            .O(N__18368),
            .I(N__18365));
    Span12Mux_h I__3985 (
            .O(N__18365),
            .I(N__18362));
    Span12Mux_v I__3984 (
            .O(N__18362),
            .I(N__18359));
    Odrv12 I__3983 (
            .O(N__18359),
            .I(\line_buffer.n598 ));
    CascadeMux I__3982 (
            .O(N__18356),
            .I(N__18353));
    InMux I__3981 (
            .O(N__18353),
            .I(N__18350));
    LocalMux I__3980 (
            .O(N__18350),
            .I(N__18347));
    Span4Mux_v I__3979 (
            .O(N__18347),
            .I(N__18344));
    Span4Mux_h I__3978 (
            .O(N__18344),
            .I(N__18341));
    Odrv4 I__3977 (
            .O(N__18341),
            .I(\line_buffer.n606 ));
    InMux I__3976 (
            .O(N__18338),
            .I(N__18335));
    LocalMux I__3975 (
            .O(N__18335),
            .I(\line_buffer.n3767 ));
    InMux I__3974 (
            .O(N__18332),
            .I(N__18329));
    LocalMux I__3973 (
            .O(N__18329),
            .I(N__18326));
    Span4Mux_v I__3972 (
            .O(N__18326),
            .I(N__18323));
    Sp12to4 I__3971 (
            .O(N__18323),
            .I(N__18320));
    Odrv12 I__3970 (
            .O(N__18320),
            .I(\line_buffer.n506 ));
    InMux I__3969 (
            .O(N__18317),
            .I(N__18314));
    LocalMux I__3968 (
            .O(N__18314),
            .I(N__18311));
    Span4Mux_v I__3967 (
            .O(N__18311),
            .I(N__18308));
    Sp12to4 I__3966 (
            .O(N__18308),
            .I(N__18305));
    Span12Mux_h I__3965 (
            .O(N__18305),
            .I(N__18302));
    Odrv12 I__3964 (
            .O(N__18302),
            .I(\line_buffer.n498 ));
    InMux I__3963 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__3962 (
            .O(N__18296),
            .I(N__18293));
    Span4Mux_v I__3961 (
            .O(N__18293),
            .I(N__18290));
    Odrv4 I__3960 (
            .O(N__18290),
            .I(\line_buffer.n3714 ));
    InMux I__3959 (
            .O(N__18287),
            .I(N__18284));
    LocalMux I__3958 (
            .O(N__18284),
            .I(N__18281));
    Span12Mux_h I__3957 (
            .O(N__18281),
            .I(N__18278));
    Odrv12 I__3956 (
            .O(N__18278),
            .I(\line_buffer.n510 ));
    InMux I__3955 (
            .O(N__18275),
            .I(N__18272));
    LocalMux I__3954 (
            .O(N__18272),
            .I(N__18269));
    Span4Mux_h I__3953 (
            .O(N__18269),
            .I(N__18266));
    Span4Mux_h I__3952 (
            .O(N__18266),
            .I(N__18263));
    Odrv4 I__3951 (
            .O(N__18263),
            .I(\line_buffer.n502 ));
    InMux I__3950 (
            .O(N__18260),
            .I(N__18257));
    LocalMux I__3949 (
            .O(N__18257),
            .I(N__18254));
    Span4Mux_v I__3948 (
            .O(N__18254),
            .I(N__18251));
    Odrv4 I__3947 (
            .O(N__18251),
            .I(\line_buffer.n3717 ));
    InMux I__3946 (
            .O(N__18248),
            .I(N__18245));
    LocalMux I__3945 (
            .O(N__18245),
            .I(N__18242));
    Odrv4 I__3944 (
            .O(N__18242),
            .I(\line_buffer.n3715 ));
    CascadeMux I__3943 (
            .O(N__18239),
            .I(\line_buffer.n3773_cascade_ ));
    InMux I__3942 (
            .O(N__18236),
            .I(N__18233));
    LocalMux I__3941 (
            .O(N__18233),
            .I(N__18230));
    Odrv4 I__3940 (
            .O(N__18230),
            .I(TX_DATA_3));
    InMux I__3939 (
            .O(N__18227),
            .I(N__18224));
    LocalMux I__3938 (
            .O(N__18224),
            .I(N__18221));
    Span12Mux_h I__3937 (
            .O(N__18221),
            .I(N__18218));
    Odrv12 I__3936 (
            .O(N__18218),
            .I(\line_buffer.n594 ));
    CascadeMux I__3935 (
            .O(N__18215),
            .I(N__18212));
    InMux I__3934 (
            .O(N__18212),
            .I(N__18209));
    LocalMux I__3933 (
            .O(N__18209),
            .I(N__18206));
    Span4Mux_v I__3932 (
            .O(N__18206),
            .I(N__18203));
    Span4Mux_h I__3931 (
            .O(N__18203),
            .I(N__18200));
    Span4Mux_h I__3930 (
            .O(N__18200),
            .I(N__18197));
    Odrv4 I__3929 (
            .O(N__18197),
            .I(\line_buffer.n602 ));
    InMux I__3928 (
            .O(N__18194),
            .I(N__18191));
    LocalMux I__3927 (
            .O(N__18191),
            .I(N__18188));
    Span4Mux_h I__3926 (
            .O(N__18188),
            .I(N__18185));
    Span4Mux_v I__3925 (
            .O(N__18185),
            .I(N__18182));
    Sp12to4 I__3924 (
            .O(N__18182),
            .I(N__18179));
    Span12Mux_v I__3923 (
            .O(N__18179),
            .I(N__18176));
    Odrv12 I__3922 (
            .O(N__18176),
            .I(\line_buffer.n497 ));
    CascadeMux I__3921 (
            .O(N__18173),
            .I(\line_buffer.n3803_cascade_ ));
    InMux I__3920 (
            .O(N__18170),
            .I(N__18167));
    LocalMux I__3919 (
            .O(N__18167),
            .I(N__18164));
    Span4Mux_v I__3918 (
            .O(N__18164),
            .I(N__18161));
    Span4Mux_v I__3917 (
            .O(N__18161),
            .I(N__18158));
    Sp12to4 I__3916 (
            .O(N__18158),
            .I(N__18155));
    Odrv12 I__3915 (
            .O(N__18155),
            .I(\line_buffer.n505 ));
    CascadeMux I__3914 (
            .O(N__18152),
            .I(\line_buffer.n3806_cascade_ ));
    InMux I__3913 (
            .O(N__18149),
            .I(N__18146));
    LocalMux I__3912 (
            .O(N__18146),
            .I(\line_buffer.n3782 ));
    InMux I__3911 (
            .O(N__18143),
            .I(N__18140));
    LocalMux I__3910 (
            .O(N__18140),
            .I(N__18137));
    Odrv12 I__3909 (
            .O(N__18137),
            .I(TX_DATA_2));
    InMux I__3908 (
            .O(N__18134),
            .I(N__18131));
    LocalMux I__3907 (
            .O(N__18131),
            .I(N__18128));
    Odrv12 I__3906 (
            .O(N__18128),
            .I(\line_buffer.n635 ));
    InMux I__3905 (
            .O(N__18125),
            .I(N__18122));
    LocalMux I__3904 (
            .O(N__18122),
            .I(N__18119));
    Span12Mux_h I__3903 (
            .O(N__18119),
            .I(N__18116));
    Span12Mux_v I__3902 (
            .O(N__18116),
            .I(N__18113));
    Odrv12 I__3901 (
            .O(N__18113),
            .I(\line_buffer.n627 ));
    InMux I__3900 (
            .O(N__18110),
            .I(N__18107));
    LocalMux I__3899 (
            .O(N__18107),
            .I(\line_buffer.n3706 ));
    InMux I__3898 (
            .O(N__18104),
            .I(N__18101));
    LocalMux I__3897 (
            .O(N__18101),
            .I(N__18098));
    Span4Mux_v I__3896 (
            .O(N__18098),
            .I(N__18095));
    Sp12to4 I__3895 (
            .O(N__18095),
            .I(N__18092));
    Span12Mux_h I__3894 (
            .O(N__18092),
            .I(N__18089));
    Span12Mux_v I__3893 (
            .O(N__18089),
            .I(N__18086));
    Odrv12 I__3892 (
            .O(N__18086),
            .I(\line_buffer.n626 ));
    CascadeMux I__3891 (
            .O(N__18083),
            .I(N__18080));
    InMux I__3890 (
            .O(N__18080),
            .I(N__18077));
    LocalMux I__3889 (
            .O(N__18077),
            .I(N__18074));
    Span4Mux_h I__3888 (
            .O(N__18074),
            .I(N__18071));
    Span4Mux_h I__3887 (
            .O(N__18071),
            .I(N__18068));
    Odrv4 I__3886 (
            .O(N__18068),
            .I(\line_buffer.n634 ));
    InMux I__3885 (
            .O(N__18065),
            .I(N__18062));
    LocalMux I__3884 (
            .O(N__18062),
            .I(\line_buffer.n3779 ));
    InMux I__3883 (
            .O(N__18059),
            .I(N__18056));
    LocalMux I__3882 (
            .O(N__18056),
            .I(N__18053));
    Odrv12 I__3881 (
            .O(N__18053),
            .I(\line_buffer.n3703 ));
    CascadeMux I__3880 (
            .O(N__18050),
            .I(\line_buffer.n3791_cascade_ ));
    InMux I__3879 (
            .O(N__18047),
            .I(N__18044));
    LocalMux I__3878 (
            .O(N__18044),
            .I(N__18041));
    Span4Mux_h I__3877 (
            .O(N__18041),
            .I(N__18038));
    Odrv4 I__3876 (
            .O(N__18038),
            .I(TX_DATA_7));
    InMux I__3875 (
            .O(N__18035),
            .I(N__18032));
    LocalMux I__3874 (
            .O(N__18032),
            .I(\transmit_module.Y_DELTA_PATTERN_38 ));
    InMux I__3873 (
            .O(N__18029),
            .I(N__18026));
    LocalMux I__3872 (
            .O(N__18026),
            .I(\transmit_module.Y_DELTA_PATTERN_35 ));
    InMux I__3871 (
            .O(N__18023),
            .I(N__18020));
    LocalMux I__3870 (
            .O(N__18020),
            .I(\transmit_module.Y_DELTA_PATTERN_37 ));
    InMux I__3869 (
            .O(N__18017),
            .I(N__18014));
    LocalMux I__3868 (
            .O(N__18014),
            .I(\transmit_module.Y_DELTA_PATTERN_36 ));
    InMux I__3867 (
            .O(N__18011),
            .I(N__18008));
    LocalMux I__3866 (
            .O(N__18008),
            .I(N__18005));
    Span4Mux_h I__3865 (
            .O(N__18005),
            .I(N__18002));
    Span4Mux_h I__3864 (
            .O(N__18002),
            .I(N__17999));
    Odrv4 I__3863 (
            .O(N__17999),
            .I(\transmit_module.Y_DELTA_PATTERN_40 ));
    InMux I__3862 (
            .O(N__17996),
            .I(N__17993));
    LocalMux I__3861 (
            .O(N__17993),
            .I(\transmit_module.Y_DELTA_PATTERN_39 ));
    InMux I__3860 (
            .O(N__17990),
            .I(N__17987));
    LocalMux I__3859 (
            .O(N__17987),
            .I(\transmit_module.Y_DELTA_PATTERN_34 ));
    CEMux I__3858 (
            .O(N__17984),
            .I(N__17977));
    CEMux I__3857 (
            .O(N__17983),
            .I(N__17974));
    CEMux I__3856 (
            .O(N__17982),
            .I(N__17971));
    CEMux I__3855 (
            .O(N__17981),
            .I(N__17966));
    CEMux I__3854 (
            .O(N__17980),
            .I(N__17963));
    LocalMux I__3853 (
            .O(N__17977),
            .I(N__17959));
    LocalMux I__3852 (
            .O(N__17974),
            .I(N__17954));
    LocalMux I__3851 (
            .O(N__17971),
            .I(N__17954));
    CEMux I__3850 (
            .O(N__17970),
            .I(N__17951));
    CEMux I__3849 (
            .O(N__17969),
            .I(N__17948));
    LocalMux I__3848 (
            .O(N__17966),
            .I(N__17943));
    LocalMux I__3847 (
            .O(N__17963),
            .I(N__17943));
    CEMux I__3846 (
            .O(N__17962),
            .I(N__17940));
    Span4Mux_v I__3845 (
            .O(N__17959),
            .I(N__17936));
    Span4Mux_v I__3844 (
            .O(N__17954),
            .I(N__17931));
    LocalMux I__3843 (
            .O(N__17951),
            .I(N__17931));
    LocalMux I__3842 (
            .O(N__17948),
            .I(N__17928));
    Span4Mux_v I__3841 (
            .O(N__17943),
            .I(N__17925));
    LocalMux I__3840 (
            .O(N__17940),
            .I(N__17922));
    CEMux I__3839 (
            .O(N__17939),
            .I(N__17919));
    Span4Mux_h I__3838 (
            .O(N__17936),
            .I(N__17914));
    Span4Mux_h I__3837 (
            .O(N__17931),
            .I(N__17914));
    Span4Mux_h I__3836 (
            .O(N__17928),
            .I(N__17910));
    Span4Mux_h I__3835 (
            .O(N__17925),
            .I(N__17905));
    Span4Mux_v I__3834 (
            .O(N__17922),
            .I(N__17905));
    LocalMux I__3833 (
            .O(N__17919),
            .I(N__17902));
    Span4Mux_h I__3832 (
            .O(N__17914),
            .I(N__17899));
    CEMux I__3831 (
            .O(N__17913),
            .I(N__17896));
    Odrv4 I__3830 (
            .O(N__17910),
            .I(\transmit_module.n3865 ));
    Odrv4 I__3829 (
            .O(N__17905),
            .I(\transmit_module.n3865 ));
    Odrv12 I__3828 (
            .O(N__17902),
            .I(\transmit_module.n3865 ));
    Odrv4 I__3827 (
            .O(N__17899),
            .I(\transmit_module.n3865 ));
    LocalMux I__3826 (
            .O(N__17896),
            .I(\transmit_module.n3865 ));
    InMux I__3825 (
            .O(N__17885),
            .I(N__17882));
    LocalMux I__3824 (
            .O(N__17882),
            .I(N__17879));
    Span12Mux_h I__3823 (
            .O(N__17879),
            .I(N__17876));
    Span12Mux_v I__3822 (
            .O(N__17876),
            .I(N__17873));
    Odrv12 I__3821 (
            .O(N__17873),
            .I(\line_buffer.n570 ));
    CascadeMux I__3820 (
            .O(N__17870),
            .I(N__17867));
    InMux I__3819 (
            .O(N__17867),
            .I(N__17864));
    LocalMux I__3818 (
            .O(N__17864),
            .I(N__17861));
    Span4Mux_v I__3817 (
            .O(N__17861),
            .I(N__17858));
    Span4Mux_v I__3816 (
            .O(N__17858),
            .I(N__17855));
    Sp12to4 I__3815 (
            .O(N__17855),
            .I(N__17852));
    Odrv12 I__3814 (
            .O(N__17852),
            .I(\line_buffer.n562 ));
    InMux I__3813 (
            .O(N__17849),
            .I(N__17846));
    LocalMux I__3812 (
            .O(N__17846),
            .I(N__17843));
    Odrv12 I__3811 (
            .O(N__17843),
            .I(\line_buffer.n3705 ));
    CascadeMux I__3810 (
            .O(N__17840),
            .I(N__17829));
    CascadeMux I__3809 (
            .O(N__17839),
            .I(N__17826));
    CascadeMux I__3808 (
            .O(N__17838),
            .I(N__17823));
    CascadeMux I__3807 (
            .O(N__17837),
            .I(N__17820));
    CascadeMux I__3806 (
            .O(N__17836),
            .I(N__17817));
    CascadeMux I__3805 (
            .O(N__17835),
            .I(N__17814));
    CascadeMux I__3804 (
            .O(N__17834),
            .I(N__17808));
    CascadeMux I__3803 (
            .O(N__17833),
            .I(N__17805));
    CascadeMux I__3802 (
            .O(N__17832),
            .I(N__17802));
    InMux I__3801 (
            .O(N__17829),
            .I(N__17792));
    InMux I__3800 (
            .O(N__17826),
            .I(N__17792));
    InMux I__3799 (
            .O(N__17823),
            .I(N__17792));
    InMux I__3798 (
            .O(N__17820),
            .I(N__17792));
    InMux I__3797 (
            .O(N__17817),
            .I(N__17785));
    InMux I__3796 (
            .O(N__17814),
            .I(N__17785));
    InMux I__3795 (
            .O(N__17813),
            .I(N__17785));
    InMux I__3794 (
            .O(N__17812),
            .I(N__17774));
    InMux I__3793 (
            .O(N__17811),
            .I(N__17774));
    InMux I__3792 (
            .O(N__17808),
            .I(N__17774));
    InMux I__3791 (
            .O(N__17805),
            .I(N__17774));
    InMux I__3790 (
            .O(N__17802),
            .I(N__17774));
    InMux I__3789 (
            .O(N__17801),
            .I(N__17767));
    LocalMux I__3788 (
            .O(N__17792),
            .I(N__17762));
    LocalMux I__3787 (
            .O(N__17785),
            .I(N__17762));
    LocalMux I__3786 (
            .O(N__17774),
            .I(N__17759));
    InMux I__3785 (
            .O(N__17773),
            .I(N__17753));
    InMux I__3784 (
            .O(N__17772),
            .I(N__17753));
    InMux I__3783 (
            .O(N__17771),
            .I(N__17750));
    InMux I__3782 (
            .O(N__17770),
            .I(N__17747));
    LocalMux I__3781 (
            .O(N__17767),
            .I(N__17742));
    Span4Mux_h I__3780 (
            .O(N__17762),
            .I(N__17742));
    Span4Mux_h I__3779 (
            .O(N__17759),
            .I(N__17739));
    InMux I__3778 (
            .O(N__17758),
            .I(N__17736));
    LocalMux I__3777 (
            .O(N__17753),
            .I(N__17731));
    LocalMux I__3776 (
            .O(N__17750),
            .I(N__17731));
    LocalMux I__3775 (
            .O(N__17747),
            .I(N__17728));
    Span4Mux_v I__3774 (
            .O(N__17742),
            .I(N__17723));
    Span4Mux_v I__3773 (
            .O(N__17739),
            .I(N__17723));
    LocalMux I__3772 (
            .O(N__17736),
            .I(N__17720));
    Span4Mux_v I__3771 (
            .O(N__17731),
            .I(N__17715));
    Span4Mux_h I__3770 (
            .O(N__17728),
            .I(N__17715));
    Sp12to4 I__3769 (
            .O(N__17723),
            .I(N__17710));
    Span12Mux_h I__3768 (
            .O(N__17720),
            .I(N__17710));
    Span4Mux_v I__3767 (
            .O(N__17715),
            .I(N__17707));
    Odrv12 I__3766 (
            .O(N__17710),
            .I(TVP_VSYNC_c));
    Odrv4 I__3765 (
            .O(N__17707),
            .I(TVP_VSYNC_c));
    SRMux I__3764 (
            .O(N__17702),
            .I(N__17699));
    LocalMux I__3763 (
            .O(N__17699),
            .I(N__17694));
    SRMux I__3762 (
            .O(N__17698),
            .I(N__17691));
    SRMux I__3761 (
            .O(N__17697),
            .I(N__17687));
    Span4Mux_v I__3760 (
            .O(N__17694),
            .I(N__17682));
    LocalMux I__3759 (
            .O(N__17691),
            .I(N__17682));
    SRMux I__3758 (
            .O(N__17690),
            .I(N__17679));
    LocalMux I__3757 (
            .O(N__17687),
            .I(N__17676));
    Span4Mux_v I__3756 (
            .O(N__17682),
            .I(N__17670));
    LocalMux I__3755 (
            .O(N__17679),
            .I(N__17670));
    Span4Mux_v I__3754 (
            .O(N__17676),
            .I(N__17667));
    SRMux I__3753 (
            .O(N__17675),
            .I(N__17664));
    Span4Mux_h I__3752 (
            .O(N__17670),
            .I(N__17661));
    Span4Mux_v I__3751 (
            .O(N__17667),
            .I(N__17656));
    LocalMux I__3750 (
            .O(N__17664),
            .I(N__17656));
    Span4Mux_v I__3749 (
            .O(N__17661),
            .I(N__17653));
    Span4Mux_v I__3748 (
            .O(N__17656),
            .I(N__17650));
    Odrv4 I__3747 (
            .O(N__17653),
            .I(\receive_module.BRAM_ADDR_13__N_31 ));
    Odrv4 I__3746 (
            .O(N__17650),
            .I(\receive_module.BRAM_ADDR_13__N_31 ));
    SRMux I__3745 (
            .O(N__17645),
            .I(N__17640));
    SRMux I__3744 (
            .O(N__17644),
            .I(N__17635));
    CEMux I__3743 (
            .O(N__17643),
            .I(N__17632));
    LocalMux I__3742 (
            .O(N__17640),
            .I(N__17629));
    InMux I__3741 (
            .O(N__17639),
            .I(N__17626));
    CEMux I__3740 (
            .O(N__17638),
            .I(N__17623));
    LocalMux I__3739 (
            .O(N__17635),
            .I(N__17620));
    LocalMux I__3738 (
            .O(N__17632),
            .I(N__17617));
    Span4Mux_v I__3737 (
            .O(N__17629),
            .I(N__17612));
    LocalMux I__3736 (
            .O(N__17626),
            .I(N__17612));
    LocalMux I__3735 (
            .O(N__17623),
            .I(N__17609));
    Sp12to4 I__3734 (
            .O(N__17620),
            .I(N__17606));
    Span4Mux_h I__3733 (
            .O(N__17617),
            .I(N__17601));
    Span4Mux_h I__3732 (
            .O(N__17612),
            .I(N__17601));
    Odrv12 I__3731 (
            .O(N__17609),
            .I(\transmit_module.video_signal_controller.n2030 ));
    Odrv12 I__3730 (
            .O(N__17606),
            .I(\transmit_module.video_signal_controller.n2030 ));
    Odrv4 I__3729 (
            .O(N__17601),
            .I(\transmit_module.video_signal_controller.n2030 ));
    SRMux I__3728 (
            .O(N__17594),
            .I(N__17590));
    SRMux I__3727 (
            .O(N__17593),
            .I(N__17587));
    LocalMux I__3726 (
            .O(N__17590),
            .I(N__17584));
    LocalMux I__3725 (
            .O(N__17587),
            .I(N__17581));
    Span4Mux_h I__3724 (
            .O(N__17584),
            .I(N__17578));
    Odrv4 I__3723 (
            .O(N__17581),
            .I(\transmit_module.video_signal_controller.n2551 ));
    Odrv4 I__3722 (
            .O(N__17578),
            .I(\transmit_module.video_signal_controller.n2551 ));
    IoInMux I__3721 (
            .O(N__17573),
            .I(N__17570));
    LocalMux I__3720 (
            .O(N__17570),
            .I(N__17567));
    Span4Mux_s2_h I__3719 (
            .O(N__17567),
            .I(N__17564));
    Span4Mux_h I__3718 (
            .O(N__17564),
            .I(N__17561));
    Span4Mux_h I__3717 (
            .O(N__17561),
            .I(N__17557));
    InMux I__3716 (
            .O(N__17560),
            .I(N__17554));
    Span4Mux_v I__3715 (
            .O(N__17557),
            .I(N__17551));
    LocalMux I__3714 (
            .O(N__17554),
            .I(N__17548));
    Span4Mux_v I__3713 (
            .O(N__17551),
            .I(N__17543));
    Span4Mux_v I__3712 (
            .O(N__17548),
            .I(N__17543));
    Odrv4 I__3711 (
            .O(N__17543),
            .I(DEBUG_c_6));
    InMux I__3710 (
            .O(N__17540),
            .I(N__17537));
    LocalMux I__3709 (
            .O(N__17537),
            .I(\transmit_module.video_signal_controller.SYNC_BUFF1 ));
    InMux I__3708 (
            .O(N__17534),
            .I(N__17531));
    LocalMux I__3707 (
            .O(N__17531),
            .I(\transmit_module.video_signal_controller.SYNC_BUFF2 ));
    IoInMux I__3706 (
            .O(N__17528),
            .I(N__17525));
    LocalMux I__3705 (
            .O(N__17525),
            .I(N__17522));
    IoSpan4Mux I__3704 (
            .O(N__17522),
            .I(N__17519));
    Span4Mux_s3_h I__3703 (
            .O(N__17519),
            .I(N__17515));
    InMux I__3702 (
            .O(N__17518),
            .I(N__17512));
    Span4Mux_h I__3701 (
            .O(N__17515),
            .I(N__17509));
    LocalMux I__3700 (
            .O(N__17512),
            .I(N__17506));
    Span4Mux_h I__3699 (
            .O(N__17509),
            .I(N__17501));
    Span4Mux_v I__3698 (
            .O(N__17506),
            .I(N__17501));
    Odrv4 I__3697 (
            .O(N__17501),
            .I(n3852));
    CEMux I__3696 (
            .O(N__17498),
            .I(N__17494));
    CEMux I__3695 (
            .O(N__17497),
            .I(N__17491));
    LocalMux I__3694 (
            .O(N__17494),
            .I(N__17487));
    LocalMux I__3693 (
            .O(N__17491),
            .I(N__17484));
    InMux I__3692 (
            .O(N__17490),
            .I(N__17481));
    Span4Mux_h I__3691 (
            .O(N__17487),
            .I(N__17478));
    Span4Mux_h I__3690 (
            .O(N__17484),
            .I(N__17475));
    LocalMux I__3689 (
            .O(N__17481),
            .I(N__17472));
    Span4Mux_h I__3688 (
            .O(N__17478),
            .I(N__17469));
    Span4Mux_h I__3687 (
            .O(N__17475),
            .I(N__17464));
    Span4Mux_h I__3686 (
            .O(N__17472),
            .I(N__17464));
    Odrv4 I__3685 (
            .O(N__17469),
            .I(\transmit_module.n2039 ));
    Odrv4 I__3684 (
            .O(N__17464),
            .I(\transmit_module.n2039 ));
    InMux I__3683 (
            .O(N__17459),
            .I(N__17456));
    LocalMux I__3682 (
            .O(N__17456),
            .I(N__17453));
    Span4Mux_v I__3681 (
            .O(N__17453),
            .I(N__17450));
    Span4Mux_h I__3680 (
            .O(N__17450),
            .I(N__17447));
    Span4Mux_h I__3679 (
            .O(N__17447),
            .I(N__17444));
    Odrv4 I__3678 (
            .O(N__17444),
            .I(\line_buffer.n603 ));
    InMux I__3677 (
            .O(N__17441),
            .I(N__17438));
    LocalMux I__3676 (
            .O(N__17438),
            .I(N__17435));
    Span4Mux_v I__3675 (
            .O(N__17435),
            .I(N__17432));
    Sp12to4 I__3674 (
            .O(N__17432),
            .I(N__17429));
    Odrv12 I__3673 (
            .O(N__17429),
            .I(\line_buffer.n595 ));
    InMux I__3672 (
            .O(N__17426),
            .I(N__17423));
    LocalMux I__3671 (
            .O(N__17423),
            .I(N__17420));
    Span4Mux_v I__3670 (
            .O(N__17420),
            .I(N__17417));
    Span4Mux_h I__3669 (
            .O(N__17417),
            .I(N__17414));
    Span4Mux_h I__3668 (
            .O(N__17414),
            .I(N__17411));
    Span4Mux_v I__3667 (
            .O(N__17411),
            .I(N__17408));
    Odrv4 I__3666 (
            .O(N__17408),
            .I(\line_buffer.n569 ));
    CascadeMux I__3665 (
            .O(N__17405),
            .I(N__17402));
    InMux I__3664 (
            .O(N__17402),
            .I(N__17399));
    LocalMux I__3663 (
            .O(N__17399),
            .I(N__17396));
    Span4Mux_h I__3662 (
            .O(N__17396),
            .I(N__17393));
    Span4Mux_h I__3661 (
            .O(N__17393),
            .I(N__17390));
    Span4Mux_h I__3660 (
            .O(N__17390),
            .I(N__17387));
    Odrv4 I__3659 (
            .O(N__17387),
            .I(\line_buffer.n561 ));
    CascadeMux I__3658 (
            .O(N__17384),
            .I(\line_buffer.n3830_cascade_ ));
    InMux I__3657 (
            .O(N__17381),
            .I(N__17378));
    LocalMux I__3656 (
            .O(N__17378),
            .I(N__17375));
    Span4Mux_h I__3655 (
            .O(N__17375),
            .I(N__17372));
    Odrv4 I__3654 (
            .O(N__17372),
            .I(TX_DATA_1));
    InMux I__3653 (
            .O(N__17369),
            .I(N__17365));
    InMux I__3652 (
            .O(N__17368),
            .I(N__17361));
    LocalMux I__3651 (
            .O(N__17365),
            .I(N__17358));
    InMux I__3650 (
            .O(N__17364),
            .I(N__17355));
    LocalMux I__3649 (
            .O(N__17361),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    Odrv4 I__3648 (
            .O(N__17358),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    LocalMux I__3647 (
            .O(N__17355),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    InMux I__3646 (
            .O(N__17348),
            .I(N__17343));
    InMux I__3645 (
            .O(N__17347),
            .I(N__17340));
    InMux I__3644 (
            .O(N__17346),
            .I(N__17337));
    LocalMux I__3643 (
            .O(N__17343),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__3642 (
            .O(N__17340),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__3641 (
            .O(N__17337),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    InMux I__3640 (
            .O(N__17330),
            .I(N__17327));
    LocalMux I__3639 (
            .O(N__17327),
            .I(N__17324));
    Odrv4 I__3638 (
            .O(N__17324),
            .I(\transmit_module.video_signal_controller.n3858 ));
    CascadeMux I__3637 (
            .O(N__17321),
            .I(\transmit_module.n213_cascade_ ));
    InMux I__3636 (
            .O(N__17318),
            .I(N__17312));
    InMux I__3635 (
            .O(N__17317),
            .I(N__17307));
    InMux I__3634 (
            .O(N__17316),
            .I(N__17307));
    InMux I__3633 (
            .O(N__17315),
            .I(N__17304));
    LocalMux I__3632 (
            .O(N__17312),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__3631 (
            .O(N__17307),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__3630 (
            .O(N__17304),
            .I(\transmit_module.TX_ADDR_7 ));
    InMux I__3629 (
            .O(N__17297),
            .I(N__17294));
    LocalMux I__3628 (
            .O(N__17294),
            .I(\transmit_module.n184 ));
    InMux I__3627 (
            .O(N__17291),
            .I(N__17287));
    InMux I__3626 (
            .O(N__17290),
            .I(N__17284));
    LocalMux I__3625 (
            .O(N__17287),
            .I(\transmit_module.n216 ));
    LocalMux I__3624 (
            .O(N__17284),
            .I(\transmit_module.n216 ));
    CascadeMux I__3623 (
            .O(N__17279),
            .I(N__17275));
    CascadeMux I__3622 (
            .O(N__17278),
            .I(N__17272));
    CascadeBuf I__3621 (
            .O(N__17275),
            .I(N__17269));
    CascadeBuf I__3620 (
            .O(N__17272),
            .I(N__17266));
    CascadeMux I__3619 (
            .O(N__17269),
            .I(N__17263));
    CascadeMux I__3618 (
            .O(N__17266),
            .I(N__17260));
    CascadeBuf I__3617 (
            .O(N__17263),
            .I(N__17257));
    CascadeBuf I__3616 (
            .O(N__17260),
            .I(N__17254));
    CascadeMux I__3615 (
            .O(N__17257),
            .I(N__17251));
    CascadeMux I__3614 (
            .O(N__17254),
            .I(N__17248));
    CascadeBuf I__3613 (
            .O(N__17251),
            .I(N__17245));
    CascadeBuf I__3612 (
            .O(N__17248),
            .I(N__17242));
    CascadeMux I__3611 (
            .O(N__17245),
            .I(N__17239));
    CascadeMux I__3610 (
            .O(N__17242),
            .I(N__17236));
    CascadeBuf I__3609 (
            .O(N__17239),
            .I(N__17233));
    CascadeBuf I__3608 (
            .O(N__17236),
            .I(N__17230));
    CascadeMux I__3607 (
            .O(N__17233),
            .I(N__17227));
    CascadeMux I__3606 (
            .O(N__17230),
            .I(N__17224));
    CascadeBuf I__3605 (
            .O(N__17227),
            .I(N__17221));
    CascadeBuf I__3604 (
            .O(N__17224),
            .I(N__17218));
    CascadeMux I__3603 (
            .O(N__17221),
            .I(N__17215));
    CascadeMux I__3602 (
            .O(N__17218),
            .I(N__17212));
    CascadeBuf I__3601 (
            .O(N__17215),
            .I(N__17209));
    CascadeBuf I__3600 (
            .O(N__17212),
            .I(N__17206));
    CascadeMux I__3599 (
            .O(N__17209),
            .I(N__17203));
    CascadeMux I__3598 (
            .O(N__17206),
            .I(N__17200));
    CascadeBuf I__3597 (
            .O(N__17203),
            .I(N__17197));
    CascadeBuf I__3596 (
            .O(N__17200),
            .I(N__17194));
    CascadeMux I__3595 (
            .O(N__17197),
            .I(N__17191));
    CascadeMux I__3594 (
            .O(N__17194),
            .I(N__17188));
    CascadeBuf I__3593 (
            .O(N__17191),
            .I(N__17185));
    CascadeBuf I__3592 (
            .O(N__17188),
            .I(N__17182));
    CascadeMux I__3591 (
            .O(N__17185),
            .I(N__17179));
    CascadeMux I__3590 (
            .O(N__17182),
            .I(N__17176));
    CascadeBuf I__3589 (
            .O(N__17179),
            .I(N__17173));
    CascadeBuf I__3588 (
            .O(N__17176),
            .I(N__17170));
    CascadeMux I__3587 (
            .O(N__17173),
            .I(N__17167));
    CascadeMux I__3586 (
            .O(N__17170),
            .I(N__17164));
    CascadeBuf I__3585 (
            .O(N__17167),
            .I(N__17161));
    CascadeBuf I__3584 (
            .O(N__17164),
            .I(N__17158));
    CascadeMux I__3583 (
            .O(N__17161),
            .I(N__17155));
    CascadeMux I__3582 (
            .O(N__17158),
            .I(N__17152));
    CascadeBuf I__3581 (
            .O(N__17155),
            .I(N__17149));
    CascadeBuf I__3580 (
            .O(N__17152),
            .I(N__17146));
    CascadeMux I__3579 (
            .O(N__17149),
            .I(N__17143));
    CascadeMux I__3578 (
            .O(N__17146),
            .I(N__17140));
    CascadeBuf I__3577 (
            .O(N__17143),
            .I(N__17137));
    CascadeBuf I__3576 (
            .O(N__17140),
            .I(N__17134));
    CascadeMux I__3575 (
            .O(N__17137),
            .I(N__17131));
    CascadeMux I__3574 (
            .O(N__17134),
            .I(N__17128));
    CascadeBuf I__3573 (
            .O(N__17131),
            .I(N__17125));
    CascadeBuf I__3572 (
            .O(N__17128),
            .I(N__17122));
    CascadeMux I__3571 (
            .O(N__17125),
            .I(N__17119));
    CascadeMux I__3570 (
            .O(N__17122),
            .I(N__17116));
    CascadeBuf I__3569 (
            .O(N__17119),
            .I(N__17113));
    CascadeBuf I__3568 (
            .O(N__17116),
            .I(N__17110));
    CascadeMux I__3567 (
            .O(N__17113),
            .I(N__17107));
    CascadeMux I__3566 (
            .O(N__17110),
            .I(N__17104));
    CascadeBuf I__3565 (
            .O(N__17107),
            .I(N__17101));
    CascadeBuf I__3564 (
            .O(N__17104),
            .I(N__17098));
    CascadeMux I__3563 (
            .O(N__17101),
            .I(N__17095));
    CascadeMux I__3562 (
            .O(N__17098),
            .I(N__17092));
    InMux I__3561 (
            .O(N__17095),
            .I(N__17089));
    InMux I__3560 (
            .O(N__17092),
            .I(N__17086));
    LocalMux I__3559 (
            .O(N__17089),
            .I(N__17083));
    LocalMux I__3558 (
            .O(N__17086),
            .I(N__17080));
    Span12Mux_s10_h I__3557 (
            .O(N__17083),
            .I(N__17077));
    Span12Mux_s9_h I__3556 (
            .O(N__17080),
            .I(N__17074));
    Span12Mux_v I__3555 (
            .O(N__17077),
            .I(N__17069));
    Span12Mux_v I__3554 (
            .O(N__17074),
            .I(N__17069));
    Odrv12 I__3553 (
            .O(N__17069),
            .I(n24));
    InMux I__3552 (
            .O(N__17066),
            .I(N__17063));
    LocalMux I__3551 (
            .O(N__17063),
            .I(\transmit_module.ADDR_Y_COMPONENT_9 ));
    InMux I__3550 (
            .O(N__17060),
            .I(N__17056));
    InMux I__3549 (
            .O(N__17059),
            .I(N__17053));
    LocalMux I__3548 (
            .O(N__17056),
            .I(\transmit_module.n181 ));
    LocalMux I__3547 (
            .O(N__17053),
            .I(\transmit_module.n181 ));
    InMux I__3546 (
            .O(N__17048),
            .I(N__17045));
    LocalMux I__3545 (
            .O(N__17045),
            .I(\transmit_module.n213 ));
    CascadeMux I__3544 (
            .O(N__17042),
            .I(N__17038));
    CascadeMux I__3543 (
            .O(N__17041),
            .I(N__17035));
    CascadeBuf I__3542 (
            .O(N__17038),
            .I(N__17032));
    CascadeBuf I__3541 (
            .O(N__17035),
            .I(N__17029));
    CascadeMux I__3540 (
            .O(N__17032),
            .I(N__17026));
    CascadeMux I__3539 (
            .O(N__17029),
            .I(N__17023));
    CascadeBuf I__3538 (
            .O(N__17026),
            .I(N__17020));
    CascadeBuf I__3537 (
            .O(N__17023),
            .I(N__17017));
    CascadeMux I__3536 (
            .O(N__17020),
            .I(N__17014));
    CascadeMux I__3535 (
            .O(N__17017),
            .I(N__17011));
    CascadeBuf I__3534 (
            .O(N__17014),
            .I(N__17008));
    CascadeBuf I__3533 (
            .O(N__17011),
            .I(N__17005));
    CascadeMux I__3532 (
            .O(N__17008),
            .I(N__17002));
    CascadeMux I__3531 (
            .O(N__17005),
            .I(N__16999));
    CascadeBuf I__3530 (
            .O(N__17002),
            .I(N__16996));
    CascadeBuf I__3529 (
            .O(N__16999),
            .I(N__16993));
    CascadeMux I__3528 (
            .O(N__16996),
            .I(N__16990));
    CascadeMux I__3527 (
            .O(N__16993),
            .I(N__16987));
    CascadeBuf I__3526 (
            .O(N__16990),
            .I(N__16984));
    CascadeBuf I__3525 (
            .O(N__16987),
            .I(N__16981));
    CascadeMux I__3524 (
            .O(N__16984),
            .I(N__16978));
    CascadeMux I__3523 (
            .O(N__16981),
            .I(N__16975));
    CascadeBuf I__3522 (
            .O(N__16978),
            .I(N__16972));
    CascadeBuf I__3521 (
            .O(N__16975),
            .I(N__16969));
    CascadeMux I__3520 (
            .O(N__16972),
            .I(N__16966));
    CascadeMux I__3519 (
            .O(N__16969),
            .I(N__16963));
    CascadeBuf I__3518 (
            .O(N__16966),
            .I(N__16960));
    CascadeBuf I__3517 (
            .O(N__16963),
            .I(N__16957));
    CascadeMux I__3516 (
            .O(N__16960),
            .I(N__16954));
    CascadeMux I__3515 (
            .O(N__16957),
            .I(N__16951));
    CascadeBuf I__3514 (
            .O(N__16954),
            .I(N__16948));
    CascadeBuf I__3513 (
            .O(N__16951),
            .I(N__16945));
    CascadeMux I__3512 (
            .O(N__16948),
            .I(N__16942));
    CascadeMux I__3511 (
            .O(N__16945),
            .I(N__16939));
    CascadeBuf I__3510 (
            .O(N__16942),
            .I(N__16936));
    CascadeBuf I__3509 (
            .O(N__16939),
            .I(N__16933));
    CascadeMux I__3508 (
            .O(N__16936),
            .I(N__16930));
    CascadeMux I__3507 (
            .O(N__16933),
            .I(N__16927));
    CascadeBuf I__3506 (
            .O(N__16930),
            .I(N__16924));
    CascadeBuf I__3505 (
            .O(N__16927),
            .I(N__16921));
    CascadeMux I__3504 (
            .O(N__16924),
            .I(N__16918));
    CascadeMux I__3503 (
            .O(N__16921),
            .I(N__16915));
    CascadeBuf I__3502 (
            .O(N__16918),
            .I(N__16912));
    CascadeBuf I__3501 (
            .O(N__16915),
            .I(N__16909));
    CascadeMux I__3500 (
            .O(N__16912),
            .I(N__16906));
    CascadeMux I__3499 (
            .O(N__16909),
            .I(N__16903));
    CascadeBuf I__3498 (
            .O(N__16906),
            .I(N__16900));
    CascadeBuf I__3497 (
            .O(N__16903),
            .I(N__16897));
    CascadeMux I__3496 (
            .O(N__16900),
            .I(N__16894));
    CascadeMux I__3495 (
            .O(N__16897),
            .I(N__16891));
    CascadeBuf I__3494 (
            .O(N__16894),
            .I(N__16888));
    CascadeBuf I__3493 (
            .O(N__16891),
            .I(N__16885));
    CascadeMux I__3492 (
            .O(N__16888),
            .I(N__16882));
    CascadeMux I__3491 (
            .O(N__16885),
            .I(N__16879));
    CascadeBuf I__3490 (
            .O(N__16882),
            .I(N__16876));
    CascadeBuf I__3489 (
            .O(N__16879),
            .I(N__16873));
    CascadeMux I__3488 (
            .O(N__16876),
            .I(N__16870));
    CascadeMux I__3487 (
            .O(N__16873),
            .I(N__16867));
    CascadeBuf I__3486 (
            .O(N__16870),
            .I(N__16864));
    CascadeBuf I__3485 (
            .O(N__16867),
            .I(N__16861));
    CascadeMux I__3484 (
            .O(N__16864),
            .I(N__16858));
    CascadeMux I__3483 (
            .O(N__16861),
            .I(N__16855));
    InMux I__3482 (
            .O(N__16858),
            .I(N__16852));
    InMux I__3481 (
            .O(N__16855),
            .I(N__16849));
    LocalMux I__3480 (
            .O(N__16852),
            .I(N__16846));
    LocalMux I__3479 (
            .O(N__16849),
            .I(N__16843));
    Span12Mux_h I__3478 (
            .O(N__16846),
            .I(N__16838));
    Span12Mux_h I__3477 (
            .O(N__16843),
            .I(N__16838));
    Span12Mux_v I__3476 (
            .O(N__16838),
            .I(N__16835));
    Odrv12 I__3475 (
            .O(N__16835),
            .I(n21));
    InMux I__3474 (
            .O(N__16832),
            .I(N__16829));
    LocalMux I__3473 (
            .O(N__16829),
            .I(N__16826));
    Span4Mux_h I__3472 (
            .O(N__16826),
            .I(N__16823));
    Span4Mux_v I__3471 (
            .O(N__16823),
            .I(N__16820));
    Span4Mux_h I__3470 (
            .O(N__16820),
            .I(N__16817));
    Span4Mux_h I__3469 (
            .O(N__16817),
            .I(N__16814));
    Odrv4 I__3468 (
            .O(N__16814),
            .I(\line_buffer.n509 ));
    CascadeMux I__3467 (
            .O(N__16811),
            .I(N__16808));
    InMux I__3466 (
            .O(N__16808),
            .I(N__16805));
    LocalMux I__3465 (
            .O(N__16805),
            .I(N__16802));
    Span4Mux_v I__3464 (
            .O(N__16802),
            .I(N__16799));
    Span4Mux_v I__3463 (
            .O(N__16799),
            .I(N__16796));
    Span4Mux_h I__3462 (
            .O(N__16796),
            .I(N__16793));
    Odrv4 I__3461 (
            .O(N__16793),
            .I(\line_buffer.n501 ));
    InMux I__3460 (
            .O(N__16790),
            .I(N__16787));
    LocalMux I__3459 (
            .O(N__16787),
            .I(\line_buffer.n3770 ));
    InMux I__3458 (
            .O(N__16784),
            .I(N__16781));
    LocalMux I__3457 (
            .O(N__16781),
            .I(N__16778));
    Span4Mux_v I__3456 (
            .O(N__16778),
            .I(N__16775));
    Span4Mux_h I__3455 (
            .O(N__16775),
            .I(N__16772));
    Span4Mux_h I__3454 (
            .O(N__16772),
            .I(N__16769));
    Odrv4 I__3453 (
            .O(N__16769),
            .I(\line_buffer.n571 ));
    InMux I__3452 (
            .O(N__16766),
            .I(N__16763));
    LocalMux I__3451 (
            .O(N__16763),
            .I(N__16760));
    Span12Mux_h I__3450 (
            .O(N__16760),
            .I(N__16757));
    Odrv12 I__3449 (
            .O(N__16757),
            .I(\line_buffer.n563 ));
    InMux I__3448 (
            .O(N__16754),
            .I(N__16751));
    LocalMux I__3447 (
            .O(N__16751),
            .I(\receive_module.rx_counter.n11 ));
    IoInMux I__3446 (
            .O(N__16748),
            .I(N__16745));
    LocalMux I__3445 (
            .O(N__16745),
            .I(N__16742));
    Span4Mux_s1_v I__3444 (
            .O(N__16742),
            .I(N__16739));
    Span4Mux_v I__3443 (
            .O(N__16739),
            .I(N__16736));
    Span4Mux_v I__3442 (
            .O(N__16736),
            .I(N__16733));
    Span4Mux_h I__3441 (
            .O(N__16733),
            .I(N__16729));
    InMux I__3440 (
            .O(N__16732),
            .I(N__16726));
    Odrv4 I__3439 (
            .O(N__16729),
            .I(LED_c));
    LocalMux I__3438 (
            .O(N__16726),
            .I(LED_c));
    CEMux I__3437 (
            .O(N__16721),
            .I(N__16717));
    CEMux I__3436 (
            .O(N__16720),
            .I(N__16714));
    LocalMux I__3435 (
            .O(N__16717),
            .I(\receive_module.rx_counter.n3862 ));
    LocalMux I__3434 (
            .O(N__16714),
            .I(\receive_module.rx_counter.n3862 ));
    InMux I__3433 (
            .O(N__16709),
            .I(N__16706));
    LocalMux I__3432 (
            .O(N__16706),
            .I(N__16703));
    Span4Mux_h I__3431 (
            .O(N__16703),
            .I(N__16697));
    InMux I__3430 (
            .O(N__16702),
            .I(N__16692));
    InMux I__3429 (
            .O(N__16701),
            .I(N__16692));
    InMux I__3428 (
            .O(N__16700),
            .I(N__16689));
    Odrv4 I__3427 (
            .O(N__16697),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__3426 (
            .O(N__16692),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__3425 (
            .O(N__16689),
            .I(\transmit_module.TX_ADDR_6 ));
    InMux I__3424 (
            .O(N__16682),
            .I(N__16679));
    LocalMux I__3423 (
            .O(N__16679),
            .I(N__16676));
    Span4Mux_h I__3422 (
            .O(N__16676),
            .I(N__16673));
    Odrv4 I__3421 (
            .O(N__16673),
            .I(\transmit_module.ADDR_Y_COMPONENT_6 ));
    InMux I__3420 (
            .O(N__16670),
            .I(N__16664));
    InMux I__3419 (
            .O(N__16669),
            .I(N__16659));
    InMux I__3418 (
            .O(N__16668),
            .I(N__16659));
    InMux I__3417 (
            .O(N__16667),
            .I(N__16656));
    LocalMux I__3416 (
            .O(N__16664),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__3415 (
            .O(N__16659),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__3414 (
            .O(N__16656),
            .I(\transmit_module.TX_ADDR_2 ));
    InMux I__3413 (
            .O(N__16649),
            .I(N__16646));
    LocalMux I__3412 (
            .O(N__16646),
            .I(\transmit_module.ADDR_Y_COMPONENT_2 ));
    InMux I__3411 (
            .O(N__16643),
            .I(N__16640));
    LocalMux I__3410 (
            .O(N__16640),
            .I(\transmit_module.ADDR_Y_COMPONENT_7 ));
    InMux I__3409 (
            .O(N__16637),
            .I(N__16634));
    LocalMux I__3408 (
            .O(N__16634),
            .I(\transmit_module.ADDR_Y_COMPONENT_4 ));
    CascadeMux I__3407 (
            .O(N__16631),
            .I(\transmit_module.n184_cascade_ ));
    InMux I__3406 (
            .O(N__16628),
            .I(N__16625));
    LocalMux I__3405 (
            .O(N__16625),
            .I(\transmit_module.n200 ));
    InMux I__3404 (
            .O(N__16622),
            .I(N__16616));
    InMux I__3403 (
            .O(N__16621),
            .I(N__16611));
    InMux I__3402 (
            .O(N__16620),
            .I(N__16611));
    InMux I__3401 (
            .O(N__16619),
            .I(N__16608));
    LocalMux I__3400 (
            .O(N__16616),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__3399 (
            .O(N__16611),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__3398 (
            .O(N__16608),
            .I(\transmit_module.TX_ADDR_4 ));
    InMux I__3397 (
            .O(N__16601),
            .I(N__16598));
    LocalMux I__3396 (
            .O(N__16598),
            .I(\transmit_module.n197 ));
    InMux I__3395 (
            .O(N__16595),
            .I(N__16592));
    LocalMux I__3394 (
            .O(N__16592),
            .I(N__16589));
    Span4Mux_v I__3393 (
            .O(N__16589),
            .I(N__16585));
    InMux I__3392 (
            .O(N__16588),
            .I(N__16582));
    Odrv4 I__3391 (
            .O(N__16585),
            .I(\transmit_module.n188 ));
    LocalMux I__3390 (
            .O(N__16582),
            .I(\transmit_module.n188 ));
    InMux I__3389 (
            .O(N__16577),
            .I(N__16572));
    InMux I__3388 (
            .O(N__16576),
            .I(N__16569));
    InMux I__3387 (
            .O(N__16575),
            .I(N__16565));
    LocalMux I__3386 (
            .O(N__16572),
            .I(N__16560));
    LocalMux I__3385 (
            .O(N__16569),
            .I(N__16560));
    InMux I__3384 (
            .O(N__16568),
            .I(N__16557));
    LocalMux I__3383 (
            .O(N__16565),
            .I(N__16554));
    Span4Mux_v I__3382 (
            .O(N__16560),
            .I(N__16551));
    LocalMux I__3381 (
            .O(N__16557),
            .I(\transmit_module.n3859 ));
    Odrv4 I__3380 (
            .O(N__16554),
            .I(\transmit_module.n3859 ));
    Odrv4 I__3379 (
            .O(N__16551),
            .I(\transmit_module.n3859 ));
    InMux I__3378 (
            .O(N__16544),
            .I(N__16540));
    InMux I__3377 (
            .O(N__16543),
            .I(N__16535));
    LocalMux I__3376 (
            .O(N__16540),
            .I(N__16532));
    InMux I__3375 (
            .O(N__16539),
            .I(N__16529));
    InMux I__3374 (
            .O(N__16538),
            .I(N__16526));
    LocalMux I__3373 (
            .O(N__16535),
            .I(\transmit_module.TX_ADDR_1 ));
    Odrv4 I__3372 (
            .O(N__16532),
            .I(\transmit_module.TX_ADDR_1 ));
    LocalMux I__3371 (
            .O(N__16529),
            .I(\transmit_module.TX_ADDR_1 ));
    LocalMux I__3370 (
            .O(N__16526),
            .I(\transmit_module.TX_ADDR_1 ));
    InMux I__3369 (
            .O(N__16517),
            .I(N__16514));
    LocalMux I__3368 (
            .O(N__16514),
            .I(\transmit_module.ADDR_Y_COMPONENT_1 ));
    CascadeMux I__3367 (
            .O(N__16511),
            .I(N__16508));
    InMux I__3366 (
            .O(N__16508),
            .I(N__16505));
    LocalMux I__3365 (
            .O(N__16505),
            .I(N__16502));
    Span4Mux_h I__3364 (
            .O(N__16502),
            .I(N__16499));
    Odrv4 I__3363 (
            .O(N__16499),
            .I(\transmit_module.ADDR_Y_COMPONENT_11 ));
    CascadeMux I__3362 (
            .O(N__16496),
            .I(N__16493));
    InMux I__3361 (
            .O(N__16493),
            .I(N__16490));
    LocalMux I__3360 (
            .O(N__16490),
            .I(N__16487));
    Span4Mux_h I__3359 (
            .O(N__16487),
            .I(N__16484));
    Odrv4 I__3358 (
            .O(N__16484),
            .I(\transmit_module.ADDR_Y_COMPONENT_12 ));
    InMux I__3357 (
            .O(N__16481),
            .I(N__16478));
    LocalMux I__3356 (
            .O(N__16478),
            .I(N__16475));
    Odrv12 I__3355 (
            .O(N__16475),
            .I(\transmit_module.ADDR_Y_COMPONENT_13 ));
    InMux I__3354 (
            .O(N__16472),
            .I(N__16467));
    InMux I__3353 (
            .O(N__16471),
            .I(N__16464));
    InMux I__3352 (
            .O(N__16470),
            .I(N__16460));
    LocalMux I__3351 (
            .O(N__16467),
            .I(N__16455));
    LocalMux I__3350 (
            .O(N__16464),
            .I(N__16455));
    InMux I__3349 (
            .O(N__16463),
            .I(N__16452));
    LocalMux I__3348 (
            .O(N__16460),
            .I(\transmit_module.TX_ADDR_0 ));
    Odrv4 I__3347 (
            .O(N__16455),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__3346 (
            .O(N__16452),
            .I(\transmit_module.TX_ADDR_0 ));
    InMux I__3345 (
            .O(N__16445),
            .I(N__16442));
    LocalMux I__3344 (
            .O(N__16442),
            .I(\transmit_module.ADDR_Y_COMPONENT_0 ));
    InMux I__3343 (
            .O(N__16439),
            .I(N__16436));
    LocalMux I__3342 (
            .O(N__16436),
            .I(N__16432));
    InMux I__3341 (
            .O(N__16435),
            .I(N__16428));
    Span4Mux_h I__3340 (
            .O(N__16432),
            .I(N__16424));
    InMux I__3339 (
            .O(N__16431),
            .I(N__16421));
    LocalMux I__3338 (
            .O(N__16428),
            .I(N__16418));
    InMux I__3337 (
            .O(N__16427),
            .I(N__16415));
    Odrv4 I__3336 (
            .O(N__16424),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__3335 (
            .O(N__16421),
            .I(\transmit_module.TX_ADDR_5 ));
    Odrv4 I__3334 (
            .O(N__16418),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__3333 (
            .O(N__16415),
            .I(\transmit_module.TX_ADDR_5 ));
    InMux I__3332 (
            .O(N__16406),
            .I(N__16403));
    LocalMux I__3331 (
            .O(N__16403),
            .I(N__16400));
    Odrv4 I__3330 (
            .O(N__16400),
            .I(\transmit_module.ADDR_Y_COMPONENT_5 ));
    CascadeMux I__3329 (
            .O(N__16397),
            .I(N__16394));
    InMux I__3328 (
            .O(N__16394),
            .I(N__16390));
    InMux I__3327 (
            .O(N__16393),
            .I(N__16385));
    LocalMux I__3326 (
            .O(N__16390),
            .I(N__16382));
    InMux I__3325 (
            .O(N__16389),
            .I(N__16377));
    InMux I__3324 (
            .O(N__16388),
            .I(N__16377));
    LocalMux I__3323 (
            .O(N__16385),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    Odrv4 I__3322 (
            .O(N__16382),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__3321 (
            .O(N__16377),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    InMux I__3320 (
            .O(N__16370),
            .I(\transmit_module.video_signal_controller.n3369 ));
    InMux I__3319 (
            .O(N__16367),
            .I(N__16362));
    InMux I__3318 (
            .O(N__16366),
            .I(N__16359));
    InMux I__3317 (
            .O(N__16365),
            .I(N__16356));
    LocalMux I__3316 (
            .O(N__16362),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__3315 (
            .O(N__16359),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__3314 (
            .O(N__16356),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    InMux I__3313 (
            .O(N__16349),
            .I(\transmit_module.video_signal_controller.n3370 ));
    InMux I__3312 (
            .O(N__16346),
            .I(N__16341));
    InMux I__3311 (
            .O(N__16345),
            .I(N__16338));
    InMux I__3310 (
            .O(N__16344),
            .I(N__16335));
    LocalMux I__3309 (
            .O(N__16341),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__3308 (
            .O(N__16338),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__3307 (
            .O(N__16335),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    InMux I__3306 (
            .O(N__16328),
            .I(\transmit_module.video_signal_controller.n3371 ));
    InMux I__3305 (
            .O(N__16325),
            .I(N__16321));
    InMux I__3304 (
            .O(N__16324),
            .I(N__16318));
    LocalMux I__3303 (
            .O(N__16321),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    LocalMux I__3302 (
            .O(N__16318),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    InMux I__3301 (
            .O(N__16313),
            .I(\transmit_module.video_signal_controller.n3372 ));
    InMux I__3300 (
            .O(N__16310),
            .I(N__16306));
    InMux I__3299 (
            .O(N__16309),
            .I(N__16303));
    LocalMux I__3298 (
            .O(N__16306),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    LocalMux I__3297 (
            .O(N__16303),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    InMux I__3296 (
            .O(N__16298),
            .I(bfn_14_14_0_));
    InMux I__3295 (
            .O(N__16295),
            .I(N__16290));
    InMux I__3294 (
            .O(N__16294),
            .I(N__16285));
    InMux I__3293 (
            .O(N__16293),
            .I(N__16285));
    LocalMux I__3292 (
            .O(N__16290),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    LocalMux I__3291 (
            .O(N__16285),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    InMux I__3290 (
            .O(N__16280),
            .I(\transmit_module.video_signal_controller.n3374 ));
    InMux I__3289 (
            .O(N__16277),
            .I(\transmit_module.video_signal_controller.n3375 ));
    InMux I__3288 (
            .O(N__16274),
            .I(\transmit_module.video_signal_controller.n3376 ));
    CascadeMux I__3287 (
            .O(N__16271),
            .I(N__16268));
    InMux I__3286 (
            .O(N__16268),
            .I(N__16265));
    LocalMux I__3285 (
            .O(N__16265),
            .I(N__16262));
    Span4Mux_v I__3284 (
            .O(N__16262),
            .I(N__16255));
    InMux I__3283 (
            .O(N__16261),
            .I(N__16250));
    InMux I__3282 (
            .O(N__16260),
            .I(N__16250));
    InMux I__3281 (
            .O(N__16259),
            .I(N__16247));
    InMux I__3280 (
            .O(N__16258),
            .I(N__16244));
    Odrv4 I__3279 (
            .O(N__16255),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__3278 (
            .O(N__16250),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__3277 (
            .O(N__16247),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__3276 (
            .O(N__16244),
            .I(\transmit_module.old_VGA_HS ));
    IoInMux I__3275 (
            .O(N__16235),
            .I(N__16232));
    LocalMux I__3274 (
            .O(N__16232),
            .I(N__16229));
    Span4Mux_s0_h I__3273 (
            .O(N__16229),
            .I(N__16225));
    InMux I__3272 (
            .O(N__16228),
            .I(N__16222));
    Sp12to4 I__3271 (
            .O(N__16225),
            .I(N__16217));
    LocalMux I__3270 (
            .O(N__16222),
            .I(N__16214));
    CascadeMux I__3269 (
            .O(N__16221),
            .I(N__16210));
    InMux I__3268 (
            .O(N__16220),
            .I(N__16205));
    Span12Mux_v I__3267 (
            .O(N__16217),
            .I(N__16202));
    Span4Mux_h I__3266 (
            .O(N__16214),
            .I(N__16199));
    InMux I__3265 (
            .O(N__16213),
            .I(N__16194));
    InMux I__3264 (
            .O(N__16210),
            .I(N__16194));
    InMux I__3263 (
            .O(N__16209),
            .I(N__16189));
    InMux I__3262 (
            .O(N__16208),
            .I(N__16189));
    LocalMux I__3261 (
            .O(N__16205),
            .I(N__16186));
    Odrv12 I__3260 (
            .O(N__16202),
            .I(ADV_HSYNC_c));
    Odrv4 I__3259 (
            .O(N__16199),
            .I(ADV_HSYNC_c));
    LocalMux I__3258 (
            .O(N__16194),
            .I(ADV_HSYNC_c));
    LocalMux I__3257 (
            .O(N__16189),
            .I(ADV_HSYNC_c));
    Odrv4 I__3256 (
            .O(N__16186),
            .I(ADV_HSYNC_c));
    CascadeMux I__3255 (
            .O(N__16175),
            .I(N__16171));
    CascadeMux I__3254 (
            .O(N__16174),
            .I(N__16168));
    CascadeBuf I__3253 (
            .O(N__16171),
            .I(N__16165));
    CascadeBuf I__3252 (
            .O(N__16168),
            .I(N__16162));
    CascadeMux I__3251 (
            .O(N__16165),
            .I(N__16159));
    CascadeMux I__3250 (
            .O(N__16162),
            .I(N__16156));
    CascadeBuf I__3249 (
            .O(N__16159),
            .I(N__16153));
    CascadeBuf I__3248 (
            .O(N__16156),
            .I(N__16150));
    CascadeMux I__3247 (
            .O(N__16153),
            .I(N__16147));
    CascadeMux I__3246 (
            .O(N__16150),
            .I(N__16144));
    CascadeBuf I__3245 (
            .O(N__16147),
            .I(N__16141));
    CascadeBuf I__3244 (
            .O(N__16144),
            .I(N__16138));
    CascadeMux I__3243 (
            .O(N__16141),
            .I(N__16135));
    CascadeMux I__3242 (
            .O(N__16138),
            .I(N__16132));
    CascadeBuf I__3241 (
            .O(N__16135),
            .I(N__16129));
    CascadeBuf I__3240 (
            .O(N__16132),
            .I(N__16126));
    CascadeMux I__3239 (
            .O(N__16129),
            .I(N__16123));
    CascadeMux I__3238 (
            .O(N__16126),
            .I(N__16120));
    CascadeBuf I__3237 (
            .O(N__16123),
            .I(N__16117));
    CascadeBuf I__3236 (
            .O(N__16120),
            .I(N__16114));
    CascadeMux I__3235 (
            .O(N__16117),
            .I(N__16111));
    CascadeMux I__3234 (
            .O(N__16114),
            .I(N__16108));
    CascadeBuf I__3233 (
            .O(N__16111),
            .I(N__16105));
    CascadeBuf I__3232 (
            .O(N__16108),
            .I(N__16102));
    CascadeMux I__3231 (
            .O(N__16105),
            .I(N__16099));
    CascadeMux I__3230 (
            .O(N__16102),
            .I(N__16096));
    CascadeBuf I__3229 (
            .O(N__16099),
            .I(N__16093));
    CascadeBuf I__3228 (
            .O(N__16096),
            .I(N__16090));
    CascadeMux I__3227 (
            .O(N__16093),
            .I(N__16087));
    CascadeMux I__3226 (
            .O(N__16090),
            .I(N__16084));
    CascadeBuf I__3225 (
            .O(N__16087),
            .I(N__16081));
    CascadeBuf I__3224 (
            .O(N__16084),
            .I(N__16078));
    CascadeMux I__3223 (
            .O(N__16081),
            .I(N__16075));
    CascadeMux I__3222 (
            .O(N__16078),
            .I(N__16072));
    CascadeBuf I__3221 (
            .O(N__16075),
            .I(N__16069));
    CascadeBuf I__3220 (
            .O(N__16072),
            .I(N__16066));
    CascadeMux I__3219 (
            .O(N__16069),
            .I(N__16063));
    CascadeMux I__3218 (
            .O(N__16066),
            .I(N__16060));
    CascadeBuf I__3217 (
            .O(N__16063),
            .I(N__16057));
    CascadeBuf I__3216 (
            .O(N__16060),
            .I(N__16054));
    CascadeMux I__3215 (
            .O(N__16057),
            .I(N__16051));
    CascadeMux I__3214 (
            .O(N__16054),
            .I(N__16048));
    CascadeBuf I__3213 (
            .O(N__16051),
            .I(N__16045));
    CascadeBuf I__3212 (
            .O(N__16048),
            .I(N__16042));
    CascadeMux I__3211 (
            .O(N__16045),
            .I(N__16039));
    CascadeMux I__3210 (
            .O(N__16042),
            .I(N__16036));
    CascadeBuf I__3209 (
            .O(N__16039),
            .I(N__16033));
    CascadeBuf I__3208 (
            .O(N__16036),
            .I(N__16030));
    CascadeMux I__3207 (
            .O(N__16033),
            .I(N__16027));
    CascadeMux I__3206 (
            .O(N__16030),
            .I(N__16024));
    CascadeBuf I__3205 (
            .O(N__16027),
            .I(N__16021));
    CascadeBuf I__3204 (
            .O(N__16024),
            .I(N__16018));
    CascadeMux I__3203 (
            .O(N__16021),
            .I(N__16015));
    CascadeMux I__3202 (
            .O(N__16018),
            .I(N__16012));
    CascadeBuf I__3201 (
            .O(N__16015),
            .I(N__16009));
    CascadeBuf I__3200 (
            .O(N__16012),
            .I(N__16006));
    CascadeMux I__3199 (
            .O(N__16009),
            .I(N__16003));
    CascadeMux I__3198 (
            .O(N__16006),
            .I(N__16000));
    CascadeBuf I__3197 (
            .O(N__16003),
            .I(N__15997));
    CascadeBuf I__3196 (
            .O(N__16000),
            .I(N__15994));
    CascadeMux I__3195 (
            .O(N__15997),
            .I(N__15991));
    CascadeMux I__3194 (
            .O(N__15994),
            .I(N__15988));
    InMux I__3193 (
            .O(N__15991),
            .I(N__15985));
    InMux I__3192 (
            .O(N__15988),
            .I(N__15982));
    LocalMux I__3191 (
            .O(N__15985),
            .I(N__15979));
    LocalMux I__3190 (
            .O(N__15982),
            .I(N__15976));
    Span4Mux_h I__3189 (
            .O(N__15979),
            .I(N__15972));
    Span4Mux_h I__3188 (
            .O(N__15976),
            .I(N__15969));
    InMux I__3187 (
            .O(N__15975),
            .I(N__15966));
    Sp12to4 I__3186 (
            .O(N__15972),
            .I(N__15963));
    Sp12to4 I__3185 (
            .O(N__15969),
            .I(N__15960));
    LocalMux I__3184 (
            .O(N__15966),
            .I(N__15957));
    Span12Mux_s9_v I__3183 (
            .O(N__15963),
            .I(N__15953));
    Span12Mux_s9_v I__3182 (
            .O(N__15960),
            .I(N__15950));
    Span4Mux_v I__3181 (
            .O(N__15957),
            .I(N__15947));
    InMux I__3180 (
            .O(N__15956),
            .I(N__15944));
    Span12Mux_v I__3179 (
            .O(N__15953),
            .I(N__15939));
    Span12Mux_v I__3178 (
            .O(N__15950),
            .I(N__15939));
    Odrv4 I__3177 (
            .O(N__15947),
            .I(RX_ADDR_10));
    LocalMux I__3176 (
            .O(N__15944),
            .I(RX_ADDR_10));
    Odrv12 I__3175 (
            .O(N__15939),
            .I(RX_ADDR_10));
    InMux I__3174 (
            .O(N__15932),
            .I(N__15929));
    LocalMux I__3173 (
            .O(N__15929),
            .I(N__15926));
    Span4Mux_h I__3172 (
            .O(N__15926),
            .I(N__15923));
    Odrv4 I__3171 (
            .O(N__15923),
            .I(\receive_module.n126 ));
    InMux I__3170 (
            .O(N__15920),
            .I(\receive_module.n3332 ));
    InMux I__3169 (
            .O(N__15917),
            .I(N__15900));
    InMux I__3168 (
            .O(N__15916),
            .I(N__15900));
    InMux I__3167 (
            .O(N__15915),
            .I(N__15900));
    InMux I__3166 (
            .O(N__15914),
            .I(N__15900));
    InMux I__3165 (
            .O(N__15913),
            .I(N__15895));
    InMux I__3164 (
            .O(N__15912),
            .I(N__15895));
    InMux I__3163 (
            .O(N__15911),
            .I(N__15892));
    InMux I__3162 (
            .O(N__15910),
            .I(N__15889));
    InMux I__3161 (
            .O(N__15909),
            .I(N__15886));
    LocalMux I__3160 (
            .O(N__15900),
            .I(N__15879));
    LocalMux I__3159 (
            .O(N__15895),
            .I(N__15879));
    LocalMux I__3158 (
            .O(N__15892),
            .I(N__15879));
    LocalMux I__3157 (
            .O(N__15889),
            .I(N__15876));
    LocalMux I__3156 (
            .O(N__15886),
            .I(N__15871));
    Span4Mux_v I__3155 (
            .O(N__15879),
            .I(N__15871));
    Span4Mux_h I__3154 (
            .O(N__15876),
            .I(N__15868));
    Odrv4 I__3153 (
            .O(N__15871),
            .I(RX_ADDR_11));
    Odrv4 I__3152 (
            .O(N__15868),
            .I(RX_ADDR_11));
    InMux I__3151 (
            .O(N__15863),
            .I(\receive_module.n3333 ));
    CascadeMux I__3150 (
            .O(N__15860),
            .I(N__15856));
    InMux I__3149 (
            .O(N__15859),
            .I(N__15848));
    InMux I__3148 (
            .O(N__15856),
            .I(N__15848));
    CascadeMux I__3147 (
            .O(N__15855),
            .I(N__15844));
    CascadeMux I__3146 (
            .O(N__15854),
            .I(N__15841));
    InMux I__3145 (
            .O(N__15853),
            .I(N__15836));
    LocalMux I__3144 (
            .O(N__15848),
            .I(N__15833));
    InMux I__3143 (
            .O(N__15847),
            .I(N__15830));
    InMux I__3142 (
            .O(N__15844),
            .I(N__15820));
    InMux I__3141 (
            .O(N__15841),
            .I(N__15820));
    InMux I__3140 (
            .O(N__15840),
            .I(N__15820));
    InMux I__3139 (
            .O(N__15839),
            .I(N__15820));
    LocalMux I__3138 (
            .O(N__15836),
            .I(N__15817));
    Span4Mux_v I__3137 (
            .O(N__15833),
            .I(N__15814));
    LocalMux I__3136 (
            .O(N__15830),
            .I(N__15811));
    InMux I__3135 (
            .O(N__15829),
            .I(N__15808));
    LocalMux I__3134 (
            .O(N__15820),
            .I(N__15805));
    Span4Mux_h I__3133 (
            .O(N__15817),
            .I(N__15802));
    Span4Mux_h I__3132 (
            .O(N__15814),
            .I(N__15797));
    Span4Mux_v I__3131 (
            .O(N__15811),
            .I(N__15797));
    LocalMux I__3130 (
            .O(N__15808),
            .I(RX_ADDR_12));
    Odrv4 I__3129 (
            .O(N__15805),
            .I(RX_ADDR_12));
    Odrv4 I__3128 (
            .O(N__15802),
            .I(RX_ADDR_12));
    Odrv4 I__3127 (
            .O(N__15797),
            .I(RX_ADDR_12));
    InMux I__3126 (
            .O(N__15788),
            .I(\receive_module.n3334 ));
    CEMux I__3125 (
            .O(N__15785),
            .I(N__15782));
    LocalMux I__3124 (
            .O(N__15782),
            .I(N__15779));
    Span4Mux_h I__3123 (
            .O(N__15779),
            .I(N__15776));
    Odrv4 I__3122 (
            .O(N__15776),
            .I(\receive_module.n3854 ));
    IoInMux I__3121 (
            .O(N__15773),
            .I(N__15770));
    LocalMux I__3120 (
            .O(N__15770),
            .I(N__15767));
    Span4Mux_s2_h I__3119 (
            .O(N__15767),
            .I(N__15761));
    InMux I__3118 (
            .O(N__15766),
            .I(N__15756));
    CascadeMux I__3117 (
            .O(N__15765),
            .I(N__15753));
    CascadeMux I__3116 (
            .O(N__15764),
            .I(N__15748));
    Span4Mux_h I__3115 (
            .O(N__15761),
            .I(N__15743));
    CascadeMux I__3114 (
            .O(N__15760),
            .I(N__15740));
    CascadeMux I__3113 (
            .O(N__15759),
            .I(N__15736));
    LocalMux I__3112 (
            .O(N__15756),
            .I(N__15733));
    InMux I__3111 (
            .O(N__15753),
            .I(N__15728));
    InMux I__3110 (
            .O(N__15752),
            .I(N__15728));
    InMux I__3109 (
            .O(N__15751),
            .I(N__15719));
    InMux I__3108 (
            .O(N__15748),
            .I(N__15719));
    InMux I__3107 (
            .O(N__15747),
            .I(N__15719));
    InMux I__3106 (
            .O(N__15746),
            .I(N__15719));
    Span4Mux_h I__3105 (
            .O(N__15743),
            .I(N__15716));
    InMux I__3104 (
            .O(N__15740),
            .I(N__15713));
    InMux I__3103 (
            .O(N__15739),
            .I(N__15708));
    InMux I__3102 (
            .O(N__15736),
            .I(N__15708));
    Span4Mux_h I__3101 (
            .O(N__15733),
            .I(N__15701));
    LocalMux I__3100 (
            .O(N__15728),
            .I(N__15701));
    LocalMux I__3099 (
            .O(N__15719),
            .I(N__15701));
    Odrv4 I__3098 (
            .O(N__15716),
            .I(DEBUG_c_3));
    LocalMux I__3097 (
            .O(N__15713),
            .I(DEBUG_c_3));
    LocalMux I__3096 (
            .O(N__15708),
            .I(DEBUG_c_3));
    Odrv4 I__3095 (
            .O(N__15701),
            .I(DEBUG_c_3));
    InMux I__3094 (
            .O(N__15692),
            .I(\receive_module.n3335 ));
    InMux I__3093 (
            .O(N__15689),
            .I(N__15686));
    LocalMux I__3092 (
            .O(N__15686),
            .I(N__15683));
    Span4Mux_h I__3091 (
            .O(N__15683),
            .I(N__15680));
    Odrv4 I__3090 (
            .O(N__15680),
            .I(\receive_module.n123 ));
    InMux I__3089 (
            .O(N__15677),
            .I(N__15673));
    InMux I__3088 (
            .O(N__15676),
            .I(N__15670));
    LocalMux I__3087 (
            .O(N__15673),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    LocalMux I__3086 (
            .O(N__15670),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    InMux I__3085 (
            .O(N__15665),
            .I(bfn_14_13_0_));
    InMux I__3084 (
            .O(N__15662),
            .I(N__15656));
    InMux I__3083 (
            .O(N__15661),
            .I(N__15649));
    InMux I__3082 (
            .O(N__15660),
            .I(N__15649));
    InMux I__3081 (
            .O(N__15659),
            .I(N__15649));
    LocalMux I__3080 (
            .O(N__15656),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__3079 (
            .O(N__15649),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    InMux I__3078 (
            .O(N__15644),
            .I(\transmit_module.video_signal_controller.n3366 ));
    InMux I__3077 (
            .O(N__15641),
            .I(N__15635));
    InMux I__3076 (
            .O(N__15640),
            .I(N__15628));
    InMux I__3075 (
            .O(N__15639),
            .I(N__15628));
    InMux I__3074 (
            .O(N__15638),
            .I(N__15628));
    LocalMux I__3073 (
            .O(N__15635),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__3072 (
            .O(N__15628),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    InMux I__3071 (
            .O(N__15623),
            .I(\transmit_module.video_signal_controller.n3367 ));
    CascadeMux I__3070 (
            .O(N__15620),
            .I(N__15615));
    InMux I__3069 (
            .O(N__15619),
            .I(N__15611));
    InMux I__3068 (
            .O(N__15618),
            .I(N__15604));
    InMux I__3067 (
            .O(N__15615),
            .I(N__15604));
    InMux I__3066 (
            .O(N__15614),
            .I(N__15604));
    LocalMux I__3065 (
            .O(N__15611),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    LocalMux I__3064 (
            .O(N__15604),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    InMux I__3063 (
            .O(N__15599),
            .I(\transmit_module.video_signal_controller.n3368 ));
    CascadeMux I__3062 (
            .O(N__15596),
            .I(N__15592));
    CascadeMux I__3061 (
            .O(N__15595),
            .I(N__15589));
    CascadeBuf I__3060 (
            .O(N__15592),
            .I(N__15586));
    CascadeBuf I__3059 (
            .O(N__15589),
            .I(N__15583));
    CascadeMux I__3058 (
            .O(N__15586),
            .I(N__15580));
    CascadeMux I__3057 (
            .O(N__15583),
            .I(N__15577));
    CascadeBuf I__3056 (
            .O(N__15580),
            .I(N__15574));
    CascadeBuf I__3055 (
            .O(N__15577),
            .I(N__15571));
    CascadeMux I__3054 (
            .O(N__15574),
            .I(N__15568));
    CascadeMux I__3053 (
            .O(N__15571),
            .I(N__15565));
    CascadeBuf I__3052 (
            .O(N__15568),
            .I(N__15562));
    CascadeBuf I__3051 (
            .O(N__15565),
            .I(N__15559));
    CascadeMux I__3050 (
            .O(N__15562),
            .I(N__15556));
    CascadeMux I__3049 (
            .O(N__15559),
            .I(N__15553));
    CascadeBuf I__3048 (
            .O(N__15556),
            .I(N__15550));
    CascadeBuf I__3047 (
            .O(N__15553),
            .I(N__15547));
    CascadeMux I__3046 (
            .O(N__15550),
            .I(N__15544));
    CascadeMux I__3045 (
            .O(N__15547),
            .I(N__15541));
    CascadeBuf I__3044 (
            .O(N__15544),
            .I(N__15538));
    CascadeBuf I__3043 (
            .O(N__15541),
            .I(N__15535));
    CascadeMux I__3042 (
            .O(N__15538),
            .I(N__15532));
    CascadeMux I__3041 (
            .O(N__15535),
            .I(N__15529));
    CascadeBuf I__3040 (
            .O(N__15532),
            .I(N__15526));
    CascadeBuf I__3039 (
            .O(N__15529),
            .I(N__15523));
    CascadeMux I__3038 (
            .O(N__15526),
            .I(N__15520));
    CascadeMux I__3037 (
            .O(N__15523),
            .I(N__15517));
    CascadeBuf I__3036 (
            .O(N__15520),
            .I(N__15514));
    CascadeBuf I__3035 (
            .O(N__15517),
            .I(N__15511));
    CascadeMux I__3034 (
            .O(N__15514),
            .I(N__15508));
    CascadeMux I__3033 (
            .O(N__15511),
            .I(N__15505));
    CascadeBuf I__3032 (
            .O(N__15508),
            .I(N__15502));
    CascadeBuf I__3031 (
            .O(N__15505),
            .I(N__15499));
    CascadeMux I__3030 (
            .O(N__15502),
            .I(N__15496));
    CascadeMux I__3029 (
            .O(N__15499),
            .I(N__15493));
    CascadeBuf I__3028 (
            .O(N__15496),
            .I(N__15490));
    CascadeBuf I__3027 (
            .O(N__15493),
            .I(N__15487));
    CascadeMux I__3026 (
            .O(N__15490),
            .I(N__15484));
    CascadeMux I__3025 (
            .O(N__15487),
            .I(N__15481));
    CascadeBuf I__3024 (
            .O(N__15484),
            .I(N__15478));
    CascadeBuf I__3023 (
            .O(N__15481),
            .I(N__15475));
    CascadeMux I__3022 (
            .O(N__15478),
            .I(N__15472));
    CascadeMux I__3021 (
            .O(N__15475),
            .I(N__15469));
    CascadeBuf I__3020 (
            .O(N__15472),
            .I(N__15466));
    CascadeBuf I__3019 (
            .O(N__15469),
            .I(N__15463));
    CascadeMux I__3018 (
            .O(N__15466),
            .I(N__15460));
    CascadeMux I__3017 (
            .O(N__15463),
            .I(N__15457));
    CascadeBuf I__3016 (
            .O(N__15460),
            .I(N__15454));
    CascadeBuf I__3015 (
            .O(N__15457),
            .I(N__15451));
    CascadeMux I__3014 (
            .O(N__15454),
            .I(N__15448));
    CascadeMux I__3013 (
            .O(N__15451),
            .I(N__15445));
    CascadeBuf I__3012 (
            .O(N__15448),
            .I(N__15442));
    CascadeBuf I__3011 (
            .O(N__15445),
            .I(N__15439));
    CascadeMux I__3010 (
            .O(N__15442),
            .I(N__15436));
    CascadeMux I__3009 (
            .O(N__15439),
            .I(N__15433));
    CascadeBuf I__3008 (
            .O(N__15436),
            .I(N__15430));
    CascadeBuf I__3007 (
            .O(N__15433),
            .I(N__15427));
    CascadeMux I__3006 (
            .O(N__15430),
            .I(N__15424));
    CascadeMux I__3005 (
            .O(N__15427),
            .I(N__15421));
    CascadeBuf I__3004 (
            .O(N__15424),
            .I(N__15418));
    CascadeBuf I__3003 (
            .O(N__15421),
            .I(N__15415));
    CascadeMux I__3002 (
            .O(N__15418),
            .I(N__15412));
    CascadeMux I__3001 (
            .O(N__15415),
            .I(N__15409));
    InMux I__3000 (
            .O(N__15412),
            .I(N__15406));
    InMux I__2999 (
            .O(N__15409),
            .I(N__15403));
    LocalMux I__2998 (
            .O(N__15406),
            .I(N__15400));
    LocalMux I__2997 (
            .O(N__15403),
            .I(N__15397));
    Span4Mux_s2_v I__2996 (
            .O(N__15400),
            .I(N__15394));
    Span4Mux_s1_v I__2995 (
            .O(N__15397),
            .I(N__15391));
    Span4Mux_v I__2994 (
            .O(N__15394),
            .I(N__15388));
    Span4Mux_h I__2993 (
            .O(N__15391),
            .I(N__15384));
    Span4Mux_v I__2992 (
            .O(N__15388),
            .I(N__15381));
    InMux I__2991 (
            .O(N__15387),
            .I(N__15378));
    Sp12to4 I__2990 (
            .O(N__15384),
            .I(N__15374));
    Sp12to4 I__2989 (
            .O(N__15381),
            .I(N__15371));
    LocalMux I__2988 (
            .O(N__15378),
            .I(N__15368));
    InMux I__2987 (
            .O(N__15377),
            .I(N__15365));
    Span12Mux_s10_v I__2986 (
            .O(N__15374),
            .I(N__15360));
    Span12Mux_h I__2985 (
            .O(N__15371),
            .I(N__15360));
    Odrv4 I__2984 (
            .O(N__15368),
            .I(RX_ADDR_2));
    LocalMux I__2983 (
            .O(N__15365),
            .I(RX_ADDR_2));
    Odrv12 I__2982 (
            .O(N__15360),
            .I(RX_ADDR_2));
    InMux I__2981 (
            .O(N__15353),
            .I(N__15350));
    LocalMux I__2980 (
            .O(N__15350),
            .I(N__15347));
    Span4Mux_h I__2979 (
            .O(N__15347),
            .I(N__15344));
    Odrv4 I__2978 (
            .O(N__15344),
            .I(\receive_module.n134 ));
    InMux I__2977 (
            .O(N__15341),
            .I(\receive_module.n3324 ));
    CascadeMux I__2976 (
            .O(N__15338),
            .I(N__15334));
    CascadeMux I__2975 (
            .O(N__15337),
            .I(N__15331));
    CascadeBuf I__2974 (
            .O(N__15334),
            .I(N__15328));
    CascadeBuf I__2973 (
            .O(N__15331),
            .I(N__15325));
    CascadeMux I__2972 (
            .O(N__15328),
            .I(N__15322));
    CascadeMux I__2971 (
            .O(N__15325),
            .I(N__15319));
    CascadeBuf I__2970 (
            .O(N__15322),
            .I(N__15316));
    CascadeBuf I__2969 (
            .O(N__15319),
            .I(N__15313));
    CascadeMux I__2968 (
            .O(N__15316),
            .I(N__15310));
    CascadeMux I__2967 (
            .O(N__15313),
            .I(N__15307));
    CascadeBuf I__2966 (
            .O(N__15310),
            .I(N__15304));
    CascadeBuf I__2965 (
            .O(N__15307),
            .I(N__15301));
    CascadeMux I__2964 (
            .O(N__15304),
            .I(N__15298));
    CascadeMux I__2963 (
            .O(N__15301),
            .I(N__15295));
    CascadeBuf I__2962 (
            .O(N__15298),
            .I(N__15292));
    CascadeBuf I__2961 (
            .O(N__15295),
            .I(N__15289));
    CascadeMux I__2960 (
            .O(N__15292),
            .I(N__15286));
    CascadeMux I__2959 (
            .O(N__15289),
            .I(N__15283));
    CascadeBuf I__2958 (
            .O(N__15286),
            .I(N__15280));
    CascadeBuf I__2957 (
            .O(N__15283),
            .I(N__15277));
    CascadeMux I__2956 (
            .O(N__15280),
            .I(N__15274));
    CascadeMux I__2955 (
            .O(N__15277),
            .I(N__15271));
    CascadeBuf I__2954 (
            .O(N__15274),
            .I(N__15268));
    CascadeBuf I__2953 (
            .O(N__15271),
            .I(N__15265));
    CascadeMux I__2952 (
            .O(N__15268),
            .I(N__15262));
    CascadeMux I__2951 (
            .O(N__15265),
            .I(N__15259));
    CascadeBuf I__2950 (
            .O(N__15262),
            .I(N__15256));
    CascadeBuf I__2949 (
            .O(N__15259),
            .I(N__15253));
    CascadeMux I__2948 (
            .O(N__15256),
            .I(N__15250));
    CascadeMux I__2947 (
            .O(N__15253),
            .I(N__15247));
    CascadeBuf I__2946 (
            .O(N__15250),
            .I(N__15244));
    CascadeBuf I__2945 (
            .O(N__15247),
            .I(N__15241));
    CascadeMux I__2944 (
            .O(N__15244),
            .I(N__15238));
    CascadeMux I__2943 (
            .O(N__15241),
            .I(N__15235));
    CascadeBuf I__2942 (
            .O(N__15238),
            .I(N__15232));
    CascadeBuf I__2941 (
            .O(N__15235),
            .I(N__15229));
    CascadeMux I__2940 (
            .O(N__15232),
            .I(N__15226));
    CascadeMux I__2939 (
            .O(N__15229),
            .I(N__15223));
    CascadeBuf I__2938 (
            .O(N__15226),
            .I(N__15220));
    CascadeBuf I__2937 (
            .O(N__15223),
            .I(N__15217));
    CascadeMux I__2936 (
            .O(N__15220),
            .I(N__15214));
    CascadeMux I__2935 (
            .O(N__15217),
            .I(N__15211));
    CascadeBuf I__2934 (
            .O(N__15214),
            .I(N__15208));
    CascadeBuf I__2933 (
            .O(N__15211),
            .I(N__15205));
    CascadeMux I__2932 (
            .O(N__15208),
            .I(N__15202));
    CascadeMux I__2931 (
            .O(N__15205),
            .I(N__15199));
    CascadeBuf I__2930 (
            .O(N__15202),
            .I(N__15196));
    CascadeBuf I__2929 (
            .O(N__15199),
            .I(N__15193));
    CascadeMux I__2928 (
            .O(N__15196),
            .I(N__15190));
    CascadeMux I__2927 (
            .O(N__15193),
            .I(N__15187));
    CascadeBuf I__2926 (
            .O(N__15190),
            .I(N__15184));
    CascadeBuf I__2925 (
            .O(N__15187),
            .I(N__15181));
    CascadeMux I__2924 (
            .O(N__15184),
            .I(N__15178));
    CascadeMux I__2923 (
            .O(N__15181),
            .I(N__15175));
    CascadeBuf I__2922 (
            .O(N__15178),
            .I(N__15172));
    CascadeBuf I__2921 (
            .O(N__15175),
            .I(N__15169));
    CascadeMux I__2920 (
            .O(N__15172),
            .I(N__15166));
    CascadeMux I__2919 (
            .O(N__15169),
            .I(N__15163));
    CascadeBuf I__2918 (
            .O(N__15166),
            .I(N__15160));
    CascadeBuf I__2917 (
            .O(N__15163),
            .I(N__15157));
    CascadeMux I__2916 (
            .O(N__15160),
            .I(N__15154));
    CascadeMux I__2915 (
            .O(N__15157),
            .I(N__15151));
    InMux I__2914 (
            .O(N__15154),
            .I(N__15148));
    InMux I__2913 (
            .O(N__15151),
            .I(N__15145));
    LocalMux I__2912 (
            .O(N__15148),
            .I(N__15142));
    LocalMux I__2911 (
            .O(N__15145),
            .I(N__15139));
    Span4Mux_s1_v I__2910 (
            .O(N__15142),
            .I(N__15136));
    Span4Mux_s1_v I__2909 (
            .O(N__15139),
            .I(N__15133));
    Span4Mux_v I__2908 (
            .O(N__15136),
            .I(N__15130));
    Span4Mux_h I__2907 (
            .O(N__15133),
            .I(N__15127));
    Span4Mux_v I__2906 (
            .O(N__15130),
            .I(N__15124));
    Span4Mux_h I__2905 (
            .O(N__15127),
            .I(N__15121));
    Sp12to4 I__2904 (
            .O(N__15124),
            .I(N__15117));
    Sp12to4 I__2903 (
            .O(N__15121),
            .I(N__15114));
    InMux I__2902 (
            .O(N__15120),
            .I(N__15110));
    Span12Mux_h I__2901 (
            .O(N__15117),
            .I(N__15105));
    Span12Mux_s9_v I__2900 (
            .O(N__15114),
            .I(N__15105));
    InMux I__2899 (
            .O(N__15113),
            .I(N__15102));
    LocalMux I__2898 (
            .O(N__15110),
            .I(N__15099));
    Span12Mux_v I__2897 (
            .O(N__15105),
            .I(N__15096));
    LocalMux I__2896 (
            .O(N__15102),
            .I(RX_ADDR_3));
    Odrv4 I__2895 (
            .O(N__15099),
            .I(RX_ADDR_3));
    Odrv12 I__2894 (
            .O(N__15096),
            .I(RX_ADDR_3));
    InMux I__2893 (
            .O(N__15089),
            .I(N__15086));
    LocalMux I__2892 (
            .O(N__15086),
            .I(N__15083));
    Odrv12 I__2891 (
            .O(N__15083),
            .I(\receive_module.n133 ));
    InMux I__2890 (
            .O(N__15080),
            .I(\receive_module.n3325 ));
    CascadeMux I__2889 (
            .O(N__15077),
            .I(N__15074));
    CascadeBuf I__2888 (
            .O(N__15074),
            .I(N__15071));
    CascadeMux I__2887 (
            .O(N__15071),
            .I(N__15067));
    CascadeMux I__2886 (
            .O(N__15070),
            .I(N__15064));
    CascadeBuf I__2885 (
            .O(N__15067),
            .I(N__15061));
    CascadeBuf I__2884 (
            .O(N__15064),
            .I(N__15058));
    CascadeMux I__2883 (
            .O(N__15061),
            .I(N__15055));
    CascadeMux I__2882 (
            .O(N__15058),
            .I(N__15052));
    CascadeBuf I__2881 (
            .O(N__15055),
            .I(N__15049));
    CascadeBuf I__2880 (
            .O(N__15052),
            .I(N__15046));
    CascadeMux I__2879 (
            .O(N__15049),
            .I(N__15043));
    CascadeMux I__2878 (
            .O(N__15046),
            .I(N__15040));
    CascadeBuf I__2877 (
            .O(N__15043),
            .I(N__15037));
    CascadeBuf I__2876 (
            .O(N__15040),
            .I(N__15034));
    CascadeMux I__2875 (
            .O(N__15037),
            .I(N__15031));
    CascadeMux I__2874 (
            .O(N__15034),
            .I(N__15028));
    CascadeBuf I__2873 (
            .O(N__15031),
            .I(N__15025));
    CascadeBuf I__2872 (
            .O(N__15028),
            .I(N__15022));
    CascadeMux I__2871 (
            .O(N__15025),
            .I(N__15019));
    CascadeMux I__2870 (
            .O(N__15022),
            .I(N__15016));
    CascadeBuf I__2869 (
            .O(N__15019),
            .I(N__15013));
    CascadeBuf I__2868 (
            .O(N__15016),
            .I(N__15010));
    CascadeMux I__2867 (
            .O(N__15013),
            .I(N__15007));
    CascadeMux I__2866 (
            .O(N__15010),
            .I(N__15004));
    CascadeBuf I__2865 (
            .O(N__15007),
            .I(N__15001));
    CascadeBuf I__2864 (
            .O(N__15004),
            .I(N__14998));
    CascadeMux I__2863 (
            .O(N__15001),
            .I(N__14995));
    CascadeMux I__2862 (
            .O(N__14998),
            .I(N__14992));
    CascadeBuf I__2861 (
            .O(N__14995),
            .I(N__14989));
    CascadeBuf I__2860 (
            .O(N__14992),
            .I(N__14986));
    CascadeMux I__2859 (
            .O(N__14989),
            .I(N__14983));
    CascadeMux I__2858 (
            .O(N__14986),
            .I(N__14980));
    CascadeBuf I__2857 (
            .O(N__14983),
            .I(N__14977));
    CascadeBuf I__2856 (
            .O(N__14980),
            .I(N__14974));
    CascadeMux I__2855 (
            .O(N__14977),
            .I(N__14971));
    CascadeMux I__2854 (
            .O(N__14974),
            .I(N__14968));
    CascadeBuf I__2853 (
            .O(N__14971),
            .I(N__14965));
    CascadeBuf I__2852 (
            .O(N__14968),
            .I(N__14962));
    CascadeMux I__2851 (
            .O(N__14965),
            .I(N__14959));
    CascadeMux I__2850 (
            .O(N__14962),
            .I(N__14956));
    CascadeBuf I__2849 (
            .O(N__14959),
            .I(N__14953));
    CascadeBuf I__2848 (
            .O(N__14956),
            .I(N__14950));
    CascadeMux I__2847 (
            .O(N__14953),
            .I(N__14947));
    CascadeMux I__2846 (
            .O(N__14950),
            .I(N__14944));
    CascadeBuf I__2845 (
            .O(N__14947),
            .I(N__14941));
    CascadeBuf I__2844 (
            .O(N__14944),
            .I(N__14938));
    CascadeMux I__2843 (
            .O(N__14941),
            .I(N__14935));
    CascadeMux I__2842 (
            .O(N__14938),
            .I(N__14932));
    CascadeBuf I__2841 (
            .O(N__14935),
            .I(N__14929));
    CascadeBuf I__2840 (
            .O(N__14932),
            .I(N__14926));
    CascadeMux I__2839 (
            .O(N__14929),
            .I(N__14923));
    CascadeMux I__2838 (
            .O(N__14926),
            .I(N__14920));
    CascadeBuf I__2837 (
            .O(N__14923),
            .I(N__14917));
    CascadeBuf I__2836 (
            .O(N__14920),
            .I(N__14914));
    CascadeMux I__2835 (
            .O(N__14917),
            .I(N__14911));
    CascadeMux I__2834 (
            .O(N__14914),
            .I(N__14908));
    CascadeBuf I__2833 (
            .O(N__14911),
            .I(N__14905));
    CascadeBuf I__2832 (
            .O(N__14908),
            .I(N__14902));
    CascadeMux I__2831 (
            .O(N__14905),
            .I(N__14899));
    CascadeMux I__2830 (
            .O(N__14902),
            .I(N__14896));
    InMux I__2829 (
            .O(N__14899),
            .I(N__14893));
    CascadeBuf I__2828 (
            .O(N__14896),
            .I(N__14890));
    LocalMux I__2827 (
            .O(N__14893),
            .I(N__14887));
    CascadeMux I__2826 (
            .O(N__14890),
            .I(N__14884));
    Span4Mux_s1_v I__2825 (
            .O(N__14887),
            .I(N__14881));
    InMux I__2824 (
            .O(N__14884),
            .I(N__14878));
    Span4Mux_h I__2823 (
            .O(N__14881),
            .I(N__14875));
    LocalMux I__2822 (
            .O(N__14878),
            .I(N__14872));
    Sp12to4 I__2821 (
            .O(N__14875),
            .I(N__14867));
    Span12Mux_s10_v I__2820 (
            .O(N__14872),
            .I(N__14864));
    InMux I__2819 (
            .O(N__14871),
            .I(N__14861));
    InMux I__2818 (
            .O(N__14870),
            .I(N__14858));
    Span12Mux_s10_v I__2817 (
            .O(N__14867),
            .I(N__14853));
    Span12Mux_h I__2816 (
            .O(N__14864),
            .I(N__14853));
    LocalMux I__2815 (
            .O(N__14861),
            .I(RX_ADDR_4));
    LocalMux I__2814 (
            .O(N__14858),
            .I(RX_ADDR_4));
    Odrv12 I__2813 (
            .O(N__14853),
            .I(RX_ADDR_4));
    CascadeMux I__2812 (
            .O(N__14846),
            .I(N__14843));
    InMux I__2811 (
            .O(N__14843),
            .I(N__14840));
    LocalMux I__2810 (
            .O(N__14840),
            .I(\receive_module.n132 ));
    InMux I__2809 (
            .O(N__14837),
            .I(\receive_module.n3326 ));
    CascadeMux I__2808 (
            .O(N__14834),
            .I(N__14831));
    CascadeBuf I__2807 (
            .O(N__14831),
            .I(N__14828));
    CascadeMux I__2806 (
            .O(N__14828),
            .I(N__14824));
    CascadeMux I__2805 (
            .O(N__14827),
            .I(N__14821));
    CascadeBuf I__2804 (
            .O(N__14824),
            .I(N__14818));
    CascadeBuf I__2803 (
            .O(N__14821),
            .I(N__14815));
    CascadeMux I__2802 (
            .O(N__14818),
            .I(N__14812));
    CascadeMux I__2801 (
            .O(N__14815),
            .I(N__14809));
    CascadeBuf I__2800 (
            .O(N__14812),
            .I(N__14806));
    CascadeBuf I__2799 (
            .O(N__14809),
            .I(N__14803));
    CascadeMux I__2798 (
            .O(N__14806),
            .I(N__14800));
    CascadeMux I__2797 (
            .O(N__14803),
            .I(N__14797));
    CascadeBuf I__2796 (
            .O(N__14800),
            .I(N__14794));
    CascadeBuf I__2795 (
            .O(N__14797),
            .I(N__14791));
    CascadeMux I__2794 (
            .O(N__14794),
            .I(N__14788));
    CascadeMux I__2793 (
            .O(N__14791),
            .I(N__14785));
    CascadeBuf I__2792 (
            .O(N__14788),
            .I(N__14782));
    CascadeBuf I__2791 (
            .O(N__14785),
            .I(N__14779));
    CascadeMux I__2790 (
            .O(N__14782),
            .I(N__14776));
    CascadeMux I__2789 (
            .O(N__14779),
            .I(N__14773));
    CascadeBuf I__2788 (
            .O(N__14776),
            .I(N__14770));
    CascadeBuf I__2787 (
            .O(N__14773),
            .I(N__14767));
    CascadeMux I__2786 (
            .O(N__14770),
            .I(N__14764));
    CascadeMux I__2785 (
            .O(N__14767),
            .I(N__14761));
    CascadeBuf I__2784 (
            .O(N__14764),
            .I(N__14758));
    CascadeBuf I__2783 (
            .O(N__14761),
            .I(N__14755));
    CascadeMux I__2782 (
            .O(N__14758),
            .I(N__14752));
    CascadeMux I__2781 (
            .O(N__14755),
            .I(N__14749));
    CascadeBuf I__2780 (
            .O(N__14752),
            .I(N__14746));
    CascadeBuf I__2779 (
            .O(N__14749),
            .I(N__14743));
    CascadeMux I__2778 (
            .O(N__14746),
            .I(N__14740));
    CascadeMux I__2777 (
            .O(N__14743),
            .I(N__14737));
    CascadeBuf I__2776 (
            .O(N__14740),
            .I(N__14734));
    CascadeBuf I__2775 (
            .O(N__14737),
            .I(N__14731));
    CascadeMux I__2774 (
            .O(N__14734),
            .I(N__14728));
    CascadeMux I__2773 (
            .O(N__14731),
            .I(N__14725));
    CascadeBuf I__2772 (
            .O(N__14728),
            .I(N__14722));
    CascadeBuf I__2771 (
            .O(N__14725),
            .I(N__14719));
    CascadeMux I__2770 (
            .O(N__14722),
            .I(N__14716));
    CascadeMux I__2769 (
            .O(N__14719),
            .I(N__14713));
    CascadeBuf I__2768 (
            .O(N__14716),
            .I(N__14710));
    CascadeBuf I__2767 (
            .O(N__14713),
            .I(N__14707));
    CascadeMux I__2766 (
            .O(N__14710),
            .I(N__14704));
    CascadeMux I__2765 (
            .O(N__14707),
            .I(N__14701));
    CascadeBuf I__2764 (
            .O(N__14704),
            .I(N__14698));
    CascadeBuf I__2763 (
            .O(N__14701),
            .I(N__14695));
    CascadeMux I__2762 (
            .O(N__14698),
            .I(N__14692));
    CascadeMux I__2761 (
            .O(N__14695),
            .I(N__14689));
    CascadeBuf I__2760 (
            .O(N__14692),
            .I(N__14686));
    CascadeBuf I__2759 (
            .O(N__14689),
            .I(N__14683));
    CascadeMux I__2758 (
            .O(N__14686),
            .I(N__14680));
    CascadeMux I__2757 (
            .O(N__14683),
            .I(N__14677));
    CascadeBuf I__2756 (
            .O(N__14680),
            .I(N__14674));
    CascadeBuf I__2755 (
            .O(N__14677),
            .I(N__14671));
    CascadeMux I__2754 (
            .O(N__14674),
            .I(N__14668));
    CascadeMux I__2753 (
            .O(N__14671),
            .I(N__14665));
    CascadeBuf I__2752 (
            .O(N__14668),
            .I(N__14662));
    CascadeBuf I__2751 (
            .O(N__14665),
            .I(N__14659));
    CascadeMux I__2750 (
            .O(N__14662),
            .I(N__14656));
    CascadeMux I__2749 (
            .O(N__14659),
            .I(N__14653));
    InMux I__2748 (
            .O(N__14656),
            .I(N__14650));
    CascadeBuf I__2747 (
            .O(N__14653),
            .I(N__14647));
    LocalMux I__2746 (
            .O(N__14650),
            .I(N__14644));
    CascadeMux I__2745 (
            .O(N__14647),
            .I(N__14641));
    Span4Mux_s2_v I__2744 (
            .O(N__14644),
            .I(N__14638));
    InMux I__2743 (
            .O(N__14641),
            .I(N__14635));
    Span4Mux_h I__2742 (
            .O(N__14638),
            .I(N__14632));
    LocalMux I__2741 (
            .O(N__14635),
            .I(N__14629));
    Span4Mux_h I__2740 (
            .O(N__14632),
            .I(N__14626));
    Span4Mux_s2_v I__2739 (
            .O(N__14629),
            .I(N__14623));
    Span4Mux_h I__2738 (
            .O(N__14626),
            .I(N__14618));
    Span4Mux_h I__2737 (
            .O(N__14623),
            .I(N__14618));
    Span4Mux_v I__2736 (
            .O(N__14618),
            .I(N__14615));
    Span4Mux_v I__2735 (
            .O(N__14615),
            .I(N__14612));
    Span4Mux_v I__2734 (
            .O(N__14612),
            .I(N__14607));
    InMux I__2733 (
            .O(N__14611),
            .I(N__14604));
    InMux I__2732 (
            .O(N__14610),
            .I(N__14601));
    Span4Mux_v I__2731 (
            .O(N__14607),
            .I(N__14598));
    LocalMux I__2730 (
            .O(N__14604),
            .I(RX_ADDR_5));
    LocalMux I__2729 (
            .O(N__14601),
            .I(RX_ADDR_5));
    Odrv4 I__2728 (
            .O(N__14598),
            .I(RX_ADDR_5));
    InMux I__2727 (
            .O(N__14591),
            .I(N__14588));
    LocalMux I__2726 (
            .O(N__14588),
            .I(\receive_module.n131 ));
    InMux I__2725 (
            .O(N__14585),
            .I(\receive_module.n3327 ));
    CascadeMux I__2724 (
            .O(N__14582),
            .I(N__14578));
    CascadeMux I__2723 (
            .O(N__14581),
            .I(N__14575));
    CascadeBuf I__2722 (
            .O(N__14578),
            .I(N__14572));
    CascadeBuf I__2721 (
            .O(N__14575),
            .I(N__14569));
    CascadeMux I__2720 (
            .O(N__14572),
            .I(N__14566));
    CascadeMux I__2719 (
            .O(N__14569),
            .I(N__14563));
    CascadeBuf I__2718 (
            .O(N__14566),
            .I(N__14560));
    CascadeBuf I__2717 (
            .O(N__14563),
            .I(N__14557));
    CascadeMux I__2716 (
            .O(N__14560),
            .I(N__14554));
    CascadeMux I__2715 (
            .O(N__14557),
            .I(N__14551));
    CascadeBuf I__2714 (
            .O(N__14554),
            .I(N__14548));
    CascadeBuf I__2713 (
            .O(N__14551),
            .I(N__14545));
    CascadeMux I__2712 (
            .O(N__14548),
            .I(N__14542));
    CascadeMux I__2711 (
            .O(N__14545),
            .I(N__14539));
    CascadeBuf I__2710 (
            .O(N__14542),
            .I(N__14536));
    CascadeBuf I__2709 (
            .O(N__14539),
            .I(N__14533));
    CascadeMux I__2708 (
            .O(N__14536),
            .I(N__14530));
    CascadeMux I__2707 (
            .O(N__14533),
            .I(N__14527));
    CascadeBuf I__2706 (
            .O(N__14530),
            .I(N__14524));
    CascadeBuf I__2705 (
            .O(N__14527),
            .I(N__14521));
    CascadeMux I__2704 (
            .O(N__14524),
            .I(N__14518));
    CascadeMux I__2703 (
            .O(N__14521),
            .I(N__14515));
    CascadeBuf I__2702 (
            .O(N__14518),
            .I(N__14512));
    CascadeBuf I__2701 (
            .O(N__14515),
            .I(N__14509));
    CascadeMux I__2700 (
            .O(N__14512),
            .I(N__14506));
    CascadeMux I__2699 (
            .O(N__14509),
            .I(N__14503));
    CascadeBuf I__2698 (
            .O(N__14506),
            .I(N__14500));
    CascadeBuf I__2697 (
            .O(N__14503),
            .I(N__14497));
    CascadeMux I__2696 (
            .O(N__14500),
            .I(N__14494));
    CascadeMux I__2695 (
            .O(N__14497),
            .I(N__14491));
    CascadeBuf I__2694 (
            .O(N__14494),
            .I(N__14488));
    CascadeBuf I__2693 (
            .O(N__14491),
            .I(N__14485));
    CascadeMux I__2692 (
            .O(N__14488),
            .I(N__14482));
    CascadeMux I__2691 (
            .O(N__14485),
            .I(N__14479));
    CascadeBuf I__2690 (
            .O(N__14482),
            .I(N__14476));
    CascadeBuf I__2689 (
            .O(N__14479),
            .I(N__14473));
    CascadeMux I__2688 (
            .O(N__14476),
            .I(N__14470));
    CascadeMux I__2687 (
            .O(N__14473),
            .I(N__14467));
    CascadeBuf I__2686 (
            .O(N__14470),
            .I(N__14464));
    CascadeBuf I__2685 (
            .O(N__14467),
            .I(N__14461));
    CascadeMux I__2684 (
            .O(N__14464),
            .I(N__14458));
    CascadeMux I__2683 (
            .O(N__14461),
            .I(N__14455));
    CascadeBuf I__2682 (
            .O(N__14458),
            .I(N__14452));
    CascadeBuf I__2681 (
            .O(N__14455),
            .I(N__14449));
    CascadeMux I__2680 (
            .O(N__14452),
            .I(N__14446));
    CascadeMux I__2679 (
            .O(N__14449),
            .I(N__14443));
    CascadeBuf I__2678 (
            .O(N__14446),
            .I(N__14440));
    CascadeBuf I__2677 (
            .O(N__14443),
            .I(N__14437));
    CascadeMux I__2676 (
            .O(N__14440),
            .I(N__14434));
    CascadeMux I__2675 (
            .O(N__14437),
            .I(N__14431));
    CascadeBuf I__2674 (
            .O(N__14434),
            .I(N__14428));
    CascadeBuf I__2673 (
            .O(N__14431),
            .I(N__14425));
    CascadeMux I__2672 (
            .O(N__14428),
            .I(N__14422));
    CascadeMux I__2671 (
            .O(N__14425),
            .I(N__14419));
    CascadeBuf I__2670 (
            .O(N__14422),
            .I(N__14416));
    CascadeBuf I__2669 (
            .O(N__14419),
            .I(N__14413));
    CascadeMux I__2668 (
            .O(N__14416),
            .I(N__14410));
    CascadeMux I__2667 (
            .O(N__14413),
            .I(N__14407));
    CascadeBuf I__2666 (
            .O(N__14410),
            .I(N__14404));
    CascadeBuf I__2665 (
            .O(N__14407),
            .I(N__14401));
    CascadeMux I__2664 (
            .O(N__14404),
            .I(N__14398));
    CascadeMux I__2663 (
            .O(N__14401),
            .I(N__14395));
    InMux I__2662 (
            .O(N__14398),
            .I(N__14392));
    InMux I__2661 (
            .O(N__14395),
            .I(N__14389));
    LocalMux I__2660 (
            .O(N__14392),
            .I(N__14386));
    LocalMux I__2659 (
            .O(N__14389),
            .I(N__14383));
    Span12Mux_h I__2658 (
            .O(N__14386),
            .I(N__14378));
    Span12Mux_v I__2657 (
            .O(N__14383),
            .I(N__14375));
    InMux I__2656 (
            .O(N__14382),
            .I(N__14372));
    InMux I__2655 (
            .O(N__14381),
            .I(N__14369));
    Span12Mux_v I__2654 (
            .O(N__14378),
            .I(N__14364));
    Span12Mux_h I__2653 (
            .O(N__14375),
            .I(N__14364));
    LocalMux I__2652 (
            .O(N__14372),
            .I(RX_ADDR_6));
    LocalMux I__2651 (
            .O(N__14369),
            .I(RX_ADDR_6));
    Odrv12 I__2650 (
            .O(N__14364),
            .I(RX_ADDR_6));
    CascadeMux I__2649 (
            .O(N__14357),
            .I(N__14354));
    InMux I__2648 (
            .O(N__14354),
            .I(N__14351));
    LocalMux I__2647 (
            .O(N__14351),
            .I(\receive_module.n130 ));
    InMux I__2646 (
            .O(N__14348),
            .I(\receive_module.n3328 ));
    CascadeMux I__2645 (
            .O(N__14345),
            .I(N__14341));
    CascadeMux I__2644 (
            .O(N__14344),
            .I(N__14338));
    CascadeBuf I__2643 (
            .O(N__14341),
            .I(N__14335));
    CascadeBuf I__2642 (
            .O(N__14338),
            .I(N__14332));
    CascadeMux I__2641 (
            .O(N__14335),
            .I(N__14329));
    CascadeMux I__2640 (
            .O(N__14332),
            .I(N__14326));
    CascadeBuf I__2639 (
            .O(N__14329),
            .I(N__14323));
    CascadeBuf I__2638 (
            .O(N__14326),
            .I(N__14320));
    CascadeMux I__2637 (
            .O(N__14323),
            .I(N__14317));
    CascadeMux I__2636 (
            .O(N__14320),
            .I(N__14314));
    CascadeBuf I__2635 (
            .O(N__14317),
            .I(N__14311));
    CascadeBuf I__2634 (
            .O(N__14314),
            .I(N__14308));
    CascadeMux I__2633 (
            .O(N__14311),
            .I(N__14305));
    CascadeMux I__2632 (
            .O(N__14308),
            .I(N__14302));
    CascadeBuf I__2631 (
            .O(N__14305),
            .I(N__14299));
    CascadeBuf I__2630 (
            .O(N__14302),
            .I(N__14296));
    CascadeMux I__2629 (
            .O(N__14299),
            .I(N__14293));
    CascadeMux I__2628 (
            .O(N__14296),
            .I(N__14290));
    CascadeBuf I__2627 (
            .O(N__14293),
            .I(N__14287));
    CascadeBuf I__2626 (
            .O(N__14290),
            .I(N__14284));
    CascadeMux I__2625 (
            .O(N__14287),
            .I(N__14281));
    CascadeMux I__2624 (
            .O(N__14284),
            .I(N__14278));
    CascadeBuf I__2623 (
            .O(N__14281),
            .I(N__14275));
    CascadeBuf I__2622 (
            .O(N__14278),
            .I(N__14272));
    CascadeMux I__2621 (
            .O(N__14275),
            .I(N__14269));
    CascadeMux I__2620 (
            .O(N__14272),
            .I(N__14266));
    CascadeBuf I__2619 (
            .O(N__14269),
            .I(N__14263));
    CascadeBuf I__2618 (
            .O(N__14266),
            .I(N__14260));
    CascadeMux I__2617 (
            .O(N__14263),
            .I(N__14257));
    CascadeMux I__2616 (
            .O(N__14260),
            .I(N__14254));
    CascadeBuf I__2615 (
            .O(N__14257),
            .I(N__14251));
    CascadeBuf I__2614 (
            .O(N__14254),
            .I(N__14248));
    CascadeMux I__2613 (
            .O(N__14251),
            .I(N__14245));
    CascadeMux I__2612 (
            .O(N__14248),
            .I(N__14242));
    CascadeBuf I__2611 (
            .O(N__14245),
            .I(N__14239));
    CascadeBuf I__2610 (
            .O(N__14242),
            .I(N__14236));
    CascadeMux I__2609 (
            .O(N__14239),
            .I(N__14233));
    CascadeMux I__2608 (
            .O(N__14236),
            .I(N__14230));
    CascadeBuf I__2607 (
            .O(N__14233),
            .I(N__14227));
    CascadeBuf I__2606 (
            .O(N__14230),
            .I(N__14224));
    CascadeMux I__2605 (
            .O(N__14227),
            .I(N__14221));
    CascadeMux I__2604 (
            .O(N__14224),
            .I(N__14218));
    CascadeBuf I__2603 (
            .O(N__14221),
            .I(N__14215));
    CascadeBuf I__2602 (
            .O(N__14218),
            .I(N__14212));
    CascadeMux I__2601 (
            .O(N__14215),
            .I(N__14209));
    CascadeMux I__2600 (
            .O(N__14212),
            .I(N__14206));
    CascadeBuf I__2599 (
            .O(N__14209),
            .I(N__14203));
    CascadeBuf I__2598 (
            .O(N__14206),
            .I(N__14200));
    CascadeMux I__2597 (
            .O(N__14203),
            .I(N__14197));
    CascadeMux I__2596 (
            .O(N__14200),
            .I(N__14194));
    CascadeBuf I__2595 (
            .O(N__14197),
            .I(N__14191));
    CascadeBuf I__2594 (
            .O(N__14194),
            .I(N__14188));
    CascadeMux I__2593 (
            .O(N__14191),
            .I(N__14185));
    CascadeMux I__2592 (
            .O(N__14188),
            .I(N__14182));
    CascadeBuf I__2591 (
            .O(N__14185),
            .I(N__14179));
    CascadeBuf I__2590 (
            .O(N__14182),
            .I(N__14176));
    CascadeMux I__2589 (
            .O(N__14179),
            .I(N__14173));
    CascadeMux I__2588 (
            .O(N__14176),
            .I(N__14170));
    CascadeBuf I__2587 (
            .O(N__14173),
            .I(N__14167));
    CascadeBuf I__2586 (
            .O(N__14170),
            .I(N__14164));
    CascadeMux I__2585 (
            .O(N__14167),
            .I(N__14161));
    CascadeMux I__2584 (
            .O(N__14164),
            .I(N__14158));
    InMux I__2583 (
            .O(N__14161),
            .I(N__14155));
    InMux I__2582 (
            .O(N__14158),
            .I(N__14152));
    LocalMux I__2581 (
            .O(N__14155),
            .I(N__14149));
    LocalMux I__2580 (
            .O(N__14152),
            .I(N__14146));
    Span4Mux_s1_v I__2579 (
            .O(N__14149),
            .I(N__14143));
    Span4Mux_s1_v I__2578 (
            .O(N__14146),
            .I(N__14140));
    Span4Mux_h I__2577 (
            .O(N__14143),
            .I(N__14137));
    Sp12to4 I__2576 (
            .O(N__14140),
            .I(N__14134));
    Sp12to4 I__2575 (
            .O(N__14137),
            .I(N__14131));
    Span12Mux_s9_v I__2574 (
            .O(N__14134),
            .I(N__14126));
    Span12Mux_s9_v I__2573 (
            .O(N__14131),
            .I(N__14123));
    InMux I__2572 (
            .O(N__14130),
            .I(N__14120));
    InMux I__2571 (
            .O(N__14129),
            .I(N__14117));
    Span12Mux_v I__2570 (
            .O(N__14126),
            .I(N__14112));
    Span12Mux_v I__2569 (
            .O(N__14123),
            .I(N__14112));
    LocalMux I__2568 (
            .O(N__14120),
            .I(RX_ADDR_7));
    LocalMux I__2567 (
            .O(N__14117),
            .I(RX_ADDR_7));
    Odrv12 I__2566 (
            .O(N__14112),
            .I(RX_ADDR_7));
    InMux I__2565 (
            .O(N__14105),
            .I(N__14102));
    LocalMux I__2564 (
            .O(N__14102),
            .I(\receive_module.n129 ));
    InMux I__2563 (
            .O(N__14099),
            .I(\receive_module.n3329 ));
    CascadeMux I__2562 (
            .O(N__14096),
            .I(N__14093));
    CascadeBuf I__2561 (
            .O(N__14093),
            .I(N__14089));
    CascadeMux I__2560 (
            .O(N__14092),
            .I(N__14086));
    CascadeMux I__2559 (
            .O(N__14089),
            .I(N__14083));
    CascadeBuf I__2558 (
            .O(N__14086),
            .I(N__14080));
    CascadeBuf I__2557 (
            .O(N__14083),
            .I(N__14077));
    CascadeMux I__2556 (
            .O(N__14080),
            .I(N__14074));
    CascadeMux I__2555 (
            .O(N__14077),
            .I(N__14071));
    CascadeBuf I__2554 (
            .O(N__14074),
            .I(N__14068));
    CascadeBuf I__2553 (
            .O(N__14071),
            .I(N__14065));
    CascadeMux I__2552 (
            .O(N__14068),
            .I(N__14062));
    CascadeMux I__2551 (
            .O(N__14065),
            .I(N__14059));
    CascadeBuf I__2550 (
            .O(N__14062),
            .I(N__14056));
    CascadeBuf I__2549 (
            .O(N__14059),
            .I(N__14053));
    CascadeMux I__2548 (
            .O(N__14056),
            .I(N__14050));
    CascadeMux I__2547 (
            .O(N__14053),
            .I(N__14047));
    CascadeBuf I__2546 (
            .O(N__14050),
            .I(N__14044));
    CascadeBuf I__2545 (
            .O(N__14047),
            .I(N__14041));
    CascadeMux I__2544 (
            .O(N__14044),
            .I(N__14038));
    CascadeMux I__2543 (
            .O(N__14041),
            .I(N__14035));
    CascadeBuf I__2542 (
            .O(N__14038),
            .I(N__14032));
    CascadeBuf I__2541 (
            .O(N__14035),
            .I(N__14029));
    CascadeMux I__2540 (
            .O(N__14032),
            .I(N__14026));
    CascadeMux I__2539 (
            .O(N__14029),
            .I(N__14023));
    CascadeBuf I__2538 (
            .O(N__14026),
            .I(N__14020));
    CascadeBuf I__2537 (
            .O(N__14023),
            .I(N__14017));
    CascadeMux I__2536 (
            .O(N__14020),
            .I(N__14014));
    CascadeMux I__2535 (
            .O(N__14017),
            .I(N__14011));
    CascadeBuf I__2534 (
            .O(N__14014),
            .I(N__14008));
    CascadeBuf I__2533 (
            .O(N__14011),
            .I(N__14005));
    CascadeMux I__2532 (
            .O(N__14008),
            .I(N__14002));
    CascadeMux I__2531 (
            .O(N__14005),
            .I(N__13999));
    CascadeBuf I__2530 (
            .O(N__14002),
            .I(N__13996));
    CascadeBuf I__2529 (
            .O(N__13999),
            .I(N__13993));
    CascadeMux I__2528 (
            .O(N__13996),
            .I(N__13990));
    CascadeMux I__2527 (
            .O(N__13993),
            .I(N__13987));
    CascadeBuf I__2526 (
            .O(N__13990),
            .I(N__13984));
    CascadeBuf I__2525 (
            .O(N__13987),
            .I(N__13981));
    CascadeMux I__2524 (
            .O(N__13984),
            .I(N__13978));
    CascadeMux I__2523 (
            .O(N__13981),
            .I(N__13975));
    CascadeBuf I__2522 (
            .O(N__13978),
            .I(N__13972));
    CascadeBuf I__2521 (
            .O(N__13975),
            .I(N__13969));
    CascadeMux I__2520 (
            .O(N__13972),
            .I(N__13966));
    CascadeMux I__2519 (
            .O(N__13969),
            .I(N__13963));
    CascadeBuf I__2518 (
            .O(N__13966),
            .I(N__13960));
    CascadeBuf I__2517 (
            .O(N__13963),
            .I(N__13957));
    CascadeMux I__2516 (
            .O(N__13960),
            .I(N__13954));
    CascadeMux I__2515 (
            .O(N__13957),
            .I(N__13951));
    CascadeBuf I__2514 (
            .O(N__13954),
            .I(N__13948));
    CascadeBuf I__2513 (
            .O(N__13951),
            .I(N__13945));
    CascadeMux I__2512 (
            .O(N__13948),
            .I(N__13942));
    CascadeMux I__2511 (
            .O(N__13945),
            .I(N__13939));
    CascadeBuf I__2510 (
            .O(N__13942),
            .I(N__13936));
    CascadeBuf I__2509 (
            .O(N__13939),
            .I(N__13933));
    CascadeMux I__2508 (
            .O(N__13936),
            .I(N__13930));
    CascadeMux I__2507 (
            .O(N__13933),
            .I(N__13927));
    CascadeBuf I__2506 (
            .O(N__13930),
            .I(N__13924));
    CascadeBuf I__2505 (
            .O(N__13927),
            .I(N__13921));
    CascadeMux I__2504 (
            .O(N__13924),
            .I(N__13918));
    CascadeMux I__2503 (
            .O(N__13921),
            .I(N__13915));
    CascadeBuf I__2502 (
            .O(N__13918),
            .I(N__13912));
    InMux I__2501 (
            .O(N__13915),
            .I(N__13909));
    CascadeMux I__2500 (
            .O(N__13912),
            .I(N__13906));
    LocalMux I__2499 (
            .O(N__13909),
            .I(N__13903));
    InMux I__2498 (
            .O(N__13906),
            .I(N__13900));
    Span4Mux_s2_v I__2497 (
            .O(N__13903),
            .I(N__13896));
    LocalMux I__2496 (
            .O(N__13900),
            .I(N__13893));
    InMux I__2495 (
            .O(N__13899),
            .I(N__13890));
    Sp12to4 I__2494 (
            .O(N__13896),
            .I(N__13887));
    Span12Mux_s9_v I__2493 (
            .O(N__13893),
            .I(N__13884));
    LocalMux I__2492 (
            .O(N__13890),
            .I(N__13881));
    Span12Mux_s9_v I__2491 (
            .O(N__13887),
            .I(N__13877));
    Span12Mux_v I__2490 (
            .O(N__13884),
            .I(N__13874));
    Span4Mux_h I__2489 (
            .O(N__13881),
            .I(N__13871));
    InMux I__2488 (
            .O(N__13880),
            .I(N__13868));
    Span12Mux_v I__2487 (
            .O(N__13877),
            .I(N__13865));
    Span12Mux_h I__2486 (
            .O(N__13874),
            .I(N__13862));
    Odrv4 I__2485 (
            .O(N__13871),
            .I(RX_ADDR_8));
    LocalMux I__2484 (
            .O(N__13868),
            .I(RX_ADDR_8));
    Odrv12 I__2483 (
            .O(N__13865),
            .I(RX_ADDR_8));
    Odrv12 I__2482 (
            .O(N__13862),
            .I(RX_ADDR_8));
    InMux I__2481 (
            .O(N__13853),
            .I(N__13850));
    LocalMux I__2480 (
            .O(N__13850),
            .I(N__13847));
    Span4Mux_v I__2479 (
            .O(N__13847),
            .I(N__13844));
    Odrv4 I__2478 (
            .O(N__13844),
            .I(\receive_module.n128 ));
    InMux I__2477 (
            .O(N__13841),
            .I(bfn_14_12_0_));
    CascadeMux I__2476 (
            .O(N__13838),
            .I(N__13834));
    CascadeMux I__2475 (
            .O(N__13837),
            .I(N__13831));
    CascadeBuf I__2474 (
            .O(N__13834),
            .I(N__13828));
    CascadeBuf I__2473 (
            .O(N__13831),
            .I(N__13825));
    CascadeMux I__2472 (
            .O(N__13828),
            .I(N__13822));
    CascadeMux I__2471 (
            .O(N__13825),
            .I(N__13819));
    CascadeBuf I__2470 (
            .O(N__13822),
            .I(N__13816));
    CascadeBuf I__2469 (
            .O(N__13819),
            .I(N__13813));
    CascadeMux I__2468 (
            .O(N__13816),
            .I(N__13810));
    CascadeMux I__2467 (
            .O(N__13813),
            .I(N__13807));
    CascadeBuf I__2466 (
            .O(N__13810),
            .I(N__13804));
    CascadeBuf I__2465 (
            .O(N__13807),
            .I(N__13801));
    CascadeMux I__2464 (
            .O(N__13804),
            .I(N__13798));
    CascadeMux I__2463 (
            .O(N__13801),
            .I(N__13795));
    CascadeBuf I__2462 (
            .O(N__13798),
            .I(N__13792));
    CascadeBuf I__2461 (
            .O(N__13795),
            .I(N__13789));
    CascadeMux I__2460 (
            .O(N__13792),
            .I(N__13786));
    CascadeMux I__2459 (
            .O(N__13789),
            .I(N__13783));
    CascadeBuf I__2458 (
            .O(N__13786),
            .I(N__13780));
    CascadeBuf I__2457 (
            .O(N__13783),
            .I(N__13777));
    CascadeMux I__2456 (
            .O(N__13780),
            .I(N__13774));
    CascadeMux I__2455 (
            .O(N__13777),
            .I(N__13771));
    CascadeBuf I__2454 (
            .O(N__13774),
            .I(N__13768));
    CascadeBuf I__2453 (
            .O(N__13771),
            .I(N__13765));
    CascadeMux I__2452 (
            .O(N__13768),
            .I(N__13762));
    CascadeMux I__2451 (
            .O(N__13765),
            .I(N__13759));
    CascadeBuf I__2450 (
            .O(N__13762),
            .I(N__13756));
    CascadeBuf I__2449 (
            .O(N__13759),
            .I(N__13753));
    CascadeMux I__2448 (
            .O(N__13756),
            .I(N__13750));
    CascadeMux I__2447 (
            .O(N__13753),
            .I(N__13747));
    CascadeBuf I__2446 (
            .O(N__13750),
            .I(N__13744));
    CascadeBuf I__2445 (
            .O(N__13747),
            .I(N__13741));
    CascadeMux I__2444 (
            .O(N__13744),
            .I(N__13738));
    CascadeMux I__2443 (
            .O(N__13741),
            .I(N__13735));
    CascadeBuf I__2442 (
            .O(N__13738),
            .I(N__13732));
    CascadeBuf I__2441 (
            .O(N__13735),
            .I(N__13729));
    CascadeMux I__2440 (
            .O(N__13732),
            .I(N__13726));
    CascadeMux I__2439 (
            .O(N__13729),
            .I(N__13723));
    CascadeBuf I__2438 (
            .O(N__13726),
            .I(N__13720));
    CascadeBuf I__2437 (
            .O(N__13723),
            .I(N__13717));
    CascadeMux I__2436 (
            .O(N__13720),
            .I(N__13714));
    CascadeMux I__2435 (
            .O(N__13717),
            .I(N__13711));
    CascadeBuf I__2434 (
            .O(N__13714),
            .I(N__13708));
    CascadeBuf I__2433 (
            .O(N__13711),
            .I(N__13705));
    CascadeMux I__2432 (
            .O(N__13708),
            .I(N__13702));
    CascadeMux I__2431 (
            .O(N__13705),
            .I(N__13699));
    CascadeBuf I__2430 (
            .O(N__13702),
            .I(N__13696));
    CascadeBuf I__2429 (
            .O(N__13699),
            .I(N__13693));
    CascadeMux I__2428 (
            .O(N__13696),
            .I(N__13690));
    CascadeMux I__2427 (
            .O(N__13693),
            .I(N__13687));
    CascadeBuf I__2426 (
            .O(N__13690),
            .I(N__13684));
    CascadeBuf I__2425 (
            .O(N__13687),
            .I(N__13681));
    CascadeMux I__2424 (
            .O(N__13684),
            .I(N__13678));
    CascadeMux I__2423 (
            .O(N__13681),
            .I(N__13675));
    CascadeBuf I__2422 (
            .O(N__13678),
            .I(N__13672));
    CascadeBuf I__2421 (
            .O(N__13675),
            .I(N__13669));
    CascadeMux I__2420 (
            .O(N__13672),
            .I(N__13666));
    CascadeMux I__2419 (
            .O(N__13669),
            .I(N__13663));
    CascadeBuf I__2418 (
            .O(N__13666),
            .I(N__13660));
    CascadeBuf I__2417 (
            .O(N__13663),
            .I(N__13657));
    CascadeMux I__2416 (
            .O(N__13660),
            .I(N__13654));
    CascadeMux I__2415 (
            .O(N__13657),
            .I(N__13651));
    InMux I__2414 (
            .O(N__13654),
            .I(N__13648));
    InMux I__2413 (
            .O(N__13651),
            .I(N__13645));
    LocalMux I__2412 (
            .O(N__13648),
            .I(N__13642));
    LocalMux I__2411 (
            .O(N__13645),
            .I(N__13639));
    Span4Mux_s3_v I__2410 (
            .O(N__13642),
            .I(N__13635));
    Span4Mux_s3_v I__2409 (
            .O(N__13639),
            .I(N__13632));
    InMux I__2408 (
            .O(N__13638),
            .I(N__13629));
    Span4Mux_h I__2407 (
            .O(N__13635),
            .I(N__13626));
    Sp12to4 I__2406 (
            .O(N__13632),
            .I(N__13623));
    LocalMux I__2405 (
            .O(N__13629),
            .I(N__13620));
    Sp12to4 I__2404 (
            .O(N__13626),
            .I(N__13614));
    Span12Mux_h I__2403 (
            .O(N__13623),
            .I(N__13614));
    Span4Mux_h I__2402 (
            .O(N__13620),
            .I(N__13611));
    InMux I__2401 (
            .O(N__13619),
            .I(N__13608));
    Span12Mux_v I__2400 (
            .O(N__13614),
            .I(N__13605));
    Odrv4 I__2399 (
            .O(N__13611),
            .I(RX_ADDR_9));
    LocalMux I__2398 (
            .O(N__13608),
            .I(RX_ADDR_9));
    Odrv12 I__2397 (
            .O(N__13605),
            .I(RX_ADDR_9));
    InMux I__2396 (
            .O(N__13598),
            .I(N__13595));
    LocalMux I__2395 (
            .O(N__13595),
            .I(N__13592));
    Span4Mux_v I__2394 (
            .O(N__13592),
            .I(N__13589));
    Odrv4 I__2393 (
            .O(N__13589),
            .I(\receive_module.n127 ));
    InMux I__2392 (
            .O(N__13586),
            .I(\receive_module.n3331 ));
    InMux I__2391 (
            .O(N__13583),
            .I(N__13579));
    InMux I__2390 (
            .O(N__13582),
            .I(N__13576));
    LocalMux I__2389 (
            .O(N__13579),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    LocalMux I__2388 (
            .O(N__13576),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    InMux I__2387 (
            .O(N__13571),
            .I(N__13567));
    InMux I__2386 (
            .O(N__13570),
            .I(N__13564));
    LocalMux I__2385 (
            .O(N__13567),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    LocalMux I__2384 (
            .O(N__13564),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    InMux I__2383 (
            .O(N__13559),
            .I(N__13555));
    InMux I__2382 (
            .O(N__13558),
            .I(N__13552));
    LocalMux I__2381 (
            .O(N__13555),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    LocalMux I__2380 (
            .O(N__13552),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    InMux I__2379 (
            .O(N__13547),
            .I(N__13543));
    InMux I__2378 (
            .O(N__13546),
            .I(N__13540));
    LocalMux I__2377 (
            .O(N__13543),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    LocalMux I__2376 (
            .O(N__13540),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    InMux I__2375 (
            .O(N__13535),
            .I(N__13531));
    InMux I__2374 (
            .O(N__13534),
            .I(N__13528));
    LocalMux I__2373 (
            .O(N__13531),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    LocalMux I__2372 (
            .O(N__13528),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    InMux I__2371 (
            .O(N__13523),
            .I(N__13519));
    InMux I__2370 (
            .O(N__13522),
            .I(N__13516));
    LocalMux I__2369 (
            .O(N__13519),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    LocalMux I__2368 (
            .O(N__13516),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    CascadeMux I__2367 (
            .O(N__13511),
            .I(\receive_module.rx_counter.n3693_cascade_ ));
    InMux I__2366 (
            .O(N__13508),
            .I(N__13505));
    LocalMux I__2365 (
            .O(N__13505),
            .I(\receive_module.rx_counter.n7 ));
    CascadeMux I__2364 (
            .O(N__13502),
            .I(\receive_module.rx_counter.n11_cascade_ ));
    InMux I__2363 (
            .O(N__13499),
            .I(N__13493));
    InMux I__2362 (
            .O(N__13498),
            .I(N__13493));
    LocalMux I__2361 (
            .O(N__13493),
            .I(N__13490));
    Odrv12 I__2360 (
            .O(N__13490),
            .I(\receive_module.rx_counter.PULSE_1HZ_N_94 ));
    SRMux I__2359 (
            .O(N__13487),
            .I(N__13484));
    LocalMux I__2358 (
            .O(N__13484),
            .I(N__13481));
    Odrv12 I__2357 (
            .O(N__13481),
            .I(\receive_module.rx_counter.n2562 ));
    CascadeMux I__2356 (
            .O(N__13478),
            .I(N__13475));
    CascadeBuf I__2355 (
            .O(N__13475),
            .I(N__13472));
    CascadeMux I__2354 (
            .O(N__13472),
            .I(N__13469));
    CascadeBuf I__2353 (
            .O(N__13469),
            .I(N__13465));
    CascadeMux I__2352 (
            .O(N__13468),
            .I(N__13462));
    CascadeMux I__2351 (
            .O(N__13465),
            .I(N__13459));
    CascadeBuf I__2350 (
            .O(N__13462),
            .I(N__13456));
    CascadeBuf I__2349 (
            .O(N__13459),
            .I(N__13453));
    CascadeMux I__2348 (
            .O(N__13456),
            .I(N__13450));
    CascadeMux I__2347 (
            .O(N__13453),
            .I(N__13447));
    CascadeBuf I__2346 (
            .O(N__13450),
            .I(N__13444));
    CascadeBuf I__2345 (
            .O(N__13447),
            .I(N__13441));
    CascadeMux I__2344 (
            .O(N__13444),
            .I(N__13438));
    CascadeMux I__2343 (
            .O(N__13441),
            .I(N__13435));
    CascadeBuf I__2342 (
            .O(N__13438),
            .I(N__13432));
    CascadeBuf I__2341 (
            .O(N__13435),
            .I(N__13429));
    CascadeMux I__2340 (
            .O(N__13432),
            .I(N__13426));
    CascadeMux I__2339 (
            .O(N__13429),
            .I(N__13423));
    CascadeBuf I__2338 (
            .O(N__13426),
            .I(N__13420));
    CascadeBuf I__2337 (
            .O(N__13423),
            .I(N__13417));
    CascadeMux I__2336 (
            .O(N__13420),
            .I(N__13414));
    CascadeMux I__2335 (
            .O(N__13417),
            .I(N__13411));
    CascadeBuf I__2334 (
            .O(N__13414),
            .I(N__13408));
    CascadeBuf I__2333 (
            .O(N__13411),
            .I(N__13405));
    CascadeMux I__2332 (
            .O(N__13408),
            .I(N__13402));
    CascadeMux I__2331 (
            .O(N__13405),
            .I(N__13399));
    CascadeBuf I__2330 (
            .O(N__13402),
            .I(N__13396));
    CascadeBuf I__2329 (
            .O(N__13399),
            .I(N__13393));
    CascadeMux I__2328 (
            .O(N__13396),
            .I(N__13390));
    CascadeMux I__2327 (
            .O(N__13393),
            .I(N__13387));
    CascadeBuf I__2326 (
            .O(N__13390),
            .I(N__13384));
    CascadeBuf I__2325 (
            .O(N__13387),
            .I(N__13381));
    CascadeMux I__2324 (
            .O(N__13384),
            .I(N__13378));
    CascadeMux I__2323 (
            .O(N__13381),
            .I(N__13375));
    CascadeBuf I__2322 (
            .O(N__13378),
            .I(N__13372));
    CascadeBuf I__2321 (
            .O(N__13375),
            .I(N__13369));
    CascadeMux I__2320 (
            .O(N__13372),
            .I(N__13366));
    CascadeMux I__2319 (
            .O(N__13369),
            .I(N__13363));
    CascadeBuf I__2318 (
            .O(N__13366),
            .I(N__13360));
    CascadeBuf I__2317 (
            .O(N__13363),
            .I(N__13357));
    CascadeMux I__2316 (
            .O(N__13360),
            .I(N__13354));
    CascadeMux I__2315 (
            .O(N__13357),
            .I(N__13351));
    CascadeBuf I__2314 (
            .O(N__13354),
            .I(N__13348));
    CascadeBuf I__2313 (
            .O(N__13351),
            .I(N__13345));
    CascadeMux I__2312 (
            .O(N__13348),
            .I(N__13342));
    CascadeMux I__2311 (
            .O(N__13345),
            .I(N__13339));
    CascadeBuf I__2310 (
            .O(N__13342),
            .I(N__13336));
    CascadeBuf I__2309 (
            .O(N__13339),
            .I(N__13333));
    CascadeMux I__2308 (
            .O(N__13336),
            .I(N__13330));
    CascadeMux I__2307 (
            .O(N__13333),
            .I(N__13327));
    CascadeBuf I__2306 (
            .O(N__13330),
            .I(N__13324));
    CascadeBuf I__2305 (
            .O(N__13327),
            .I(N__13321));
    CascadeMux I__2304 (
            .O(N__13324),
            .I(N__13318));
    CascadeMux I__2303 (
            .O(N__13321),
            .I(N__13315));
    CascadeBuf I__2302 (
            .O(N__13318),
            .I(N__13312));
    CascadeBuf I__2301 (
            .O(N__13315),
            .I(N__13309));
    CascadeMux I__2300 (
            .O(N__13312),
            .I(N__13306));
    CascadeMux I__2299 (
            .O(N__13309),
            .I(N__13303));
    CascadeBuf I__2298 (
            .O(N__13306),
            .I(N__13300));
    InMux I__2297 (
            .O(N__13303),
            .I(N__13297));
    CascadeMux I__2296 (
            .O(N__13300),
            .I(N__13294));
    LocalMux I__2295 (
            .O(N__13297),
            .I(N__13291));
    CascadeBuf I__2294 (
            .O(N__13294),
            .I(N__13288));
    Span4Mux_s1_v I__2293 (
            .O(N__13291),
            .I(N__13285));
    CascadeMux I__2292 (
            .O(N__13288),
            .I(N__13282));
    Span4Mux_h I__2291 (
            .O(N__13285),
            .I(N__13279));
    InMux I__2290 (
            .O(N__13282),
            .I(N__13276));
    Sp12to4 I__2289 (
            .O(N__13279),
            .I(N__13273));
    LocalMux I__2288 (
            .O(N__13276),
            .I(N__13270));
    Span12Mux_s9_v I__2287 (
            .O(N__13273),
            .I(N__13265));
    Span12Mux_s9_v I__2286 (
            .O(N__13270),
            .I(N__13262));
    InMux I__2285 (
            .O(N__13269),
            .I(N__13259));
    InMux I__2284 (
            .O(N__13268),
            .I(N__13256));
    Span12Mux_v I__2283 (
            .O(N__13265),
            .I(N__13253));
    Span12Mux_v I__2282 (
            .O(N__13262),
            .I(N__13250));
    LocalMux I__2281 (
            .O(N__13259),
            .I(RX_ADDR_0));
    LocalMux I__2280 (
            .O(N__13256),
            .I(RX_ADDR_0));
    Odrv12 I__2279 (
            .O(N__13253),
            .I(RX_ADDR_0));
    Odrv12 I__2278 (
            .O(N__13250),
            .I(RX_ADDR_0));
    InMux I__2277 (
            .O(N__13241),
            .I(N__13238));
    LocalMux I__2276 (
            .O(N__13238),
            .I(\receive_module.n136 ));
    InMux I__2275 (
            .O(N__13235),
            .I(bfn_14_11_0_));
    CascadeMux I__2274 (
            .O(N__13232),
            .I(N__13228));
    CascadeMux I__2273 (
            .O(N__13231),
            .I(N__13225));
    CascadeBuf I__2272 (
            .O(N__13228),
            .I(N__13222));
    CascadeBuf I__2271 (
            .O(N__13225),
            .I(N__13219));
    CascadeMux I__2270 (
            .O(N__13222),
            .I(N__13216));
    CascadeMux I__2269 (
            .O(N__13219),
            .I(N__13213));
    CascadeBuf I__2268 (
            .O(N__13216),
            .I(N__13210));
    CascadeBuf I__2267 (
            .O(N__13213),
            .I(N__13207));
    CascadeMux I__2266 (
            .O(N__13210),
            .I(N__13204));
    CascadeMux I__2265 (
            .O(N__13207),
            .I(N__13201));
    CascadeBuf I__2264 (
            .O(N__13204),
            .I(N__13198));
    CascadeBuf I__2263 (
            .O(N__13201),
            .I(N__13195));
    CascadeMux I__2262 (
            .O(N__13198),
            .I(N__13192));
    CascadeMux I__2261 (
            .O(N__13195),
            .I(N__13189));
    CascadeBuf I__2260 (
            .O(N__13192),
            .I(N__13186));
    CascadeBuf I__2259 (
            .O(N__13189),
            .I(N__13183));
    CascadeMux I__2258 (
            .O(N__13186),
            .I(N__13180));
    CascadeMux I__2257 (
            .O(N__13183),
            .I(N__13177));
    CascadeBuf I__2256 (
            .O(N__13180),
            .I(N__13174));
    CascadeBuf I__2255 (
            .O(N__13177),
            .I(N__13171));
    CascadeMux I__2254 (
            .O(N__13174),
            .I(N__13168));
    CascadeMux I__2253 (
            .O(N__13171),
            .I(N__13165));
    CascadeBuf I__2252 (
            .O(N__13168),
            .I(N__13162));
    CascadeBuf I__2251 (
            .O(N__13165),
            .I(N__13159));
    CascadeMux I__2250 (
            .O(N__13162),
            .I(N__13156));
    CascadeMux I__2249 (
            .O(N__13159),
            .I(N__13153));
    CascadeBuf I__2248 (
            .O(N__13156),
            .I(N__13150));
    CascadeBuf I__2247 (
            .O(N__13153),
            .I(N__13147));
    CascadeMux I__2246 (
            .O(N__13150),
            .I(N__13144));
    CascadeMux I__2245 (
            .O(N__13147),
            .I(N__13141));
    CascadeBuf I__2244 (
            .O(N__13144),
            .I(N__13138));
    CascadeBuf I__2243 (
            .O(N__13141),
            .I(N__13135));
    CascadeMux I__2242 (
            .O(N__13138),
            .I(N__13132));
    CascadeMux I__2241 (
            .O(N__13135),
            .I(N__13129));
    CascadeBuf I__2240 (
            .O(N__13132),
            .I(N__13126));
    CascadeBuf I__2239 (
            .O(N__13129),
            .I(N__13123));
    CascadeMux I__2238 (
            .O(N__13126),
            .I(N__13120));
    CascadeMux I__2237 (
            .O(N__13123),
            .I(N__13117));
    CascadeBuf I__2236 (
            .O(N__13120),
            .I(N__13114));
    CascadeBuf I__2235 (
            .O(N__13117),
            .I(N__13111));
    CascadeMux I__2234 (
            .O(N__13114),
            .I(N__13108));
    CascadeMux I__2233 (
            .O(N__13111),
            .I(N__13105));
    CascadeBuf I__2232 (
            .O(N__13108),
            .I(N__13102));
    CascadeBuf I__2231 (
            .O(N__13105),
            .I(N__13099));
    CascadeMux I__2230 (
            .O(N__13102),
            .I(N__13096));
    CascadeMux I__2229 (
            .O(N__13099),
            .I(N__13093));
    CascadeBuf I__2228 (
            .O(N__13096),
            .I(N__13090));
    CascadeBuf I__2227 (
            .O(N__13093),
            .I(N__13087));
    CascadeMux I__2226 (
            .O(N__13090),
            .I(N__13084));
    CascadeMux I__2225 (
            .O(N__13087),
            .I(N__13081));
    CascadeBuf I__2224 (
            .O(N__13084),
            .I(N__13078));
    CascadeBuf I__2223 (
            .O(N__13081),
            .I(N__13075));
    CascadeMux I__2222 (
            .O(N__13078),
            .I(N__13072));
    CascadeMux I__2221 (
            .O(N__13075),
            .I(N__13069));
    CascadeBuf I__2220 (
            .O(N__13072),
            .I(N__13066));
    CascadeBuf I__2219 (
            .O(N__13069),
            .I(N__13063));
    CascadeMux I__2218 (
            .O(N__13066),
            .I(N__13060));
    CascadeMux I__2217 (
            .O(N__13063),
            .I(N__13057));
    CascadeBuf I__2216 (
            .O(N__13060),
            .I(N__13054));
    CascadeBuf I__2215 (
            .O(N__13057),
            .I(N__13051));
    CascadeMux I__2214 (
            .O(N__13054),
            .I(N__13048));
    CascadeMux I__2213 (
            .O(N__13051),
            .I(N__13045));
    InMux I__2212 (
            .O(N__13048),
            .I(N__13042));
    InMux I__2211 (
            .O(N__13045),
            .I(N__13039));
    LocalMux I__2210 (
            .O(N__13042),
            .I(N__13036));
    LocalMux I__2209 (
            .O(N__13039),
            .I(N__13032));
    Span4Mux_s1_v I__2208 (
            .O(N__13036),
            .I(N__13029));
    CascadeMux I__2207 (
            .O(N__13035),
            .I(N__13026));
    Span4Mux_s1_v I__2206 (
            .O(N__13032),
            .I(N__13023));
    Span4Mux_v I__2205 (
            .O(N__13029),
            .I(N__13020));
    InMux I__2204 (
            .O(N__13026),
            .I(N__13017));
    Span4Mux_h I__2203 (
            .O(N__13023),
            .I(N__13014));
    Span4Mux_v I__2202 (
            .O(N__13020),
            .I(N__13011));
    LocalMux I__2201 (
            .O(N__13017),
            .I(N__13007));
    Sp12to4 I__2200 (
            .O(N__13014),
            .I(N__13004));
    Sp12to4 I__2199 (
            .O(N__13011),
            .I(N__13001));
    InMux I__2198 (
            .O(N__13010),
            .I(N__12998));
    Sp12to4 I__2197 (
            .O(N__13007),
            .I(N__12993));
    Span12Mux_s9_v I__2196 (
            .O(N__13004),
            .I(N__12993));
    Span12Mux_s8_h I__2195 (
            .O(N__13001),
            .I(N__12990));
    LocalMux I__2194 (
            .O(N__12998),
            .I(N__12983));
    Span12Mux_v I__2193 (
            .O(N__12993),
            .I(N__12983));
    Span12Mux_v I__2192 (
            .O(N__12990),
            .I(N__12983));
    Odrv12 I__2191 (
            .O(N__12983),
            .I(RX_ADDR_1));
    InMux I__2190 (
            .O(N__12980),
            .I(N__12977));
    LocalMux I__2189 (
            .O(N__12977),
            .I(N__12974));
    Odrv4 I__2188 (
            .O(N__12974),
            .I(\receive_module.n135 ));
    InMux I__2187 (
            .O(N__12971),
            .I(\receive_module.n3323 ));
    InMux I__2186 (
            .O(N__12968),
            .I(\transmit_module.n3348 ));
    InMux I__2185 (
            .O(N__12965),
            .I(N__12962));
    LocalMux I__2184 (
            .O(N__12962),
            .I(N__12959));
    Odrv4 I__2183 (
            .O(N__12959),
            .I(\transmit_module.n191 ));
    InMux I__2182 (
            .O(N__12956),
            .I(N__12948));
    InMux I__2181 (
            .O(N__12955),
            .I(N__12948));
    InMux I__2180 (
            .O(N__12954),
            .I(N__12943));
    InMux I__2179 (
            .O(N__12953),
            .I(N__12943));
    LocalMux I__2178 (
            .O(N__12948),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__2177 (
            .O(N__12943),
            .I(\transmit_module.TX_ADDR_8 ));
    InMux I__2176 (
            .O(N__12938),
            .I(N__12935));
    LocalMux I__2175 (
            .O(N__12935),
            .I(\transmit_module.ADDR_Y_COMPONENT_8 ));
    CascadeMux I__2174 (
            .O(N__12932),
            .I(N__12928));
    InMux I__2173 (
            .O(N__12931),
            .I(N__12925));
    InMux I__2172 (
            .O(N__12928),
            .I(N__12922));
    LocalMux I__2171 (
            .O(N__12925),
            .I(N__12919));
    LocalMux I__2170 (
            .O(N__12922),
            .I(N__12916));
    Odrv4 I__2169 (
            .O(N__12919),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    Odrv4 I__2168 (
            .O(N__12916),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    InMux I__2167 (
            .O(N__12911),
            .I(N__12908));
    LocalMux I__2166 (
            .O(N__12908),
            .I(\transmit_module.X_DELTA_PATTERN_1 ));
    InMux I__2165 (
            .O(N__12905),
            .I(N__12902));
    LocalMux I__2164 (
            .O(N__12902),
            .I(\transmit_module.X_DELTA_PATTERN_2 ));
    InMux I__2163 (
            .O(N__12899),
            .I(N__12896));
    LocalMux I__2162 (
            .O(N__12896),
            .I(\transmit_module.X_DELTA_PATTERN_5 ));
    InMux I__2161 (
            .O(N__12893),
            .I(N__12890));
    LocalMux I__2160 (
            .O(N__12890),
            .I(\transmit_module.X_DELTA_PATTERN_4 ));
    InMux I__2159 (
            .O(N__12887),
            .I(N__12884));
    LocalMux I__2158 (
            .O(N__12884),
            .I(\transmit_module.X_DELTA_PATTERN_3 ));
    CEMux I__2157 (
            .O(N__12881),
            .I(N__12875));
    CEMux I__2156 (
            .O(N__12880),
            .I(N__12871));
    CEMux I__2155 (
            .O(N__12879),
            .I(N__12868));
    CEMux I__2154 (
            .O(N__12878),
            .I(N__12864));
    LocalMux I__2153 (
            .O(N__12875),
            .I(N__12861));
    CEMux I__2152 (
            .O(N__12874),
            .I(N__12858));
    LocalMux I__2151 (
            .O(N__12871),
            .I(N__12855));
    LocalMux I__2150 (
            .O(N__12868),
            .I(N__12852));
    CEMux I__2149 (
            .O(N__12867),
            .I(N__12849));
    LocalMux I__2148 (
            .O(N__12864),
            .I(N__12846));
    Span4Mux_v I__2147 (
            .O(N__12861),
            .I(N__12843));
    LocalMux I__2146 (
            .O(N__12858),
            .I(N__12840));
    Span4Mux_v I__2145 (
            .O(N__12855),
            .I(N__12833));
    Span4Mux_h I__2144 (
            .O(N__12852),
            .I(N__12833));
    LocalMux I__2143 (
            .O(N__12849),
            .I(N__12833));
    Span4Mux_v I__2142 (
            .O(N__12846),
            .I(N__12830));
    Span4Mux_h I__2141 (
            .O(N__12843),
            .I(N__12827));
    Span4Mux_h I__2140 (
            .O(N__12840),
            .I(N__12822));
    Span4Mux_h I__2139 (
            .O(N__12833),
            .I(N__12822));
    Odrv4 I__2138 (
            .O(N__12830),
            .I(\transmit_module.n2099 ));
    Odrv4 I__2137 (
            .O(N__12827),
            .I(\transmit_module.n2099 ));
    Odrv4 I__2136 (
            .O(N__12822),
            .I(\transmit_module.n2099 ));
    InMux I__2135 (
            .O(N__12815),
            .I(N__12812));
    LocalMux I__2134 (
            .O(N__12812),
            .I(\line_buffer.n3788 ));
    InMux I__2133 (
            .O(N__12809),
            .I(N__12806));
    LocalMux I__2132 (
            .O(N__12806),
            .I(N__12803));
    Span4Mux_v I__2131 (
            .O(N__12803),
            .I(N__12800));
    Odrv4 I__2130 (
            .O(N__12800),
            .I(TX_DATA_6));
    InMux I__2129 (
            .O(N__12797),
            .I(\transmit_module.n3339 ));
    InMux I__2128 (
            .O(N__12794),
            .I(N__12791));
    LocalMux I__2127 (
            .O(N__12791),
            .I(\transmit_module.n199 ));
    InMux I__2126 (
            .O(N__12788),
            .I(\transmit_module.n3340 ));
    InMux I__2125 (
            .O(N__12785),
            .I(N__12782));
    LocalMux I__2124 (
            .O(N__12782),
            .I(\transmit_module.n198 ));
    InMux I__2123 (
            .O(N__12779),
            .I(\transmit_module.n3341 ));
    InMux I__2122 (
            .O(N__12776),
            .I(\transmit_module.n3342 ));
    CascadeMux I__2121 (
            .O(N__12773),
            .I(N__12770));
    InMux I__2120 (
            .O(N__12770),
            .I(N__12767));
    LocalMux I__2119 (
            .O(N__12767),
            .I(\transmit_module.n196 ));
    InMux I__2118 (
            .O(N__12764),
            .I(bfn_13_19_0_));
    InMux I__2117 (
            .O(N__12761),
            .I(\transmit_module.n3344 ));
    InMux I__2116 (
            .O(N__12758),
            .I(\transmit_module.n3345 ));
    InMux I__2115 (
            .O(N__12755),
            .I(N__12752));
    LocalMux I__2114 (
            .O(N__12752),
            .I(N__12749));
    Span4Mux_h I__2113 (
            .O(N__12749),
            .I(N__12746));
    Odrv4 I__2112 (
            .O(N__12746),
            .I(\transmit_module.n193 ));
    InMux I__2111 (
            .O(N__12743),
            .I(\transmit_module.n3346 ));
    InMux I__2110 (
            .O(N__12740),
            .I(N__12737));
    LocalMux I__2109 (
            .O(N__12737),
            .I(N__12734));
    Odrv12 I__2108 (
            .O(N__12734),
            .I(\transmit_module.n192 ));
    InMux I__2107 (
            .O(N__12731),
            .I(\transmit_module.n3347 ));
    InMux I__2106 (
            .O(N__12728),
            .I(N__12725));
    LocalMux I__2105 (
            .O(N__12725),
            .I(N__12722));
    Span4Mux_v I__2104 (
            .O(N__12722),
            .I(N__12719));
    Odrv4 I__2103 (
            .O(N__12719),
            .I(\transmit_module.n187 ));
    InMux I__2102 (
            .O(N__12716),
            .I(N__12713));
    LocalMux I__2101 (
            .O(N__12713),
            .I(N__12710));
    Odrv4 I__2100 (
            .O(N__12710),
            .I(\transmit_module.n219 ));
    CascadeMux I__2099 (
            .O(N__12707),
            .I(\transmit_module.n187_cascade_ ));
    InMux I__2098 (
            .O(N__12704),
            .I(N__12701));
    LocalMux I__2097 (
            .O(N__12701),
            .I(\transmit_module.n218 ));
    CascadeMux I__2096 (
            .O(N__12698),
            .I(N__12695));
    InMux I__2095 (
            .O(N__12695),
            .I(N__12689));
    InMux I__2094 (
            .O(N__12694),
            .I(N__12689));
    LocalMux I__2093 (
            .O(N__12689),
            .I(\transmit_module.n186 ));
    CascadeMux I__2092 (
            .O(N__12686),
            .I(N__12683));
    InMux I__2091 (
            .O(N__12683),
            .I(N__12680));
    LocalMux I__2090 (
            .O(N__12680),
            .I(N__12677));
    Odrv4 I__2089 (
            .O(N__12677),
            .I(\transmit_module.n204 ));
    CascadeMux I__2088 (
            .O(N__12674),
            .I(N__12671));
    InMux I__2087 (
            .O(N__12671),
            .I(N__12668));
    LocalMux I__2086 (
            .O(N__12668),
            .I(N__12665));
    Span4Mux_h I__2085 (
            .O(N__12665),
            .I(N__12662));
    Odrv4 I__2084 (
            .O(N__12662),
            .I(\transmit_module.n203 ));
    InMux I__2083 (
            .O(N__12659),
            .I(\transmit_module.n3336 ));
    CascadeMux I__2082 (
            .O(N__12656),
            .I(N__12653));
    InMux I__2081 (
            .O(N__12653),
            .I(N__12650));
    LocalMux I__2080 (
            .O(N__12650),
            .I(N__12647));
    Odrv4 I__2079 (
            .O(N__12647),
            .I(\transmit_module.n202 ));
    InMux I__2078 (
            .O(N__12644),
            .I(\transmit_module.n3337 ));
    InMux I__2077 (
            .O(N__12641),
            .I(\transmit_module.n3338 ));
    IoInMux I__2076 (
            .O(N__12638),
            .I(N__12633));
    IoInMux I__2075 (
            .O(N__12637),
            .I(N__12630));
    IoInMux I__2074 (
            .O(N__12636),
            .I(N__12627));
    LocalMux I__2073 (
            .O(N__12633),
            .I(N__12624));
    LocalMux I__2072 (
            .O(N__12630),
            .I(N__12621));
    LocalMux I__2071 (
            .O(N__12627),
            .I(N__12618));
    Span4Mux_s2_v I__2070 (
            .O(N__12624),
            .I(N__12615));
    Span4Mux_s2_v I__2069 (
            .O(N__12621),
            .I(N__12612));
    Span4Mux_s0_h I__2068 (
            .O(N__12618),
            .I(N__12609));
    Span4Mux_v I__2067 (
            .O(N__12615),
            .I(N__12606));
    Span4Mux_v I__2066 (
            .O(N__12612),
            .I(N__12603));
    Sp12to4 I__2065 (
            .O(N__12609),
            .I(N__12600));
    Sp12to4 I__2064 (
            .O(N__12606),
            .I(N__12597));
    Sp12to4 I__2063 (
            .O(N__12603),
            .I(N__12594));
    Span12Mux_v I__2062 (
            .O(N__12600),
            .I(N__12591));
    Span12Mux_h I__2061 (
            .O(N__12597),
            .I(N__12584));
    Span12Mux_h I__2060 (
            .O(N__12594),
            .I(N__12584));
    Span12Mux_h I__2059 (
            .O(N__12591),
            .I(N__12584));
    Odrv12 I__2058 (
            .O(N__12584),
            .I(n1848));
    IoInMux I__2057 (
            .O(N__12581),
            .I(N__12576));
    IoInMux I__2056 (
            .O(N__12580),
            .I(N__12573));
    IoInMux I__2055 (
            .O(N__12579),
            .I(N__12570));
    LocalMux I__2054 (
            .O(N__12576),
            .I(N__12567));
    LocalMux I__2053 (
            .O(N__12573),
            .I(N__12564));
    LocalMux I__2052 (
            .O(N__12570),
            .I(N__12561));
    Span4Mux_s1_v I__2051 (
            .O(N__12567),
            .I(N__12558));
    IoSpan4Mux I__2050 (
            .O(N__12564),
            .I(N__12555));
    Span4Mux_s1_h I__2049 (
            .O(N__12561),
            .I(N__12552));
    Span4Mux_v I__2048 (
            .O(N__12558),
            .I(N__12549));
    Span4Mux_s3_v I__2047 (
            .O(N__12555),
            .I(N__12546));
    Span4Mux_h I__2046 (
            .O(N__12552),
            .I(N__12543));
    Sp12to4 I__2045 (
            .O(N__12549),
            .I(N__12540));
    Sp12to4 I__2044 (
            .O(N__12546),
            .I(N__12535));
    Sp12to4 I__2043 (
            .O(N__12543),
            .I(N__12535));
    Span12Mux_h I__2042 (
            .O(N__12540),
            .I(N__12532));
    Span12Mux_v I__2041 (
            .O(N__12535),
            .I(N__12529));
    Odrv12 I__2040 (
            .O(N__12532),
            .I(n1847));
    Odrv12 I__2039 (
            .O(N__12529),
            .I(n1847));
    IoInMux I__2038 (
            .O(N__12524),
            .I(N__12520));
    IoInMux I__2037 (
            .O(N__12523),
            .I(N__12517));
    LocalMux I__2036 (
            .O(N__12520),
            .I(N__12513));
    LocalMux I__2035 (
            .O(N__12517),
            .I(N__12510));
    IoInMux I__2034 (
            .O(N__12516),
            .I(N__12507));
    Span4Mux_s0_v I__2033 (
            .O(N__12513),
            .I(N__12504));
    IoSpan4Mux I__2032 (
            .O(N__12510),
            .I(N__12501));
    LocalMux I__2031 (
            .O(N__12507),
            .I(N__12498));
    Sp12to4 I__2030 (
            .O(N__12504),
            .I(N__12495));
    IoSpan4Mux I__2029 (
            .O(N__12501),
            .I(N__12492));
    Span12Mux_s4_v I__2028 (
            .O(N__12498),
            .I(N__12489));
    Span12Mux_h I__2027 (
            .O(N__12495),
            .I(N__12486));
    Sp12to4 I__2026 (
            .O(N__12492),
            .I(N__12483));
    Span12Mux_v I__2025 (
            .O(N__12489),
            .I(N__12480));
    Span12Mux_v I__2024 (
            .O(N__12486),
            .I(N__12475));
    Span12Mux_h I__2023 (
            .O(N__12483),
            .I(N__12475));
    Odrv12 I__2022 (
            .O(N__12480),
            .I(n1846));
    Odrv12 I__2021 (
            .O(N__12475),
            .I(n1846));
    IoInMux I__2020 (
            .O(N__12470),
            .I(N__12465));
    IoInMux I__2019 (
            .O(N__12469),
            .I(N__12462));
    IoInMux I__2018 (
            .O(N__12468),
            .I(N__12459));
    LocalMux I__2017 (
            .O(N__12465),
            .I(N__12456));
    LocalMux I__2016 (
            .O(N__12462),
            .I(N__12453));
    LocalMux I__2015 (
            .O(N__12459),
            .I(N__12450));
    Span4Mux_s2_v I__2014 (
            .O(N__12456),
            .I(N__12447));
    Span12Mux_s4_v I__2013 (
            .O(N__12453),
            .I(N__12444));
    Span4Mux_s3_h I__2012 (
            .O(N__12450),
            .I(N__12441));
    Span4Mux_h I__2011 (
            .O(N__12447),
            .I(N__12438));
    Span12Mux_v I__2010 (
            .O(N__12444),
            .I(N__12435));
    Sp12to4 I__2009 (
            .O(N__12441),
            .I(N__12432));
    Sp12to4 I__2008 (
            .O(N__12438),
            .I(N__12429));
    Span12Mux_h I__2007 (
            .O(N__12435),
            .I(N__12424));
    Span12Mux_v I__2006 (
            .O(N__12432),
            .I(N__12424));
    Span12Mux_s11_v I__2005 (
            .O(N__12429),
            .I(N__12421));
    Odrv12 I__2004 (
            .O(N__12424),
            .I(n1845));
    Odrv12 I__2003 (
            .O(N__12421),
            .I(n1845));
    IoInMux I__2002 (
            .O(N__12416),
            .I(N__12413));
    LocalMux I__2001 (
            .O(N__12413),
            .I(N__12408));
    IoInMux I__2000 (
            .O(N__12412),
            .I(N__12405));
    IoInMux I__1999 (
            .O(N__12411),
            .I(N__12402));
    Span4Mux_s0_v I__1998 (
            .O(N__12408),
            .I(N__12399));
    LocalMux I__1997 (
            .O(N__12405),
            .I(N__12396));
    LocalMux I__1996 (
            .O(N__12402),
            .I(N__12393));
    Span4Mux_v I__1995 (
            .O(N__12399),
            .I(N__12390));
    Span4Mux_s0_h I__1994 (
            .O(N__12396),
            .I(N__12387));
    IoSpan4Mux I__1993 (
            .O(N__12393),
            .I(N__12384));
    Sp12to4 I__1992 (
            .O(N__12390),
            .I(N__12381));
    Sp12to4 I__1991 (
            .O(N__12387),
            .I(N__12378));
    Span4Mux_s2_v I__1990 (
            .O(N__12384),
            .I(N__12375));
    Span12Mux_s9_h I__1989 (
            .O(N__12381),
            .I(N__12372));
    Span12Mux_s10_v I__1988 (
            .O(N__12378),
            .I(N__12369));
    Sp12to4 I__1987 (
            .O(N__12375),
            .I(N__12366));
    Span12Mux_v I__1986 (
            .O(N__12372),
            .I(N__12363));
    Span12Mux_h I__1985 (
            .O(N__12369),
            .I(N__12358));
    Span12Mux_s10_v I__1984 (
            .O(N__12366),
            .I(N__12358));
    Odrv12 I__1983 (
            .O(N__12363),
            .I(n1844));
    Odrv12 I__1982 (
            .O(N__12358),
            .I(n1844));
    IoInMux I__1981 (
            .O(N__12353),
            .I(N__12350));
    LocalMux I__1980 (
            .O(N__12350),
            .I(N__12346));
    IoInMux I__1979 (
            .O(N__12349),
            .I(N__12342));
    IoSpan4Mux I__1978 (
            .O(N__12346),
            .I(N__12339));
    IoInMux I__1977 (
            .O(N__12345),
            .I(N__12336));
    LocalMux I__1976 (
            .O(N__12342),
            .I(N__12333));
    Span4Mux_s0_v I__1975 (
            .O(N__12339),
            .I(N__12330));
    LocalMux I__1974 (
            .O(N__12336),
            .I(N__12327));
    Span4Mux_s0_h I__1973 (
            .O(N__12333),
            .I(N__12324));
    Span4Mux_v I__1972 (
            .O(N__12330),
            .I(N__12321));
    IoSpan4Mux I__1971 (
            .O(N__12327),
            .I(N__12318));
    Sp12to4 I__1970 (
            .O(N__12324),
            .I(N__12315));
    Sp12to4 I__1969 (
            .O(N__12321),
            .I(N__12312));
    Span4Mux_s3_v I__1968 (
            .O(N__12318),
            .I(N__12309));
    Span12Mux_s9_v I__1967 (
            .O(N__12315),
            .I(N__12306));
    Span12Mux_h I__1966 (
            .O(N__12312),
            .I(N__12301));
    Sp12to4 I__1965 (
            .O(N__12309),
            .I(N__12301));
    Span12Mux_h I__1964 (
            .O(N__12306),
            .I(N__12298));
    Span12Mux_v I__1963 (
            .O(N__12301),
            .I(N__12295));
    Odrv12 I__1962 (
            .O(N__12298),
            .I(ADV_B_c));
    Odrv12 I__1961 (
            .O(N__12295),
            .I(ADV_B_c));
    SRMux I__1960 (
            .O(N__12290),
            .I(N__12287));
    LocalMux I__1959 (
            .O(N__12287),
            .I(N__12284));
    Span4Mux_h I__1958 (
            .O(N__12284),
            .I(N__12281));
    Odrv4 I__1957 (
            .O(N__12281),
            .I(n2404));
    InMux I__1956 (
            .O(N__12278),
            .I(N__12275));
    LocalMux I__1955 (
            .O(N__12275),
            .I(N__12272));
    Odrv4 I__1954 (
            .O(N__12272),
            .I(\transmit_module.n220 ));
    CascadeMux I__1953 (
            .O(N__12269),
            .I(\transmit_module.n218_cascade_ ));
    CascadeMux I__1952 (
            .O(N__12266),
            .I(N__12263));
    CascadeBuf I__1951 (
            .O(N__12263),
            .I(N__12259));
    CascadeMux I__1950 (
            .O(N__12262),
            .I(N__12256));
    CascadeMux I__1949 (
            .O(N__12259),
            .I(N__12253));
    CascadeBuf I__1948 (
            .O(N__12256),
            .I(N__12250));
    CascadeBuf I__1947 (
            .O(N__12253),
            .I(N__12247));
    CascadeMux I__1946 (
            .O(N__12250),
            .I(N__12244));
    CascadeMux I__1945 (
            .O(N__12247),
            .I(N__12241));
    CascadeBuf I__1944 (
            .O(N__12244),
            .I(N__12238));
    CascadeBuf I__1943 (
            .O(N__12241),
            .I(N__12235));
    CascadeMux I__1942 (
            .O(N__12238),
            .I(N__12232));
    CascadeMux I__1941 (
            .O(N__12235),
            .I(N__12229));
    CascadeBuf I__1940 (
            .O(N__12232),
            .I(N__12226));
    CascadeBuf I__1939 (
            .O(N__12229),
            .I(N__12223));
    CascadeMux I__1938 (
            .O(N__12226),
            .I(N__12220));
    CascadeMux I__1937 (
            .O(N__12223),
            .I(N__12217));
    CascadeBuf I__1936 (
            .O(N__12220),
            .I(N__12214));
    CascadeBuf I__1935 (
            .O(N__12217),
            .I(N__12211));
    CascadeMux I__1934 (
            .O(N__12214),
            .I(N__12208));
    CascadeMux I__1933 (
            .O(N__12211),
            .I(N__12205));
    CascadeBuf I__1932 (
            .O(N__12208),
            .I(N__12202));
    CascadeBuf I__1931 (
            .O(N__12205),
            .I(N__12199));
    CascadeMux I__1930 (
            .O(N__12202),
            .I(N__12196));
    CascadeMux I__1929 (
            .O(N__12199),
            .I(N__12193));
    CascadeBuf I__1928 (
            .O(N__12196),
            .I(N__12190));
    CascadeBuf I__1927 (
            .O(N__12193),
            .I(N__12187));
    CascadeMux I__1926 (
            .O(N__12190),
            .I(N__12184));
    CascadeMux I__1925 (
            .O(N__12187),
            .I(N__12181));
    CascadeBuf I__1924 (
            .O(N__12184),
            .I(N__12178));
    CascadeBuf I__1923 (
            .O(N__12181),
            .I(N__12175));
    CascadeMux I__1922 (
            .O(N__12178),
            .I(N__12172));
    CascadeMux I__1921 (
            .O(N__12175),
            .I(N__12169));
    CascadeBuf I__1920 (
            .O(N__12172),
            .I(N__12166));
    CascadeBuf I__1919 (
            .O(N__12169),
            .I(N__12163));
    CascadeMux I__1918 (
            .O(N__12166),
            .I(N__12160));
    CascadeMux I__1917 (
            .O(N__12163),
            .I(N__12157));
    CascadeBuf I__1916 (
            .O(N__12160),
            .I(N__12154));
    CascadeBuf I__1915 (
            .O(N__12157),
            .I(N__12151));
    CascadeMux I__1914 (
            .O(N__12154),
            .I(N__12148));
    CascadeMux I__1913 (
            .O(N__12151),
            .I(N__12145));
    CascadeBuf I__1912 (
            .O(N__12148),
            .I(N__12142));
    CascadeBuf I__1911 (
            .O(N__12145),
            .I(N__12139));
    CascadeMux I__1910 (
            .O(N__12142),
            .I(N__12136));
    CascadeMux I__1909 (
            .O(N__12139),
            .I(N__12133));
    CascadeBuf I__1908 (
            .O(N__12136),
            .I(N__12130));
    CascadeBuf I__1907 (
            .O(N__12133),
            .I(N__12127));
    CascadeMux I__1906 (
            .O(N__12130),
            .I(N__12124));
    CascadeMux I__1905 (
            .O(N__12127),
            .I(N__12121));
    CascadeBuf I__1904 (
            .O(N__12124),
            .I(N__12118));
    CascadeBuf I__1903 (
            .O(N__12121),
            .I(N__12115));
    CascadeMux I__1902 (
            .O(N__12118),
            .I(N__12112));
    CascadeMux I__1901 (
            .O(N__12115),
            .I(N__12109));
    CascadeBuf I__1900 (
            .O(N__12112),
            .I(N__12106));
    CascadeBuf I__1899 (
            .O(N__12109),
            .I(N__12103));
    CascadeMux I__1898 (
            .O(N__12106),
            .I(N__12100));
    CascadeMux I__1897 (
            .O(N__12103),
            .I(N__12097));
    CascadeBuf I__1896 (
            .O(N__12100),
            .I(N__12094));
    CascadeBuf I__1895 (
            .O(N__12097),
            .I(N__12091));
    CascadeMux I__1894 (
            .O(N__12094),
            .I(N__12088));
    CascadeMux I__1893 (
            .O(N__12091),
            .I(N__12085));
    CascadeBuf I__1892 (
            .O(N__12088),
            .I(N__12082));
    InMux I__1891 (
            .O(N__12085),
            .I(N__12079));
    CascadeMux I__1890 (
            .O(N__12082),
            .I(N__12076));
    LocalMux I__1889 (
            .O(N__12079),
            .I(N__12073));
    InMux I__1888 (
            .O(N__12076),
            .I(N__12070));
    Span12Mux_v I__1887 (
            .O(N__12073),
            .I(N__12067));
    LocalMux I__1886 (
            .O(N__12070),
            .I(N__12064));
    Span12Mux_h I__1885 (
            .O(N__12067),
            .I(N__12059));
    Span12Mux_h I__1884 (
            .O(N__12064),
            .I(N__12059));
    Span12Mux_v I__1883 (
            .O(N__12059),
            .I(N__12056));
    Odrv12 I__1882 (
            .O(N__12056),
            .I(n26));
    CascadeMux I__1881 (
            .O(N__12053),
            .I(N__12050));
    InMux I__1880 (
            .O(N__12050),
            .I(N__12046));
    InMux I__1879 (
            .O(N__12049),
            .I(N__12041));
    LocalMux I__1878 (
            .O(N__12046),
            .I(N__12038));
    InMux I__1877 (
            .O(N__12045),
            .I(N__12035));
    InMux I__1876 (
            .O(N__12044),
            .I(N__12032));
    LocalMux I__1875 (
            .O(N__12041),
            .I(\transmit_module.video_signal_controller.n3857 ));
    Odrv4 I__1874 (
            .O(N__12038),
            .I(\transmit_module.video_signal_controller.n3857 ));
    LocalMux I__1873 (
            .O(N__12035),
            .I(\transmit_module.video_signal_controller.n3857 ));
    LocalMux I__1872 (
            .O(N__12032),
            .I(\transmit_module.video_signal_controller.n3857 ));
    InMux I__1871 (
            .O(N__12023),
            .I(N__12020));
    LocalMux I__1870 (
            .O(N__12020),
            .I(N__12013));
    InMux I__1869 (
            .O(N__12019),
            .I(N__12006));
    InMux I__1868 (
            .O(N__12018),
            .I(N__12006));
    InMux I__1867 (
            .O(N__12017),
            .I(N__12003));
    InMux I__1866 (
            .O(N__12016),
            .I(N__12000));
    Span4Mux_v I__1865 (
            .O(N__12013),
            .I(N__11997));
    InMux I__1864 (
            .O(N__12012),
            .I(N__11994));
    InMux I__1863 (
            .O(N__12011),
            .I(N__11991));
    LocalMux I__1862 (
            .O(N__12006),
            .I(N__11988));
    LocalMux I__1861 (
            .O(N__12003),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    LocalMux I__1860 (
            .O(N__12000),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    Odrv4 I__1859 (
            .O(N__11997),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    LocalMux I__1858 (
            .O(N__11994),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    LocalMux I__1857 (
            .O(N__11991),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    Odrv4 I__1856 (
            .O(N__11988),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    CascadeMux I__1855 (
            .O(N__11975),
            .I(N__11971));
    CascadeMux I__1854 (
            .O(N__11974),
            .I(N__11968));
    InMux I__1853 (
            .O(N__11971),
            .I(N__11965));
    InMux I__1852 (
            .O(N__11968),
            .I(N__11962));
    LocalMux I__1851 (
            .O(N__11965),
            .I(\transmit_module.video_signal_controller.n3856 ));
    LocalMux I__1850 (
            .O(N__11962),
            .I(\transmit_module.video_signal_controller.n3856 ));
    CascadeMux I__1849 (
            .O(N__11957),
            .I(\transmit_module.n220_cascade_ ));
    CascadeMux I__1848 (
            .O(N__11954),
            .I(N__11951));
    CascadeBuf I__1847 (
            .O(N__11951),
            .I(N__11947));
    CascadeMux I__1846 (
            .O(N__11950),
            .I(N__11944));
    CascadeMux I__1845 (
            .O(N__11947),
            .I(N__11941));
    CascadeBuf I__1844 (
            .O(N__11944),
            .I(N__11938));
    CascadeBuf I__1843 (
            .O(N__11941),
            .I(N__11935));
    CascadeMux I__1842 (
            .O(N__11938),
            .I(N__11932));
    CascadeMux I__1841 (
            .O(N__11935),
            .I(N__11929));
    CascadeBuf I__1840 (
            .O(N__11932),
            .I(N__11926));
    CascadeBuf I__1839 (
            .O(N__11929),
            .I(N__11923));
    CascadeMux I__1838 (
            .O(N__11926),
            .I(N__11920));
    CascadeMux I__1837 (
            .O(N__11923),
            .I(N__11917));
    CascadeBuf I__1836 (
            .O(N__11920),
            .I(N__11914));
    CascadeBuf I__1835 (
            .O(N__11917),
            .I(N__11911));
    CascadeMux I__1834 (
            .O(N__11914),
            .I(N__11908));
    CascadeMux I__1833 (
            .O(N__11911),
            .I(N__11905));
    CascadeBuf I__1832 (
            .O(N__11908),
            .I(N__11902));
    CascadeBuf I__1831 (
            .O(N__11905),
            .I(N__11899));
    CascadeMux I__1830 (
            .O(N__11902),
            .I(N__11896));
    CascadeMux I__1829 (
            .O(N__11899),
            .I(N__11893));
    CascadeBuf I__1828 (
            .O(N__11896),
            .I(N__11890));
    CascadeBuf I__1827 (
            .O(N__11893),
            .I(N__11887));
    CascadeMux I__1826 (
            .O(N__11890),
            .I(N__11884));
    CascadeMux I__1825 (
            .O(N__11887),
            .I(N__11881));
    CascadeBuf I__1824 (
            .O(N__11884),
            .I(N__11878));
    CascadeBuf I__1823 (
            .O(N__11881),
            .I(N__11875));
    CascadeMux I__1822 (
            .O(N__11878),
            .I(N__11872));
    CascadeMux I__1821 (
            .O(N__11875),
            .I(N__11869));
    CascadeBuf I__1820 (
            .O(N__11872),
            .I(N__11866));
    CascadeBuf I__1819 (
            .O(N__11869),
            .I(N__11863));
    CascadeMux I__1818 (
            .O(N__11866),
            .I(N__11860));
    CascadeMux I__1817 (
            .O(N__11863),
            .I(N__11857));
    CascadeBuf I__1816 (
            .O(N__11860),
            .I(N__11854));
    CascadeBuf I__1815 (
            .O(N__11857),
            .I(N__11851));
    CascadeMux I__1814 (
            .O(N__11854),
            .I(N__11848));
    CascadeMux I__1813 (
            .O(N__11851),
            .I(N__11845));
    CascadeBuf I__1812 (
            .O(N__11848),
            .I(N__11842));
    CascadeBuf I__1811 (
            .O(N__11845),
            .I(N__11839));
    CascadeMux I__1810 (
            .O(N__11842),
            .I(N__11836));
    CascadeMux I__1809 (
            .O(N__11839),
            .I(N__11833));
    CascadeBuf I__1808 (
            .O(N__11836),
            .I(N__11830));
    CascadeBuf I__1807 (
            .O(N__11833),
            .I(N__11827));
    CascadeMux I__1806 (
            .O(N__11830),
            .I(N__11824));
    CascadeMux I__1805 (
            .O(N__11827),
            .I(N__11821));
    CascadeBuf I__1804 (
            .O(N__11824),
            .I(N__11818));
    CascadeBuf I__1803 (
            .O(N__11821),
            .I(N__11815));
    CascadeMux I__1802 (
            .O(N__11818),
            .I(N__11812));
    CascadeMux I__1801 (
            .O(N__11815),
            .I(N__11809));
    CascadeBuf I__1800 (
            .O(N__11812),
            .I(N__11806));
    CascadeBuf I__1799 (
            .O(N__11809),
            .I(N__11803));
    CascadeMux I__1798 (
            .O(N__11806),
            .I(N__11800));
    CascadeMux I__1797 (
            .O(N__11803),
            .I(N__11797));
    CascadeBuf I__1796 (
            .O(N__11800),
            .I(N__11794));
    CascadeBuf I__1795 (
            .O(N__11797),
            .I(N__11791));
    CascadeMux I__1794 (
            .O(N__11794),
            .I(N__11788));
    CascadeMux I__1793 (
            .O(N__11791),
            .I(N__11785));
    CascadeBuf I__1792 (
            .O(N__11788),
            .I(N__11782));
    CascadeBuf I__1791 (
            .O(N__11785),
            .I(N__11779));
    CascadeMux I__1790 (
            .O(N__11782),
            .I(N__11776));
    CascadeMux I__1789 (
            .O(N__11779),
            .I(N__11773));
    CascadeBuf I__1788 (
            .O(N__11776),
            .I(N__11770));
    InMux I__1787 (
            .O(N__11773),
            .I(N__11767));
    CascadeMux I__1786 (
            .O(N__11770),
            .I(N__11764));
    LocalMux I__1785 (
            .O(N__11767),
            .I(N__11761));
    InMux I__1784 (
            .O(N__11764),
            .I(N__11758));
    Span4Mux_h I__1783 (
            .O(N__11761),
            .I(N__11755));
    LocalMux I__1782 (
            .O(N__11758),
            .I(N__11752));
    Span4Mux_h I__1781 (
            .O(N__11755),
            .I(N__11749));
    Span12Mux_s7_v I__1780 (
            .O(N__11752),
            .I(N__11746));
    Sp12to4 I__1779 (
            .O(N__11749),
            .I(N__11743));
    Span12Mux_h I__1778 (
            .O(N__11746),
            .I(N__11738));
    Span12Mux_s7_v I__1777 (
            .O(N__11743),
            .I(N__11738));
    Odrv12 I__1776 (
            .O(N__11738),
            .I(n28));
    InMux I__1775 (
            .O(N__11735),
            .I(N__11732));
    LocalMux I__1774 (
            .O(N__11732),
            .I(\transmit_module.BRAM_ADDR_13_N_256_13 ));
    CascadeMux I__1773 (
            .O(N__11729),
            .I(\transmit_module.n219_cascade_ ));
    CascadeMux I__1772 (
            .O(N__11726),
            .I(N__11722));
    CascadeMux I__1771 (
            .O(N__11725),
            .I(N__11719));
    CascadeBuf I__1770 (
            .O(N__11722),
            .I(N__11716));
    CascadeBuf I__1769 (
            .O(N__11719),
            .I(N__11713));
    CascadeMux I__1768 (
            .O(N__11716),
            .I(N__11710));
    CascadeMux I__1767 (
            .O(N__11713),
            .I(N__11707));
    CascadeBuf I__1766 (
            .O(N__11710),
            .I(N__11704));
    CascadeBuf I__1765 (
            .O(N__11707),
            .I(N__11701));
    CascadeMux I__1764 (
            .O(N__11704),
            .I(N__11698));
    CascadeMux I__1763 (
            .O(N__11701),
            .I(N__11695));
    CascadeBuf I__1762 (
            .O(N__11698),
            .I(N__11692));
    CascadeBuf I__1761 (
            .O(N__11695),
            .I(N__11689));
    CascadeMux I__1760 (
            .O(N__11692),
            .I(N__11686));
    CascadeMux I__1759 (
            .O(N__11689),
            .I(N__11683));
    CascadeBuf I__1758 (
            .O(N__11686),
            .I(N__11680));
    CascadeBuf I__1757 (
            .O(N__11683),
            .I(N__11677));
    CascadeMux I__1756 (
            .O(N__11680),
            .I(N__11674));
    CascadeMux I__1755 (
            .O(N__11677),
            .I(N__11671));
    CascadeBuf I__1754 (
            .O(N__11674),
            .I(N__11668));
    CascadeBuf I__1753 (
            .O(N__11671),
            .I(N__11665));
    CascadeMux I__1752 (
            .O(N__11668),
            .I(N__11662));
    CascadeMux I__1751 (
            .O(N__11665),
            .I(N__11659));
    CascadeBuf I__1750 (
            .O(N__11662),
            .I(N__11656));
    CascadeBuf I__1749 (
            .O(N__11659),
            .I(N__11653));
    CascadeMux I__1748 (
            .O(N__11656),
            .I(N__11650));
    CascadeMux I__1747 (
            .O(N__11653),
            .I(N__11647));
    CascadeBuf I__1746 (
            .O(N__11650),
            .I(N__11644));
    CascadeBuf I__1745 (
            .O(N__11647),
            .I(N__11641));
    CascadeMux I__1744 (
            .O(N__11644),
            .I(N__11638));
    CascadeMux I__1743 (
            .O(N__11641),
            .I(N__11635));
    CascadeBuf I__1742 (
            .O(N__11638),
            .I(N__11632));
    CascadeBuf I__1741 (
            .O(N__11635),
            .I(N__11629));
    CascadeMux I__1740 (
            .O(N__11632),
            .I(N__11626));
    CascadeMux I__1739 (
            .O(N__11629),
            .I(N__11623));
    CascadeBuf I__1738 (
            .O(N__11626),
            .I(N__11620));
    CascadeBuf I__1737 (
            .O(N__11623),
            .I(N__11617));
    CascadeMux I__1736 (
            .O(N__11620),
            .I(N__11614));
    CascadeMux I__1735 (
            .O(N__11617),
            .I(N__11611));
    CascadeBuf I__1734 (
            .O(N__11614),
            .I(N__11608));
    CascadeBuf I__1733 (
            .O(N__11611),
            .I(N__11605));
    CascadeMux I__1732 (
            .O(N__11608),
            .I(N__11602));
    CascadeMux I__1731 (
            .O(N__11605),
            .I(N__11599));
    CascadeBuf I__1730 (
            .O(N__11602),
            .I(N__11596));
    CascadeBuf I__1729 (
            .O(N__11599),
            .I(N__11593));
    CascadeMux I__1728 (
            .O(N__11596),
            .I(N__11590));
    CascadeMux I__1727 (
            .O(N__11593),
            .I(N__11587));
    CascadeBuf I__1726 (
            .O(N__11590),
            .I(N__11584));
    CascadeBuf I__1725 (
            .O(N__11587),
            .I(N__11581));
    CascadeMux I__1724 (
            .O(N__11584),
            .I(N__11578));
    CascadeMux I__1723 (
            .O(N__11581),
            .I(N__11575));
    CascadeBuf I__1722 (
            .O(N__11578),
            .I(N__11572));
    CascadeBuf I__1721 (
            .O(N__11575),
            .I(N__11569));
    CascadeMux I__1720 (
            .O(N__11572),
            .I(N__11566));
    CascadeMux I__1719 (
            .O(N__11569),
            .I(N__11563));
    CascadeBuf I__1718 (
            .O(N__11566),
            .I(N__11560));
    CascadeBuf I__1717 (
            .O(N__11563),
            .I(N__11557));
    CascadeMux I__1716 (
            .O(N__11560),
            .I(N__11554));
    CascadeMux I__1715 (
            .O(N__11557),
            .I(N__11551));
    CascadeBuf I__1714 (
            .O(N__11554),
            .I(N__11548));
    CascadeBuf I__1713 (
            .O(N__11551),
            .I(N__11545));
    CascadeMux I__1712 (
            .O(N__11548),
            .I(N__11542));
    CascadeMux I__1711 (
            .O(N__11545),
            .I(N__11539));
    InMux I__1710 (
            .O(N__11542),
            .I(N__11536));
    InMux I__1709 (
            .O(N__11539),
            .I(N__11533));
    LocalMux I__1708 (
            .O(N__11536),
            .I(N__11530));
    LocalMux I__1707 (
            .O(N__11533),
            .I(N__11527));
    Span4Mux_h I__1706 (
            .O(N__11530),
            .I(N__11524));
    Span12Mux_s11_v I__1705 (
            .O(N__11527),
            .I(N__11521));
    Span4Mux_h I__1704 (
            .O(N__11524),
            .I(N__11518));
    Span12Mux_h I__1703 (
            .O(N__11521),
            .I(N__11513));
    Sp12to4 I__1702 (
            .O(N__11518),
            .I(N__11513));
    Span12Mux_s11_v I__1701 (
            .O(N__11513),
            .I(N__11510));
    Odrv12 I__1700 (
            .O(N__11510),
            .I(n27));
    IoInMux I__1699 (
            .O(N__11507),
            .I(N__11503));
    IoInMux I__1698 (
            .O(N__11506),
            .I(N__11500));
    LocalMux I__1697 (
            .O(N__11503),
            .I(N__11497));
    LocalMux I__1696 (
            .O(N__11500),
            .I(N__11493));
    IoSpan4Mux I__1695 (
            .O(N__11497),
            .I(N__11490));
    IoInMux I__1694 (
            .O(N__11496),
            .I(N__11487));
    IoSpan4Mux I__1693 (
            .O(N__11493),
            .I(N__11484));
    IoSpan4Mux I__1692 (
            .O(N__11490),
            .I(N__11479));
    LocalMux I__1691 (
            .O(N__11487),
            .I(N__11479));
    Span4Mux_s0_h I__1690 (
            .O(N__11484),
            .I(N__11476));
    IoSpan4Mux I__1689 (
            .O(N__11479),
            .I(N__11473));
    Sp12to4 I__1688 (
            .O(N__11476),
            .I(N__11470));
    Span4Mux_s2_v I__1687 (
            .O(N__11473),
            .I(N__11467));
    Span12Mux_v I__1686 (
            .O(N__11470),
            .I(N__11464));
    Sp12to4 I__1685 (
            .O(N__11467),
            .I(N__11461));
    Span12Mux_h I__1684 (
            .O(N__11464),
            .I(N__11456));
    Span12Mux_s8_v I__1683 (
            .O(N__11461),
            .I(N__11456));
    Odrv12 I__1682 (
            .O(N__11456),
            .I(n1850));
    IoInMux I__1681 (
            .O(N__11453),
            .I(N__11450));
    LocalMux I__1680 (
            .O(N__11450),
            .I(N__11445));
    IoInMux I__1679 (
            .O(N__11449),
            .I(N__11442));
    IoInMux I__1678 (
            .O(N__11448),
            .I(N__11439));
    IoSpan4Mux I__1677 (
            .O(N__11445),
            .I(N__11436));
    LocalMux I__1676 (
            .O(N__11442),
            .I(N__11433));
    LocalMux I__1675 (
            .O(N__11439),
            .I(N__11430));
    IoSpan4Mux I__1674 (
            .O(N__11436),
            .I(N__11427));
    Span4Mux_s3_h I__1673 (
            .O(N__11433),
            .I(N__11424));
    Span4Mux_s3_v I__1672 (
            .O(N__11430),
            .I(N__11421));
    Span4Mux_s3_v I__1671 (
            .O(N__11427),
            .I(N__11418));
    Span4Mux_h I__1670 (
            .O(N__11424),
            .I(N__11415));
    Span4Mux_v I__1669 (
            .O(N__11421),
            .I(N__11412));
    Sp12to4 I__1668 (
            .O(N__11418),
            .I(N__11407));
    Sp12to4 I__1667 (
            .O(N__11415),
            .I(N__11407));
    Sp12to4 I__1666 (
            .O(N__11412),
            .I(N__11404));
    Span12Mux_v I__1665 (
            .O(N__11407),
            .I(N__11401));
    Span12Mux_h I__1664 (
            .O(N__11404),
            .I(N__11398));
    Odrv12 I__1663 (
            .O(N__11401),
            .I(n1849));
    Odrv12 I__1662 (
            .O(N__11398),
            .I(n1849));
    CascadeMux I__1661 (
            .O(N__11393),
            .I(\transmit_module.video_signal_controller.n3023_cascade_ ));
    CascadeMux I__1660 (
            .O(N__11390),
            .I(\transmit_module.video_signal_controller.n3697_cascade_ ));
    InMux I__1659 (
            .O(N__11387),
            .I(N__11384));
    LocalMux I__1658 (
            .O(N__11384),
            .I(\transmit_module.video_signal_controller.n8 ));
    InMux I__1657 (
            .O(N__11381),
            .I(N__11378));
    LocalMux I__1656 (
            .O(N__11378),
            .I(\transmit_module.video_signal_controller.n3577 ));
    CascadeMux I__1655 (
            .O(N__11375),
            .I(\transmit_module.video_signal_controller.n6_adj_568_cascade_ ));
    InMux I__1654 (
            .O(N__11372),
            .I(N__11369));
    LocalMux I__1653 (
            .O(N__11369),
            .I(\transmit_module.video_signal_controller.n3603 ));
    CascadeMux I__1652 (
            .O(N__11366),
            .I(\transmit_module.video_signal_controller.n6_cascade_ ));
    InMux I__1651 (
            .O(N__11363),
            .I(N__11359));
    InMux I__1650 (
            .O(N__11362),
            .I(N__11356));
    LocalMux I__1649 (
            .O(N__11359),
            .I(\transmit_module.video_signal_controller.n3575 ));
    LocalMux I__1648 (
            .O(N__11356),
            .I(\transmit_module.video_signal_controller.n3575 ));
    InMux I__1647 (
            .O(N__11351),
            .I(N__11347));
    InMux I__1646 (
            .O(N__11350),
            .I(N__11344));
    LocalMux I__1645 (
            .O(N__11347),
            .I(\transmit_module.video_signal_controller.n2015 ));
    LocalMux I__1644 (
            .O(N__11344),
            .I(\transmit_module.video_signal_controller.n2015 ));
    InMux I__1643 (
            .O(N__11339),
            .I(\receive_module.rx_counter.n3390 ));
    InMux I__1642 (
            .O(N__11336),
            .I(\receive_module.rx_counter.n3391 ));
    IoInMux I__1641 (
            .O(N__11333),
            .I(N__11330));
    LocalMux I__1640 (
            .O(N__11330),
            .I(N__11327));
    IoSpan4Mux I__1639 (
            .O(N__11327),
            .I(N__11324));
    IoSpan4Mux I__1638 (
            .O(N__11324),
            .I(N__11321));
    Sp12to4 I__1637 (
            .O(N__11321),
            .I(N__11305));
    InMux I__1636 (
            .O(N__11320),
            .I(N__11287));
    InMux I__1635 (
            .O(N__11319),
            .I(N__11287));
    InMux I__1634 (
            .O(N__11318),
            .I(N__11287));
    InMux I__1633 (
            .O(N__11317),
            .I(N__11287));
    InMux I__1632 (
            .O(N__11316),
            .I(N__11287));
    InMux I__1631 (
            .O(N__11315),
            .I(N__11270));
    InMux I__1630 (
            .O(N__11314),
            .I(N__11270));
    InMux I__1629 (
            .O(N__11313),
            .I(N__11270));
    InMux I__1628 (
            .O(N__11312),
            .I(N__11270));
    InMux I__1627 (
            .O(N__11311),
            .I(N__11270));
    InMux I__1626 (
            .O(N__11310),
            .I(N__11270));
    InMux I__1625 (
            .O(N__11309),
            .I(N__11270));
    InMux I__1624 (
            .O(N__11308),
            .I(N__11270));
    Span12Mux_h I__1623 (
            .O(N__11305),
            .I(N__11267));
    InMux I__1622 (
            .O(N__11304),
            .I(N__11264));
    InMux I__1621 (
            .O(N__11303),
            .I(N__11259));
    InMux I__1620 (
            .O(N__11302),
            .I(N__11259));
    InMux I__1619 (
            .O(N__11301),
            .I(N__11250));
    InMux I__1618 (
            .O(N__11300),
            .I(N__11250));
    InMux I__1617 (
            .O(N__11299),
            .I(N__11250));
    InMux I__1616 (
            .O(N__11298),
            .I(N__11250));
    LocalMux I__1615 (
            .O(N__11287),
            .I(N__11245));
    LocalMux I__1614 (
            .O(N__11270),
            .I(N__11245));
    Odrv12 I__1613 (
            .O(N__11267),
            .I(DEBUG_c_5));
    LocalMux I__1612 (
            .O(N__11264),
            .I(DEBUG_c_5));
    LocalMux I__1611 (
            .O(N__11259),
            .I(DEBUG_c_5));
    LocalMux I__1610 (
            .O(N__11250),
            .I(DEBUG_c_5));
    Odrv4 I__1609 (
            .O(N__11245),
            .I(DEBUG_c_5));
    InMux I__1608 (
            .O(N__11234),
            .I(N__11231));
    LocalMux I__1607 (
            .O(N__11231),
            .I(N__11227));
    InMux I__1606 (
            .O(N__11230),
            .I(N__11222));
    Span4Mux_h I__1605 (
            .O(N__11227),
            .I(N__11219));
    InMux I__1604 (
            .O(N__11226),
            .I(N__11216));
    InMux I__1603 (
            .O(N__11225),
            .I(N__11213));
    LocalMux I__1602 (
            .O(N__11222),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    Odrv4 I__1601 (
            .O(N__11219),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__1600 (
            .O(N__11216),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__1599 (
            .O(N__11213),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    InMux I__1598 (
            .O(N__11204),
            .I(N__11201));
    LocalMux I__1597 (
            .O(N__11201),
            .I(N__11196));
    CascadeMux I__1596 (
            .O(N__11200),
            .I(N__11193));
    InMux I__1595 (
            .O(N__11199),
            .I(N__11190));
    Span4Mux_h I__1594 (
            .O(N__11196),
            .I(N__11187));
    InMux I__1593 (
            .O(N__11193),
            .I(N__11184));
    LocalMux I__1592 (
            .O(N__11190),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    Odrv4 I__1591 (
            .O(N__11187),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__1590 (
            .O(N__11184),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    InMux I__1589 (
            .O(N__11177),
            .I(N__11174));
    LocalMux I__1588 (
            .O(N__11174),
            .I(N__11169));
    InMux I__1587 (
            .O(N__11173),
            .I(N__11165));
    InMux I__1586 (
            .O(N__11172),
            .I(N__11162));
    Span4Mux_h I__1585 (
            .O(N__11169),
            .I(N__11159));
    InMux I__1584 (
            .O(N__11168),
            .I(N__11156));
    LocalMux I__1583 (
            .O(N__11165),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__1582 (
            .O(N__11162),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    Odrv4 I__1581 (
            .O(N__11159),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__1580 (
            .O(N__11156),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    InMux I__1579 (
            .O(N__11147),
            .I(N__11144));
    LocalMux I__1578 (
            .O(N__11144),
            .I(N__11141));
    Span4Mux_v I__1577 (
            .O(N__11141),
            .I(N__11138));
    Odrv4 I__1576 (
            .O(N__11138),
            .I(\transmit_module.video_signal_controller.n21 ));
    InMux I__1575 (
            .O(N__11135),
            .I(N__11131));
    InMux I__1574 (
            .O(N__11134),
            .I(N__11126));
    LocalMux I__1573 (
            .O(N__11131),
            .I(N__11123));
    InMux I__1572 (
            .O(N__11130),
            .I(N__11118));
    InMux I__1571 (
            .O(N__11129),
            .I(N__11118));
    LocalMux I__1570 (
            .O(N__11126),
            .I(\receive_module.rx_counter.Y_4 ));
    Odrv4 I__1569 (
            .O(N__11123),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__1568 (
            .O(N__11118),
            .I(\receive_module.rx_counter.Y_4 ));
    InMux I__1567 (
            .O(N__11111),
            .I(N__11108));
    LocalMux I__1566 (
            .O(N__11108),
            .I(\receive_module.rx_counter.n4 ));
    CascadeMux I__1565 (
            .O(N__11105),
            .I(N__11101));
    InMux I__1564 (
            .O(N__11104),
            .I(N__11097));
    InMux I__1563 (
            .O(N__11101),
            .I(N__11094));
    InMux I__1562 (
            .O(N__11100),
            .I(N__11090));
    LocalMux I__1561 (
            .O(N__11097),
            .I(N__11085));
    LocalMux I__1560 (
            .O(N__11094),
            .I(N__11085));
    InMux I__1559 (
            .O(N__11093),
            .I(N__11082));
    LocalMux I__1558 (
            .O(N__11090),
            .I(\receive_module.rx_counter.Y_3 ));
    Odrv4 I__1557 (
            .O(N__11085),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__1556 (
            .O(N__11082),
            .I(\receive_module.rx_counter.Y_3 ));
    InMux I__1555 (
            .O(N__11075),
            .I(N__11071));
    InMux I__1554 (
            .O(N__11074),
            .I(N__11066));
    LocalMux I__1553 (
            .O(N__11071),
            .I(N__11063));
    InMux I__1552 (
            .O(N__11070),
            .I(N__11058));
    InMux I__1551 (
            .O(N__11069),
            .I(N__11058));
    LocalMux I__1550 (
            .O(N__11066),
            .I(\receive_module.rx_counter.Y_1 ));
    Odrv4 I__1549 (
            .O(N__11063),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__1548 (
            .O(N__11058),
            .I(\receive_module.rx_counter.Y_1 ));
    InMux I__1547 (
            .O(N__11051),
            .I(N__11048));
    LocalMux I__1546 (
            .O(N__11048),
            .I(\receive_module.rx_counter.n3657 ));
    InMux I__1545 (
            .O(N__11045),
            .I(N__11042));
    LocalMux I__1544 (
            .O(N__11042),
            .I(\receive_module.rx_counter.n3619 ));
    CascadeMux I__1543 (
            .O(N__11039),
            .I(\receive_module.rx_counter.n3648_cascade_ ));
    CascadeMux I__1542 (
            .O(N__11036),
            .I(DEBUG_c_5_cascade_));
    SRMux I__1541 (
            .O(N__11033),
            .I(N__11030));
    LocalMux I__1540 (
            .O(N__11030),
            .I(N__11024));
    SRMux I__1539 (
            .O(N__11029),
            .I(N__11021));
    SRMux I__1538 (
            .O(N__11028),
            .I(N__11018));
    SRMux I__1537 (
            .O(N__11027),
            .I(N__11015));
    Span4Mux_v I__1536 (
            .O(N__11024),
            .I(N__11012));
    LocalMux I__1535 (
            .O(N__11021),
            .I(N__11007));
    LocalMux I__1534 (
            .O(N__11018),
            .I(N__11007));
    LocalMux I__1533 (
            .O(N__11015),
            .I(N__11004));
    Sp12to4 I__1532 (
            .O(N__11012),
            .I(N__10999));
    Span12Mux_s6_v I__1531 (
            .O(N__11007),
            .I(N__10999));
    Span4Mux_h I__1530 (
            .O(N__11004),
            .I(N__10996));
    Span12Mux_v I__1529 (
            .O(N__10999),
            .I(N__10993));
    Span4Mux_h I__1528 (
            .O(N__10996),
            .I(N__10990));
    Span12Mux_h I__1527 (
            .O(N__10993),
            .I(N__10987));
    Span4Mux_v I__1526 (
            .O(N__10990),
            .I(N__10984));
    Odrv12 I__1525 (
            .O(N__10987),
            .I(\line_buffer.n641 ));
    Odrv4 I__1524 (
            .O(N__10984),
            .I(\line_buffer.n641 ));
    SRMux I__1523 (
            .O(N__10979),
            .I(N__10974));
    SRMux I__1522 (
            .O(N__10978),
            .I(N__10971));
    SRMux I__1521 (
            .O(N__10977),
            .I(N__10967));
    LocalMux I__1520 (
            .O(N__10974),
            .I(N__10962));
    LocalMux I__1519 (
            .O(N__10971),
            .I(N__10962));
    SRMux I__1518 (
            .O(N__10970),
            .I(N__10959));
    LocalMux I__1517 (
            .O(N__10967),
            .I(N__10956));
    Span4Mux_v I__1516 (
            .O(N__10962),
            .I(N__10951));
    LocalMux I__1515 (
            .O(N__10959),
            .I(N__10951));
    Sp12to4 I__1514 (
            .O(N__10956),
            .I(N__10946));
    Sp12to4 I__1513 (
            .O(N__10951),
            .I(N__10946));
    Span12Mux_v I__1512 (
            .O(N__10946),
            .I(N__10943));
    Span12Mux_h I__1511 (
            .O(N__10943),
            .I(N__10940));
    Odrv12 I__1510 (
            .O(N__10940),
            .I(\line_buffer.n609 ));
    InMux I__1509 (
            .O(N__10937),
            .I(bfn_13_10_0_));
    InMux I__1508 (
            .O(N__10934),
            .I(\receive_module.rx_counter.n3387 ));
    InMux I__1507 (
            .O(N__10931),
            .I(\receive_module.rx_counter.n3388 ));
    InMux I__1506 (
            .O(N__10928),
            .I(\receive_module.rx_counter.n3389 ));
    InMux I__1505 (
            .O(N__10925),
            .I(N__10922));
    LocalMux I__1504 (
            .O(N__10922),
            .I(\transmit_module.n212 ));
    InMux I__1503 (
            .O(N__10919),
            .I(N__10913));
    InMux I__1502 (
            .O(N__10918),
            .I(N__10913));
    LocalMux I__1501 (
            .O(N__10913),
            .I(\transmit_module.n180 ));
    CascadeMux I__1500 (
            .O(N__10910),
            .I(\transmit_module.n212_cascade_ ));
    InMux I__1499 (
            .O(N__10907),
            .I(N__10904));
    LocalMux I__1498 (
            .O(N__10904),
            .I(N__10901));
    Span4Mux_v I__1497 (
            .O(N__10901),
            .I(N__10898));
    Span4Mux_h I__1496 (
            .O(N__10898),
            .I(N__10895));
    Odrv4 I__1495 (
            .O(N__10895),
            .I(\transmit_module.X_DELTA_PATTERN_9 ));
    InMux I__1494 (
            .O(N__10892),
            .I(N__10889));
    LocalMux I__1493 (
            .O(N__10889),
            .I(\transmit_module.X_DELTA_PATTERN_8 ));
    InMux I__1492 (
            .O(N__10886),
            .I(N__10883));
    LocalMux I__1491 (
            .O(N__10883),
            .I(\transmit_module.X_DELTA_PATTERN_7 ));
    InMux I__1490 (
            .O(N__10880),
            .I(N__10877));
    LocalMux I__1489 (
            .O(N__10877),
            .I(\transmit_module.X_DELTA_PATTERN_6 ));
    InMux I__1488 (
            .O(N__10874),
            .I(N__10871));
    LocalMux I__1487 (
            .O(N__10871),
            .I(N__10868));
    Span4Mux_h I__1486 (
            .O(N__10868),
            .I(N__10865));
    Odrv4 I__1485 (
            .O(N__10865),
            .I(\line_buffer.n574 ));
    InMux I__1484 (
            .O(N__10862),
            .I(N__10859));
    LocalMux I__1483 (
            .O(N__10859),
            .I(\line_buffer.n3785 ));
    CascadeMux I__1482 (
            .O(N__10856),
            .I(N__10853));
    InMux I__1481 (
            .O(N__10853),
            .I(N__10850));
    LocalMux I__1480 (
            .O(N__10850),
            .I(N__10847));
    Sp12to4 I__1479 (
            .O(N__10847),
            .I(N__10844));
    Span12Mux_v I__1478 (
            .O(N__10844),
            .I(N__10841));
    Span12Mux_v I__1477 (
            .O(N__10841),
            .I(N__10838));
    Span12Mux_h I__1476 (
            .O(N__10838),
            .I(N__10835));
    Odrv12 I__1475 (
            .O(N__10835),
            .I(\line_buffer.n566 ));
    SRMux I__1474 (
            .O(N__10832),
            .I(N__10828));
    SRMux I__1473 (
            .O(N__10831),
            .I(N__10825));
    LocalMux I__1472 (
            .O(N__10828),
            .I(N__10821));
    LocalMux I__1471 (
            .O(N__10825),
            .I(N__10818));
    SRMux I__1470 (
            .O(N__10824),
            .I(N__10815));
    Span4Mux_h I__1469 (
            .O(N__10821),
            .I(N__10811));
    Span4Mux_v I__1468 (
            .O(N__10818),
            .I(N__10806));
    LocalMux I__1467 (
            .O(N__10815),
            .I(N__10806));
    SRMux I__1466 (
            .O(N__10814),
            .I(N__10803));
    Span4Mux_v I__1465 (
            .O(N__10811),
            .I(N__10800));
    Span4Mux_v I__1464 (
            .O(N__10806),
            .I(N__10797));
    LocalMux I__1463 (
            .O(N__10803),
            .I(N__10794));
    Span4Mux_v I__1462 (
            .O(N__10800),
            .I(N__10787));
    Span4Mux_h I__1461 (
            .O(N__10797),
            .I(N__10787));
    Span4Mux_h I__1460 (
            .O(N__10794),
            .I(N__10787));
    Span4Mux_h I__1459 (
            .O(N__10787),
            .I(N__10784));
    Span4Mux_h I__1458 (
            .O(N__10784),
            .I(N__10781));
    Odrv4 I__1457 (
            .O(N__10781),
            .I(\line_buffer.n577 ));
    SRMux I__1456 (
            .O(N__10778),
            .I(N__10775));
    LocalMux I__1455 (
            .O(N__10775),
            .I(N__10770));
    SRMux I__1454 (
            .O(N__10774),
            .I(N__10767));
    SRMux I__1453 (
            .O(N__10773),
            .I(N__10763));
    Span4Mux_v I__1452 (
            .O(N__10770),
            .I(N__10758));
    LocalMux I__1451 (
            .O(N__10767),
            .I(N__10758));
    SRMux I__1450 (
            .O(N__10766),
            .I(N__10755));
    LocalMux I__1449 (
            .O(N__10763),
            .I(N__10748));
    Sp12to4 I__1448 (
            .O(N__10758),
            .I(N__10748));
    LocalMux I__1447 (
            .O(N__10755),
            .I(N__10748));
    Span12Mux_v I__1446 (
            .O(N__10748),
            .I(N__10745));
    Span12Mux_h I__1445 (
            .O(N__10745),
            .I(N__10742));
    Odrv12 I__1444 (
            .O(N__10742),
            .I(\line_buffer.n513 ));
    InMux I__1443 (
            .O(N__10739),
            .I(N__10733));
    InMux I__1442 (
            .O(N__10738),
            .I(N__10733));
    LocalMux I__1441 (
            .O(N__10733),
            .I(N__10726));
    InMux I__1440 (
            .O(N__10732),
            .I(N__10723));
    InMux I__1439 (
            .O(N__10731),
            .I(N__10720));
    InMux I__1438 (
            .O(N__10730),
            .I(N__10717));
    InMux I__1437 (
            .O(N__10729),
            .I(N__10714));
    Span4Mux_v I__1436 (
            .O(N__10726),
            .I(N__10711));
    LocalMux I__1435 (
            .O(N__10723),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__1434 (
            .O(N__10720),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__1433 (
            .O(N__10717),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__1432 (
            .O(N__10714),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    Odrv4 I__1431 (
            .O(N__10711),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    InMux I__1430 (
            .O(N__10700),
            .I(N__10690));
    InMux I__1429 (
            .O(N__10699),
            .I(N__10690));
    InMux I__1428 (
            .O(N__10698),
            .I(N__10687));
    InMux I__1427 (
            .O(N__10697),
            .I(N__10682));
    InMux I__1426 (
            .O(N__10696),
            .I(N__10682));
    InMux I__1425 (
            .O(N__10695),
            .I(N__10679));
    LocalMux I__1424 (
            .O(N__10690),
            .I(N__10676));
    LocalMux I__1423 (
            .O(N__10687),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    LocalMux I__1422 (
            .O(N__10682),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    LocalMux I__1421 (
            .O(N__10679),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__1420 (
            .O(N__10676),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    InMux I__1419 (
            .O(N__10667),
            .I(N__10664));
    LocalMux I__1418 (
            .O(N__10664),
            .I(\transmit_module.n214 ));
    InMux I__1417 (
            .O(N__10661),
            .I(N__10657));
    InMux I__1416 (
            .O(N__10660),
            .I(N__10654));
    LocalMux I__1415 (
            .O(N__10657),
            .I(\transmit_module.n182 ));
    LocalMux I__1414 (
            .O(N__10654),
            .I(\transmit_module.n182 ));
    CascadeMux I__1413 (
            .O(N__10649),
            .I(\transmit_module.n214_cascade_ ));
    CascadeMux I__1412 (
            .O(N__10646),
            .I(N__10643));
    CascadeBuf I__1411 (
            .O(N__10643),
            .I(N__10639));
    CascadeMux I__1410 (
            .O(N__10642),
            .I(N__10636));
    CascadeMux I__1409 (
            .O(N__10639),
            .I(N__10633));
    CascadeBuf I__1408 (
            .O(N__10636),
            .I(N__10630));
    CascadeBuf I__1407 (
            .O(N__10633),
            .I(N__10627));
    CascadeMux I__1406 (
            .O(N__10630),
            .I(N__10624));
    CascadeMux I__1405 (
            .O(N__10627),
            .I(N__10621));
    CascadeBuf I__1404 (
            .O(N__10624),
            .I(N__10618));
    CascadeBuf I__1403 (
            .O(N__10621),
            .I(N__10615));
    CascadeMux I__1402 (
            .O(N__10618),
            .I(N__10612));
    CascadeMux I__1401 (
            .O(N__10615),
            .I(N__10609));
    CascadeBuf I__1400 (
            .O(N__10612),
            .I(N__10606));
    CascadeBuf I__1399 (
            .O(N__10609),
            .I(N__10603));
    CascadeMux I__1398 (
            .O(N__10606),
            .I(N__10600));
    CascadeMux I__1397 (
            .O(N__10603),
            .I(N__10597));
    CascadeBuf I__1396 (
            .O(N__10600),
            .I(N__10594));
    CascadeBuf I__1395 (
            .O(N__10597),
            .I(N__10591));
    CascadeMux I__1394 (
            .O(N__10594),
            .I(N__10588));
    CascadeMux I__1393 (
            .O(N__10591),
            .I(N__10585));
    CascadeBuf I__1392 (
            .O(N__10588),
            .I(N__10582));
    CascadeBuf I__1391 (
            .O(N__10585),
            .I(N__10579));
    CascadeMux I__1390 (
            .O(N__10582),
            .I(N__10576));
    CascadeMux I__1389 (
            .O(N__10579),
            .I(N__10573));
    CascadeBuf I__1388 (
            .O(N__10576),
            .I(N__10570));
    CascadeBuf I__1387 (
            .O(N__10573),
            .I(N__10567));
    CascadeMux I__1386 (
            .O(N__10570),
            .I(N__10564));
    CascadeMux I__1385 (
            .O(N__10567),
            .I(N__10561));
    CascadeBuf I__1384 (
            .O(N__10564),
            .I(N__10558));
    CascadeBuf I__1383 (
            .O(N__10561),
            .I(N__10555));
    CascadeMux I__1382 (
            .O(N__10558),
            .I(N__10552));
    CascadeMux I__1381 (
            .O(N__10555),
            .I(N__10549));
    CascadeBuf I__1380 (
            .O(N__10552),
            .I(N__10546));
    CascadeBuf I__1379 (
            .O(N__10549),
            .I(N__10543));
    CascadeMux I__1378 (
            .O(N__10546),
            .I(N__10540));
    CascadeMux I__1377 (
            .O(N__10543),
            .I(N__10537));
    CascadeBuf I__1376 (
            .O(N__10540),
            .I(N__10534));
    CascadeBuf I__1375 (
            .O(N__10537),
            .I(N__10531));
    CascadeMux I__1374 (
            .O(N__10534),
            .I(N__10528));
    CascadeMux I__1373 (
            .O(N__10531),
            .I(N__10525));
    CascadeBuf I__1372 (
            .O(N__10528),
            .I(N__10522));
    CascadeBuf I__1371 (
            .O(N__10525),
            .I(N__10519));
    CascadeMux I__1370 (
            .O(N__10522),
            .I(N__10516));
    CascadeMux I__1369 (
            .O(N__10519),
            .I(N__10513));
    CascadeBuf I__1368 (
            .O(N__10516),
            .I(N__10510));
    CascadeBuf I__1367 (
            .O(N__10513),
            .I(N__10507));
    CascadeMux I__1366 (
            .O(N__10510),
            .I(N__10504));
    CascadeMux I__1365 (
            .O(N__10507),
            .I(N__10501));
    CascadeBuf I__1364 (
            .O(N__10504),
            .I(N__10498));
    CascadeBuf I__1363 (
            .O(N__10501),
            .I(N__10495));
    CascadeMux I__1362 (
            .O(N__10498),
            .I(N__10492));
    CascadeMux I__1361 (
            .O(N__10495),
            .I(N__10489));
    CascadeBuf I__1360 (
            .O(N__10492),
            .I(N__10486));
    CascadeBuf I__1359 (
            .O(N__10489),
            .I(N__10483));
    CascadeMux I__1358 (
            .O(N__10486),
            .I(N__10480));
    CascadeMux I__1357 (
            .O(N__10483),
            .I(N__10477));
    CascadeBuf I__1356 (
            .O(N__10480),
            .I(N__10474));
    CascadeBuf I__1355 (
            .O(N__10477),
            .I(N__10471));
    CascadeMux I__1354 (
            .O(N__10474),
            .I(N__10468));
    CascadeMux I__1353 (
            .O(N__10471),
            .I(N__10465));
    CascadeBuf I__1352 (
            .O(N__10468),
            .I(N__10462));
    InMux I__1351 (
            .O(N__10465),
            .I(N__10459));
    CascadeMux I__1350 (
            .O(N__10462),
            .I(N__10456));
    LocalMux I__1349 (
            .O(N__10459),
            .I(N__10453));
    InMux I__1348 (
            .O(N__10456),
            .I(N__10450));
    Span4Mux_v I__1347 (
            .O(N__10453),
            .I(N__10447));
    LocalMux I__1346 (
            .O(N__10450),
            .I(N__10444));
    Span4Mux_h I__1345 (
            .O(N__10447),
            .I(N__10441));
    Span4Mux_h I__1344 (
            .O(N__10444),
            .I(N__10438));
    Sp12to4 I__1343 (
            .O(N__10441),
            .I(N__10435));
    Sp12to4 I__1342 (
            .O(N__10438),
            .I(N__10432));
    Span12Mux_h I__1341 (
            .O(N__10435),
            .I(N__10427));
    Span12Mux_s5_v I__1340 (
            .O(N__10432),
            .I(N__10427));
    Odrv12 I__1339 (
            .O(N__10427),
            .I(n20));
    CascadeMux I__1338 (
            .O(N__10424),
            .I(\transmit_module.n215_cascade_ ));
    CascadeMux I__1337 (
            .O(N__10421),
            .I(N__10417));
    CascadeMux I__1336 (
            .O(N__10420),
            .I(N__10414));
    CascadeBuf I__1335 (
            .O(N__10417),
            .I(N__10411));
    CascadeBuf I__1334 (
            .O(N__10414),
            .I(N__10408));
    CascadeMux I__1333 (
            .O(N__10411),
            .I(N__10405));
    CascadeMux I__1332 (
            .O(N__10408),
            .I(N__10402));
    CascadeBuf I__1331 (
            .O(N__10405),
            .I(N__10399));
    CascadeBuf I__1330 (
            .O(N__10402),
            .I(N__10396));
    CascadeMux I__1329 (
            .O(N__10399),
            .I(N__10393));
    CascadeMux I__1328 (
            .O(N__10396),
            .I(N__10390));
    CascadeBuf I__1327 (
            .O(N__10393),
            .I(N__10387));
    CascadeBuf I__1326 (
            .O(N__10390),
            .I(N__10384));
    CascadeMux I__1325 (
            .O(N__10387),
            .I(N__10381));
    CascadeMux I__1324 (
            .O(N__10384),
            .I(N__10378));
    CascadeBuf I__1323 (
            .O(N__10381),
            .I(N__10375));
    CascadeBuf I__1322 (
            .O(N__10378),
            .I(N__10372));
    CascadeMux I__1321 (
            .O(N__10375),
            .I(N__10369));
    CascadeMux I__1320 (
            .O(N__10372),
            .I(N__10366));
    CascadeBuf I__1319 (
            .O(N__10369),
            .I(N__10363));
    CascadeBuf I__1318 (
            .O(N__10366),
            .I(N__10360));
    CascadeMux I__1317 (
            .O(N__10363),
            .I(N__10357));
    CascadeMux I__1316 (
            .O(N__10360),
            .I(N__10354));
    CascadeBuf I__1315 (
            .O(N__10357),
            .I(N__10351));
    CascadeBuf I__1314 (
            .O(N__10354),
            .I(N__10348));
    CascadeMux I__1313 (
            .O(N__10351),
            .I(N__10345));
    CascadeMux I__1312 (
            .O(N__10348),
            .I(N__10342));
    CascadeBuf I__1311 (
            .O(N__10345),
            .I(N__10339));
    CascadeBuf I__1310 (
            .O(N__10342),
            .I(N__10336));
    CascadeMux I__1309 (
            .O(N__10339),
            .I(N__10333));
    CascadeMux I__1308 (
            .O(N__10336),
            .I(N__10330));
    CascadeBuf I__1307 (
            .O(N__10333),
            .I(N__10327));
    CascadeBuf I__1306 (
            .O(N__10330),
            .I(N__10324));
    CascadeMux I__1305 (
            .O(N__10327),
            .I(N__10321));
    CascadeMux I__1304 (
            .O(N__10324),
            .I(N__10318));
    CascadeBuf I__1303 (
            .O(N__10321),
            .I(N__10315));
    CascadeBuf I__1302 (
            .O(N__10318),
            .I(N__10312));
    CascadeMux I__1301 (
            .O(N__10315),
            .I(N__10309));
    CascadeMux I__1300 (
            .O(N__10312),
            .I(N__10306));
    CascadeBuf I__1299 (
            .O(N__10309),
            .I(N__10303));
    CascadeBuf I__1298 (
            .O(N__10306),
            .I(N__10300));
    CascadeMux I__1297 (
            .O(N__10303),
            .I(N__10297));
    CascadeMux I__1296 (
            .O(N__10300),
            .I(N__10294));
    CascadeBuf I__1295 (
            .O(N__10297),
            .I(N__10291));
    CascadeBuf I__1294 (
            .O(N__10294),
            .I(N__10288));
    CascadeMux I__1293 (
            .O(N__10291),
            .I(N__10285));
    CascadeMux I__1292 (
            .O(N__10288),
            .I(N__10282));
    CascadeBuf I__1291 (
            .O(N__10285),
            .I(N__10279));
    CascadeBuf I__1290 (
            .O(N__10282),
            .I(N__10276));
    CascadeMux I__1289 (
            .O(N__10279),
            .I(N__10273));
    CascadeMux I__1288 (
            .O(N__10276),
            .I(N__10270));
    CascadeBuf I__1287 (
            .O(N__10273),
            .I(N__10267));
    CascadeBuf I__1286 (
            .O(N__10270),
            .I(N__10264));
    CascadeMux I__1285 (
            .O(N__10267),
            .I(N__10261));
    CascadeMux I__1284 (
            .O(N__10264),
            .I(N__10258));
    CascadeBuf I__1283 (
            .O(N__10261),
            .I(N__10255));
    CascadeBuf I__1282 (
            .O(N__10258),
            .I(N__10252));
    CascadeMux I__1281 (
            .O(N__10255),
            .I(N__10249));
    CascadeMux I__1280 (
            .O(N__10252),
            .I(N__10246));
    CascadeBuf I__1279 (
            .O(N__10249),
            .I(N__10243));
    CascadeBuf I__1278 (
            .O(N__10246),
            .I(N__10240));
    CascadeMux I__1277 (
            .O(N__10243),
            .I(N__10237));
    CascadeMux I__1276 (
            .O(N__10240),
            .I(N__10234));
    InMux I__1275 (
            .O(N__10237),
            .I(N__10231));
    InMux I__1274 (
            .O(N__10234),
            .I(N__10228));
    LocalMux I__1273 (
            .O(N__10231),
            .I(N__10225));
    LocalMux I__1272 (
            .O(N__10228),
            .I(N__10222));
    Span12Mux_h I__1271 (
            .O(N__10225),
            .I(N__10219));
    Span4Mux_h I__1270 (
            .O(N__10222),
            .I(N__10216));
    Span12Mux_v I__1269 (
            .O(N__10219),
            .I(N__10213));
    Sp12to4 I__1268 (
            .O(N__10216),
            .I(N__10210));
    Odrv12 I__1267 (
            .O(N__10213),
            .I(n23));
    Odrv12 I__1266 (
            .O(N__10210),
            .I(n23));
    InMux I__1265 (
            .O(N__10205),
            .I(N__10199));
    InMux I__1264 (
            .O(N__10204),
            .I(N__10199));
    LocalMux I__1263 (
            .O(N__10199),
            .I(N__10196));
    Odrv12 I__1262 (
            .O(N__10196),
            .I(\transmit_module.n183 ));
    InMux I__1261 (
            .O(N__10193),
            .I(N__10190));
    LocalMux I__1260 (
            .O(N__10190),
            .I(\transmit_module.n215 ));
    CascadeMux I__1259 (
            .O(N__10187),
            .I(\transmit_module.n3859_cascade_ ));
    InMux I__1258 (
            .O(N__10184),
            .I(N__10179));
    InMux I__1257 (
            .O(N__10183),
            .I(N__10176));
    InMux I__1256 (
            .O(N__10182),
            .I(N__10173));
    LocalMux I__1255 (
            .O(N__10179),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1254 (
            .O(N__10176),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1253 (
            .O(N__10173),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    CascadeMux I__1252 (
            .O(N__10166),
            .I(\transmit_module.video_signal_controller.n4_cascade_ ));
    InMux I__1251 (
            .O(N__10163),
            .I(N__10158));
    InMux I__1250 (
            .O(N__10162),
            .I(N__10155));
    InMux I__1249 (
            .O(N__10161),
            .I(N__10152));
    LocalMux I__1248 (
            .O(N__10158),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1247 (
            .O(N__10155),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1246 (
            .O(N__10152),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    CascadeMux I__1245 (
            .O(N__10145),
            .I(\transmit_module.video_signal_controller.n23_cascade_ ));
    InMux I__1244 (
            .O(N__10142),
            .I(N__10139));
    LocalMux I__1243 (
            .O(N__10139),
            .I(\transmit_module.Y_DELTA_PATTERN_98 ));
    InMux I__1242 (
            .O(N__10136),
            .I(N__10133));
    LocalMux I__1241 (
            .O(N__10133),
            .I(\transmit_module.Y_DELTA_PATTERN_97 ));
    InMux I__1240 (
            .O(N__10130),
            .I(N__10127));
    LocalMux I__1239 (
            .O(N__10127),
            .I(\transmit_module.Y_DELTA_PATTERN_96 ));
    InMux I__1238 (
            .O(N__10124),
            .I(N__10120));
    InMux I__1237 (
            .O(N__10123),
            .I(N__10117));
    LocalMux I__1236 (
            .O(N__10120),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__1235 (
            .O(N__10117),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    InMux I__1234 (
            .O(N__10112),
            .I(N__10108));
    InMux I__1233 (
            .O(N__10111),
            .I(N__10105));
    LocalMux I__1232 (
            .O(N__10108),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__1231 (
            .O(N__10105),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    InMux I__1230 (
            .O(N__10100),
            .I(N__10096));
    InMux I__1229 (
            .O(N__10099),
            .I(N__10093));
    LocalMux I__1228 (
            .O(N__10096),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    LocalMux I__1227 (
            .O(N__10093),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    CascadeMux I__1226 (
            .O(N__10088),
            .I(\transmit_module.video_signal_controller.n8_adj_569_cascade_ ));
    CascadeMux I__1225 (
            .O(N__10085),
            .I(\transmit_module.video_signal_controller.n3029_cascade_ ));
    CascadeMux I__1224 (
            .O(N__10082),
            .I(\transmit_module.video_signal_controller.n3857_cascade_ ));
    CEMux I__1223 (
            .O(N__10079),
            .I(N__10076));
    LocalMux I__1222 (
            .O(N__10076),
            .I(N__10071));
    CEMux I__1221 (
            .O(N__10075),
            .I(N__10068));
    CEMux I__1220 (
            .O(N__10074),
            .I(N__10064));
    Span4Mux_v I__1219 (
            .O(N__10071),
            .I(N__10061));
    LocalMux I__1218 (
            .O(N__10068),
            .I(N__10058));
    CEMux I__1217 (
            .O(N__10067),
            .I(N__10055));
    LocalMux I__1216 (
            .O(N__10064),
            .I(N__10052));
    Odrv4 I__1215 (
            .O(N__10061),
            .I(\transmit_module.n2125 ));
    Odrv4 I__1214 (
            .O(N__10058),
            .I(\transmit_module.n2125 ));
    LocalMux I__1213 (
            .O(N__10055),
            .I(\transmit_module.n2125 ));
    Odrv12 I__1212 (
            .O(N__10052),
            .I(\transmit_module.n2125 ));
    InMux I__1211 (
            .O(N__10043),
            .I(N__10040));
    LocalMux I__1210 (
            .O(N__10040),
            .I(\transmit_module.Y_DELTA_PATTERN_99 ));
    InMux I__1209 (
            .O(N__10037),
            .I(N__10034));
    LocalMux I__1208 (
            .O(N__10034),
            .I(\transmit_module.Y_DELTA_PATTERN_90 ));
    InMux I__1207 (
            .O(N__10031),
            .I(N__10028));
    LocalMux I__1206 (
            .O(N__10028),
            .I(\transmit_module.Y_DELTA_PATTERN_87 ));
    InMux I__1205 (
            .O(N__10025),
            .I(N__10022));
    LocalMux I__1204 (
            .O(N__10022),
            .I(\transmit_module.Y_DELTA_PATTERN_89 ));
    InMux I__1203 (
            .O(N__10019),
            .I(N__10016));
    LocalMux I__1202 (
            .O(N__10016),
            .I(\transmit_module.Y_DELTA_PATTERN_88 ));
    CascadeMux I__1201 (
            .O(N__10013),
            .I(\receive_module.rx_counter.n14_cascade_ ));
    CascadeMux I__1200 (
            .O(N__10010),
            .I(N__10006));
    InMux I__1199 (
            .O(N__10009),
            .I(N__10002));
    InMux I__1198 (
            .O(N__10006),
            .I(N__9997));
    InMux I__1197 (
            .O(N__10005),
            .I(N__9997));
    LocalMux I__1196 (
            .O(N__10002),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__1195 (
            .O(N__9997),
            .I(\receive_module.rx_counter.Y_8 ));
    InMux I__1194 (
            .O(N__9992),
            .I(N__9987));
    InMux I__1193 (
            .O(N__9991),
            .I(N__9982));
    InMux I__1192 (
            .O(N__9990),
            .I(N__9982));
    LocalMux I__1191 (
            .O(N__9987),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__1190 (
            .O(N__9982),
            .I(\receive_module.rx_counter.Y_7 ));
    CascadeMux I__1189 (
            .O(N__9977),
            .I(\receive_module.rx_counter.n15_cascade_ ));
    InMux I__1188 (
            .O(N__9974),
            .I(N__9971));
    LocalMux I__1187 (
            .O(N__9971),
            .I(\receive_module.rx_counter.n3861 ));
    InMux I__1186 (
            .O(N__9968),
            .I(N__9962));
    InMux I__1185 (
            .O(N__9967),
            .I(N__9957));
    InMux I__1184 (
            .O(N__9966),
            .I(N__9957));
    InMux I__1183 (
            .O(N__9965),
            .I(N__9954));
    LocalMux I__1182 (
            .O(N__9962),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__1181 (
            .O(N__9957),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__1180 (
            .O(N__9954),
            .I(\receive_module.rx_counter.Y_0 ));
    InMux I__1179 (
            .O(N__9947),
            .I(N__9944));
    LocalMux I__1178 (
            .O(N__9944),
            .I(\receive_module.rx_counter.n10_adj_570 ));
    InMux I__1177 (
            .O(N__9941),
            .I(N__9935));
    InMux I__1176 (
            .O(N__9940),
            .I(N__9932));
    InMux I__1175 (
            .O(N__9939),
            .I(N__9929));
    InMux I__1174 (
            .O(N__9938),
            .I(N__9926));
    LocalMux I__1173 (
            .O(N__9935),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__1172 (
            .O(N__9932),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__1171 (
            .O(N__9929),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__1170 (
            .O(N__9926),
            .I(\receive_module.rx_counter.Y_2 ));
    SRMux I__1169 (
            .O(N__9917),
            .I(N__9914));
    LocalMux I__1168 (
            .O(N__9914),
            .I(N__9911));
    Span4Mux_v I__1167 (
            .O(N__9911),
            .I(N__9908));
    Span4Mux_v I__1166 (
            .O(N__9908),
            .I(N__9903));
    SRMux I__1165 (
            .O(N__9907),
            .I(N__9900));
    SRMux I__1164 (
            .O(N__9906),
            .I(N__9897));
    Span4Mux_v I__1163 (
            .O(N__9903),
            .I(N__9893));
    LocalMux I__1162 (
            .O(N__9900),
            .I(N__9890));
    LocalMux I__1161 (
            .O(N__9897),
            .I(N__9887));
    SRMux I__1160 (
            .O(N__9896),
            .I(N__9884));
    Span4Mux_v I__1159 (
            .O(N__9893),
            .I(N__9875));
    Span4Mux_v I__1158 (
            .O(N__9890),
            .I(N__9875));
    Span4Mux_v I__1157 (
            .O(N__9887),
            .I(N__9875));
    LocalMux I__1156 (
            .O(N__9884),
            .I(N__9875));
    Span4Mux_h I__1155 (
            .O(N__9875),
            .I(N__9872));
    Odrv4 I__1154 (
            .O(N__9872),
            .I(\line_buffer.n610 ));
    SRMux I__1153 (
            .O(N__9869),
            .I(N__9865));
    SRMux I__1152 (
            .O(N__9868),
            .I(N__9862));
    LocalMux I__1151 (
            .O(N__9865),
            .I(N__9856));
    LocalMux I__1150 (
            .O(N__9862),
            .I(N__9856));
    SRMux I__1149 (
            .O(N__9861),
            .I(N__9853));
    Span4Mux_s3_v I__1148 (
            .O(N__9856),
            .I(N__9847));
    LocalMux I__1147 (
            .O(N__9853),
            .I(N__9847));
    SRMux I__1146 (
            .O(N__9852),
            .I(N__9844));
    Span4Mux_v I__1145 (
            .O(N__9847),
            .I(N__9841));
    LocalMux I__1144 (
            .O(N__9844),
            .I(N__9838));
    Span4Mux_h I__1143 (
            .O(N__9841),
            .I(N__9835));
    Span4Mux_v I__1142 (
            .O(N__9838),
            .I(N__9832));
    Span4Mux_v I__1141 (
            .O(N__9835),
            .I(N__9829));
    Span4Mux_h I__1140 (
            .O(N__9832),
            .I(N__9826));
    Span4Mux_v I__1139 (
            .O(N__9829),
            .I(N__9823));
    Span4Mux_h I__1138 (
            .O(N__9826),
            .I(N__9820));
    Span4Mux_v I__1137 (
            .O(N__9823),
            .I(N__9815));
    Span4Mux_h I__1136 (
            .O(N__9820),
            .I(N__9815));
    Odrv4 I__1135 (
            .O(N__9815),
            .I(\line_buffer.n512 ));
    CascadeMux I__1134 (
            .O(N__9812),
            .I(N__9808));
    CascadeMux I__1133 (
            .O(N__9811),
            .I(N__9805));
    CascadeBuf I__1132 (
            .O(N__9808),
            .I(N__9802));
    CascadeBuf I__1131 (
            .O(N__9805),
            .I(N__9799));
    CascadeMux I__1130 (
            .O(N__9802),
            .I(N__9796));
    CascadeMux I__1129 (
            .O(N__9799),
            .I(N__9793));
    CascadeBuf I__1128 (
            .O(N__9796),
            .I(N__9790));
    CascadeBuf I__1127 (
            .O(N__9793),
            .I(N__9787));
    CascadeMux I__1126 (
            .O(N__9790),
            .I(N__9784));
    CascadeMux I__1125 (
            .O(N__9787),
            .I(N__9781));
    CascadeBuf I__1124 (
            .O(N__9784),
            .I(N__9778));
    CascadeBuf I__1123 (
            .O(N__9781),
            .I(N__9775));
    CascadeMux I__1122 (
            .O(N__9778),
            .I(N__9772));
    CascadeMux I__1121 (
            .O(N__9775),
            .I(N__9769));
    CascadeBuf I__1120 (
            .O(N__9772),
            .I(N__9766));
    CascadeBuf I__1119 (
            .O(N__9769),
            .I(N__9763));
    CascadeMux I__1118 (
            .O(N__9766),
            .I(N__9760));
    CascadeMux I__1117 (
            .O(N__9763),
            .I(N__9757));
    CascadeBuf I__1116 (
            .O(N__9760),
            .I(N__9754));
    CascadeBuf I__1115 (
            .O(N__9757),
            .I(N__9751));
    CascadeMux I__1114 (
            .O(N__9754),
            .I(N__9748));
    CascadeMux I__1113 (
            .O(N__9751),
            .I(N__9745));
    CascadeBuf I__1112 (
            .O(N__9748),
            .I(N__9742));
    CascadeBuf I__1111 (
            .O(N__9745),
            .I(N__9739));
    CascadeMux I__1110 (
            .O(N__9742),
            .I(N__9736));
    CascadeMux I__1109 (
            .O(N__9739),
            .I(N__9733));
    CascadeBuf I__1108 (
            .O(N__9736),
            .I(N__9730));
    CascadeBuf I__1107 (
            .O(N__9733),
            .I(N__9727));
    CascadeMux I__1106 (
            .O(N__9730),
            .I(N__9724));
    CascadeMux I__1105 (
            .O(N__9727),
            .I(N__9721));
    CascadeBuf I__1104 (
            .O(N__9724),
            .I(N__9718));
    CascadeBuf I__1103 (
            .O(N__9721),
            .I(N__9715));
    CascadeMux I__1102 (
            .O(N__9718),
            .I(N__9712));
    CascadeMux I__1101 (
            .O(N__9715),
            .I(N__9709));
    CascadeBuf I__1100 (
            .O(N__9712),
            .I(N__9706));
    CascadeBuf I__1099 (
            .O(N__9709),
            .I(N__9703));
    CascadeMux I__1098 (
            .O(N__9706),
            .I(N__9700));
    CascadeMux I__1097 (
            .O(N__9703),
            .I(N__9697));
    CascadeBuf I__1096 (
            .O(N__9700),
            .I(N__9694));
    CascadeBuf I__1095 (
            .O(N__9697),
            .I(N__9691));
    CascadeMux I__1094 (
            .O(N__9694),
            .I(N__9688));
    CascadeMux I__1093 (
            .O(N__9691),
            .I(N__9685));
    CascadeBuf I__1092 (
            .O(N__9688),
            .I(N__9682));
    CascadeBuf I__1091 (
            .O(N__9685),
            .I(N__9679));
    CascadeMux I__1090 (
            .O(N__9682),
            .I(N__9676));
    CascadeMux I__1089 (
            .O(N__9679),
            .I(N__9673));
    CascadeBuf I__1088 (
            .O(N__9676),
            .I(N__9670));
    CascadeBuf I__1087 (
            .O(N__9673),
            .I(N__9667));
    CascadeMux I__1086 (
            .O(N__9670),
            .I(N__9664));
    CascadeMux I__1085 (
            .O(N__9667),
            .I(N__9661));
    CascadeBuf I__1084 (
            .O(N__9664),
            .I(N__9658));
    CascadeBuf I__1083 (
            .O(N__9661),
            .I(N__9655));
    CascadeMux I__1082 (
            .O(N__9658),
            .I(N__9652));
    CascadeMux I__1081 (
            .O(N__9655),
            .I(N__9649));
    CascadeBuf I__1080 (
            .O(N__9652),
            .I(N__9646));
    CascadeBuf I__1079 (
            .O(N__9649),
            .I(N__9643));
    CascadeMux I__1078 (
            .O(N__9646),
            .I(N__9640));
    CascadeMux I__1077 (
            .O(N__9643),
            .I(N__9637));
    CascadeBuf I__1076 (
            .O(N__9640),
            .I(N__9634));
    CascadeBuf I__1075 (
            .O(N__9637),
            .I(N__9631));
    CascadeMux I__1074 (
            .O(N__9634),
            .I(N__9628));
    CascadeMux I__1073 (
            .O(N__9631),
            .I(N__9625));
    InMux I__1072 (
            .O(N__9628),
            .I(N__9622));
    InMux I__1071 (
            .O(N__9625),
            .I(N__9619));
    LocalMux I__1070 (
            .O(N__9622),
            .I(N__9616));
    LocalMux I__1069 (
            .O(N__9619),
            .I(N__9613));
    Span12Mux_h I__1068 (
            .O(N__9616),
            .I(N__9610));
    Span12Mux_h I__1067 (
            .O(N__9613),
            .I(N__9607));
    Span12Mux_v I__1066 (
            .O(N__9610),
            .I(N__9602));
    Span12Mux_v I__1065 (
            .O(N__9607),
            .I(N__9602));
    Odrv12 I__1064 (
            .O(N__9602),
            .I(n22));
    InMux I__1063 (
            .O(N__9599),
            .I(N__9596));
    LocalMux I__1062 (
            .O(N__9596),
            .I(\transmit_module.X_DELTA_PATTERN_15 ));
    InMux I__1061 (
            .O(N__9593),
            .I(N__9590));
    LocalMux I__1060 (
            .O(N__9590),
            .I(\transmit_module.X_DELTA_PATTERN_14 ));
    InMux I__1059 (
            .O(N__9587),
            .I(N__9584));
    LocalMux I__1058 (
            .O(N__9584),
            .I(N__9581));
    Span4Mux_v I__1057 (
            .O(N__9581),
            .I(N__9578));
    Span4Mux_h I__1056 (
            .O(N__9578),
            .I(N__9575));
    Odrv4 I__1055 (
            .O(N__9575),
            .I(\line_buffer.n630 ));
    CascadeMux I__1054 (
            .O(N__9572),
            .I(N__9569));
    InMux I__1053 (
            .O(N__9569),
            .I(N__9566));
    LocalMux I__1052 (
            .O(N__9566),
            .I(N__9563));
    Span4Mux_h I__1051 (
            .O(N__9563),
            .I(N__9560));
    Span4Mux_v I__1050 (
            .O(N__9560),
            .I(N__9557));
    Odrv4 I__1049 (
            .O(N__9557),
            .I(\line_buffer.n638 ));
    InMux I__1048 (
            .O(N__9554),
            .I(N__9549));
    InMux I__1047 (
            .O(N__9553),
            .I(N__9544));
    InMux I__1046 (
            .O(N__9552),
            .I(N__9544));
    LocalMux I__1045 (
            .O(N__9549),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__1044 (
            .O(N__9544),
            .I(\receive_module.rx_counter.Y_6 ));
    InMux I__1043 (
            .O(N__9539),
            .I(N__9534));
    InMux I__1042 (
            .O(N__9538),
            .I(N__9531));
    InMux I__1041 (
            .O(N__9537),
            .I(N__9528));
    LocalMux I__1040 (
            .O(N__9534),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__1039 (
            .O(N__9531),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__1038 (
            .O(N__9528),
            .I(\receive_module.rx_counter.Y_5 ));
    CascadeMux I__1037 (
            .O(N__9521),
            .I(\receive_module.rx_counter.n3619_cascade_ ));
    SRMux I__1036 (
            .O(N__9518),
            .I(N__9515));
    LocalMux I__1035 (
            .O(N__9515),
            .I(N__9511));
    SRMux I__1034 (
            .O(N__9514),
            .I(N__9508));
    Span4Mux_v I__1033 (
            .O(N__9511),
            .I(N__9502));
    LocalMux I__1032 (
            .O(N__9508),
            .I(N__9502));
    SRMux I__1031 (
            .O(N__9507),
            .I(N__9499));
    Span4Mux_v I__1030 (
            .O(N__9502),
            .I(N__9493));
    LocalMux I__1029 (
            .O(N__9499),
            .I(N__9493));
    SRMux I__1028 (
            .O(N__9498),
            .I(N__9490));
    Span4Mux_v I__1027 (
            .O(N__9493),
            .I(N__9485));
    LocalMux I__1026 (
            .O(N__9490),
            .I(N__9485));
    Span4Mux_h I__1025 (
            .O(N__9485),
            .I(N__9482));
    Span4Mux_v I__1024 (
            .O(N__9482),
            .I(N__9479));
    Odrv4 I__1023 (
            .O(N__9479),
            .I(\line_buffer.n642 ));
    SRMux I__1022 (
            .O(N__9476),
            .I(N__9472));
    SRMux I__1021 (
            .O(N__9475),
            .I(N__9469));
    LocalMux I__1020 (
            .O(N__9472),
            .I(N__9465));
    LocalMux I__1019 (
            .O(N__9469),
            .I(N__9462));
    SRMux I__1018 (
            .O(N__9468),
            .I(N__9459));
    Span4Mux_v I__1017 (
            .O(N__9465),
            .I(N__9455));
    Span4Mux_s3_v I__1016 (
            .O(N__9462),
            .I(N__9450));
    LocalMux I__1015 (
            .O(N__9459),
            .I(N__9450));
    SRMux I__1014 (
            .O(N__9458),
            .I(N__9447));
    Span4Mux_h I__1013 (
            .O(N__9455),
            .I(N__9444));
    Span4Mux_h I__1012 (
            .O(N__9450),
            .I(N__9439));
    LocalMux I__1011 (
            .O(N__9447),
            .I(N__9439));
    Span4Mux_v I__1010 (
            .O(N__9444),
            .I(N__9436));
    Span4Mux_v I__1009 (
            .O(N__9439),
            .I(N__9433));
    Span4Mux_v I__1008 (
            .O(N__9436),
            .I(N__9428));
    Span4Mux_h I__1007 (
            .O(N__9433),
            .I(N__9428));
    Odrv4 I__1006 (
            .O(N__9428),
            .I(\line_buffer.n578 ));
    InMux I__1005 (
            .O(N__9425),
            .I(bfn_11_16_0_));
    InMux I__1004 (
            .O(N__9422),
            .I(\transmit_module.video_signal_controller.n3385 ));
    InMux I__1003 (
            .O(N__9419),
            .I(\transmit_module.video_signal_controller.n3386 ));
    InMux I__1002 (
            .O(N__9416),
            .I(N__9413));
    LocalMux I__1001 (
            .O(N__9413),
            .I(N__9410));
    Odrv12 I__1000 (
            .O(N__9410),
            .I(\transmit_module.Y_DELTA_PATTERN_28 ));
    InMux I__999 (
            .O(N__9407),
            .I(N__9404));
    LocalMux I__998 (
            .O(N__9404),
            .I(\transmit_module.Y_DELTA_PATTERN_29 ));
    InMux I__997 (
            .O(N__9401),
            .I(N__9398));
    LocalMux I__996 (
            .O(N__9398),
            .I(\transmit_module.Y_DELTA_PATTERN_30 ));
    InMux I__995 (
            .O(N__9395),
            .I(N__9392));
    LocalMux I__994 (
            .O(N__9392),
            .I(\transmit_module.Y_DELTA_PATTERN_31 ));
    InMux I__993 (
            .O(N__9389),
            .I(N__9386));
    LocalMux I__992 (
            .O(N__9386),
            .I(\transmit_module.Y_DELTA_PATTERN_73 ));
    InMux I__991 (
            .O(N__9383),
            .I(N__9380));
    LocalMux I__990 (
            .O(N__9380),
            .I(N__9377));
    Span4Mux_h I__989 (
            .O(N__9377),
            .I(N__9374));
    Odrv4 I__988 (
            .O(N__9374),
            .I(\transmit_module.Y_DELTA_PATTERN_72 ));
    InMux I__987 (
            .O(N__9371),
            .I(N__9368));
    LocalMux I__986 (
            .O(N__9368),
            .I(\transmit_module.Y_DELTA_PATTERN_92 ));
    InMux I__985 (
            .O(N__9365),
            .I(N__9362));
    LocalMux I__984 (
            .O(N__9362),
            .I(\transmit_module.Y_DELTA_PATTERN_91 ));
    InMux I__983 (
            .O(N__9359),
            .I(bfn_11_15_0_));
    InMux I__982 (
            .O(N__9356),
            .I(\transmit_module.video_signal_controller.n3377 ));
    InMux I__981 (
            .O(N__9353),
            .I(\transmit_module.video_signal_controller.n3378 ));
    InMux I__980 (
            .O(N__9350),
            .I(\transmit_module.video_signal_controller.n3379 ));
    InMux I__979 (
            .O(N__9347),
            .I(\transmit_module.video_signal_controller.n3380 ));
    InMux I__978 (
            .O(N__9344),
            .I(\transmit_module.video_signal_controller.n3381 ));
    InMux I__977 (
            .O(N__9341),
            .I(\transmit_module.video_signal_controller.n3382 ));
    InMux I__976 (
            .O(N__9338),
            .I(\transmit_module.video_signal_controller.n3383 ));
    InMux I__975 (
            .O(N__9335),
            .I(N__9332));
    LocalMux I__974 (
            .O(N__9332),
            .I(\transmit_module.Y_DELTA_PATTERN_12 ));
    InMux I__973 (
            .O(N__9329),
            .I(N__9326));
    LocalMux I__972 (
            .O(N__9326),
            .I(\transmit_module.Y_DELTA_PATTERN_11 ));
    InMux I__971 (
            .O(N__9323),
            .I(N__9320));
    LocalMux I__970 (
            .O(N__9320),
            .I(N__9317));
    Span4Mux_h I__969 (
            .O(N__9317),
            .I(N__9314));
    Odrv4 I__968 (
            .O(N__9314),
            .I(\transmit_module.Y_DELTA_PATTERN_83 ));
    InMux I__967 (
            .O(N__9311),
            .I(N__9308));
    LocalMux I__966 (
            .O(N__9308),
            .I(\transmit_module.Y_DELTA_PATTERN_84 ));
    InMux I__965 (
            .O(N__9305),
            .I(N__9302));
    LocalMux I__964 (
            .O(N__9302),
            .I(\transmit_module.Y_DELTA_PATTERN_95 ));
    InMux I__963 (
            .O(N__9299),
            .I(N__9296));
    LocalMux I__962 (
            .O(N__9296),
            .I(\transmit_module.Y_DELTA_PATTERN_94 ));
    InMux I__961 (
            .O(N__9293),
            .I(N__9290));
    LocalMux I__960 (
            .O(N__9290),
            .I(\transmit_module.Y_DELTA_PATTERN_93 ));
    InMux I__959 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__958 (
            .O(N__9284),
            .I(\transmit_module.Y_DELTA_PATTERN_85 ));
    InMux I__957 (
            .O(N__9281),
            .I(N__9278));
    LocalMux I__956 (
            .O(N__9278),
            .I(\transmit_module.Y_DELTA_PATTERN_86 ));
    InMux I__955 (
            .O(N__9275),
            .I(N__9272));
    LocalMux I__954 (
            .O(N__9272),
            .I(\transmit_module.Y_DELTA_PATTERN_26 ));
    InMux I__953 (
            .O(N__9269),
            .I(N__9266));
    LocalMux I__952 (
            .O(N__9266),
            .I(\transmit_module.Y_DELTA_PATTERN_25 ));
    InMux I__951 (
            .O(N__9263),
            .I(N__9260));
    LocalMux I__950 (
            .O(N__9260),
            .I(\transmit_module.Y_DELTA_PATTERN_7 ));
    InMux I__949 (
            .O(N__9257),
            .I(N__9254));
    LocalMux I__948 (
            .O(N__9254),
            .I(\transmit_module.Y_DELTA_PATTERN_27 ));
    InMux I__947 (
            .O(N__9251),
            .I(N__9248));
    LocalMux I__946 (
            .O(N__9248),
            .I(\transmit_module.Y_DELTA_PATTERN_10 ));
    InMux I__945 (
            .O(N__9245),
            .I(N__9242));
    LocalMux I__944 (
            .O(N__9242),
            .I(N__9239));
    Span4Mux_h I__943 (
            .O(N__9239),
            .I(N__9236));
    Odrv4 I__942 (
            .O(N__9236),
            .I(\transmit_module.Y_DELTA_PATTERN_13 ));
    InMux I__941 (
            .O(N__9233),
            .I(N__9230));
    LocalMux I__940 (
            .O(N__9230),
            .I(\transmit_module.Y_DELTA_PATTERN_9 ));
    InMux I__939 (
            .O(N__9227),
            .I(N__9224));
    LocalMux I__938 (
            .O(N__9224),
            .I(\transmit_module.Y_DELTA_PATTERN_8 ));
    InMux I__937 (
            .O(N__9221),
            .I(bfn_11_9_0_));
    InMux I__936 (
            .O(N__9218),
            .I(\receive_module.rx_counter.n3349 ));
    InMux I__935 (
            .O(N__9215),
            .I(\receive_module.rx_counter.n3350 ));
    InMux I__934 (
            .O(N__9212),
            .I(\receive_module.rx_counter.n3351 ));
    InMux I__933 (
            .O(N__9209),
            .I(\receive_module.rx_counter.n3352 ));
    InMux I__932 (
            .O(N__9206),
            .I(\receive_module.rx_counter.n3353 ));
    InMux I__931 (
            .O(N__9203),
            .I(\receive_module.rx_counter.n3354 ));
    InMux I__930 (
            .O(N__9200),
            .I(\receive_module.rx_counter.n3355 ));
    InMux I__929 (
            .O(N__9197),
            .I(bfn_11_10_0_));
    CEMux I__928 (
            .O(N__9194),
            .I(N__9191));
    LocalMux I__927 (
            .O(N__9191),
            .I(N__9187));
    CEMux I__926 (
            .O(N__9190),
            .I(N__9184));
    Sp12to4 I__925 (
            .O(N__9187),
            .I(N__9179));
    LocalMux I__924 (
            .O(N__9184),
            .I(N__9179));
    Odrv12 I__923 (
            .O(N__9179),
            .I(n2057));
    InMux I__922 (
            .O(N__9176),
            .I(N__9173));
    LocalMux I__921 (
            .O(N__9173),
            .I(N__9170));
    Odrv12 I__920 (
            .O(N__9170),
            .I(\transmit_module.Y_DELTA_PATTERN_51 ));
    InMux I__919 (
            .O(N__9167),
            .I(N__9164));
    LocalMux I__918 (
            .O(N__9164),
            .I(N__9161));
    Odrv4 I__917 (
            .O(N__9161),
            .I(\transmit_module.Y_DELTA_PATTERN_63 ));
    InMux I__916 (
            .O(N__9158),
            .I(N__9155));
    LocalMux I__915 (
            .O(N__9155),
            .I(\transmit_module.Y_DELTA_PATTERN_62 ));
    InMux I__914 (
            .O(N__9152),
            .I(N__9149));
    LocalMux I__913 (
            .O(N__9149),
            .I(\transmit_module.Y_DELTA_PATTERN_74 ));
    InMux I__912 (
            .O(N__9146),
            .I(N__9143));
    LocalMux I__911 (
            .O(N__9143),
            .I(\transmit_module.Y_DELTA_PATTERN_50 ));
    InMux I__910 (
            .O(N__9140),
            .I(N__9137));
    LocalMux I__909 (
            .O(N__9137),
            .I(\transmit_module.Y_DELTA_PATTERN_49 ));
    InMux I__908 (
            .O(N__9134),
            .I(N__9131));
    LocalMux I__907 (
            .O(N__9131),
            .I(\transmit_module.Y_DELTA_PATTERN_65 ));
    InMux I__906 (
            .O(N__9128),
            .I(N__9125));
    LocalMux I__905 (
            .O(N__9125),
            .I(N__9122));
    Odrv4 I__904 (
            .O(N__9122),
            .I(\transmit_module.Y_DELTA_PATTERN_64 ));
    InMux I__903 (
            .O(N__9119),
            .I(N__9116));
    LocalMux I__902 (
            .O(N__9116),
            .I(\transmit_module.X_DELTA_PATTERN_12 ));
    InMux I__901 (
            .O(N__9113),
            .I(N__9110));
    LocalMux I__900 (
            .O(N__9110),
            .I(\transmit_module.X_DELTA_PATTERN_13 ));
    InMux I__899 (
            .O(N__9107),
            .I(N__9104));
    LocalMux I__898 (
            .O(N__9104),
            .I(old_HS));
    InMux I__897 (
            .O(N__9101),
            .I(N__9098));
    LocalMux I__896 (
            .O(N__9098),
            .I(\transmit_module.Y_DELTA_PATTERN_79 ));
    InMux I__895 (
            .O(N__9095),
            .I(N__9092));
    LocalMux I__894 (
            .O(N__9092),
            .I(N__9089));
    Odrv4 I__893 (
            .O(N__9089),
            .I(\transmit_module.Y_DELTA_PATTERN_48 ));
    InMux I__892 (
            .O(N__9086),
            .I(N__9083));
    LocalMux I__891 (
            .O(N__9083),
            .I(\transmit_module.Y_DELTA_PATTERN_47 ));
    InMux I__890 (
            .O(N__9080),
            .I(N__9077));
    LocalMux I__889 (
            .O(N__9077),
            .I(\transmit_module.Y_DELTA_PATTERN_67 ));
    InMux I__888 (
            .O(N__9074),
            .I(N__9071));
    LocalMux I__887 (
            .O(N__9071),
            .I(\transmit_module.Y_DELTA_PATTERN_82 ));
    InMux I__886 (
            .O(N__9068),
            .I(N__9065));
    LocalMux I__885 (
            .O(N__9065),
            .I(\transmit_module.Y_DELTA_PATTERN_44 ));
    InMux I__884 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__883 (
            .O(N__9059),
            .I(\transmit_module.Y_DELTA_PATTERN_43 ));
    InMux I__882 (
            .O(N__9056),
            .I(N__9053));
    LocalMux I__881 (
            .O(N__9053),
            .I(\transmit_module.Y_DELTA_PATTERN_81 ));
    InMux I__880 (
            .O(N__9050),
            .I(N__9047));
    LocalMux I__879 (
            .O(N__9047),
            .I(\transmit_module.Y_DELTA_PATTERN_80 ));
    InMux I__878 (
            .O(N__9044),
            .I(N__9041));
    LocalMux I__877 (
            .O(N__9041),
            .I(\transmit_module.Y_DELTA_PATTERN_66 ));
    InMux I__876 (
            .O(N__9038),
            .I(N__9035));
    LocalMux I__875 (
            .O(N__9035),
            .I(N__9032));
    Odrv4 I__874 (
            .O(N__9032),
            .I(\transmit_module.Y_DELTA_PATTERN_76 ));
    InMux I__873 (
            .O(N__9029),
            .I(N__9026));
    LocalMux I__872 (
            .O(N__9026),
            .I(\transmit_module.Y_DELTA_PATTERN_75 ));
    InMux I__871 (
            .O(N__9023),
            .I(N__9020));
    LocalMux I__870 (
            .O(N__9020),
            .I(\transmit_module.Y_DELTA_PATTERN_45 ));
    InMux I__869 (
            .O(N__9017),
            .I(N__9014));
    LocalMux I__868 (
            .O(N__9014),
            .I(\transmit_module.Y_DELTA_PATTERN_77 ));
    InMux I__867 (
            .O(N__9011),
            .I(N__9008));
    LocalMux I__866 (
            .O(N__9008),
            .I(\transmit_module.Y_DELTA_PATTERN_3 ));
    InMux I__865 (
            .O(N__9005),
            .I(N__9002));
    LocalMux I__864 (
            .O(N__9002),
            .I(\transmit_module.Y_DELTA_PATTERN_2 ));
    InMux I__863 (
            .O(N__8999),
            .I(N__8996));
    LocalMux I__862 (
            .O(N__8996),
            .I(\transmit_module.Y_DELTA_PATTERN_46 ));
    InMux I__861 (
            .O(N__8993),
            .I(N__8990));
    LocalMux I__860 (
            .O(N__8990),
            .I(\transmit_module.Y_DELTA_PATTERN_78 ));
    InMux I__859 (
            .O(N__8987),
            .I(N__8984));
    LocalMux I__858 (
            .O(N__8984),
            .I(\transmit_module.Y_DELTA_PATTERN_68 ));
    InMux I__857 (
            .O(N__8981),
            .I(N__8978));
    LocalMux I__856 (
            .O(N__8978),
            .I(\transmit_module.Y_DELTA_PATTERN_6 ));
    InMux I__855 (
            .O(N__8975),
            .I(N__8972));
    LocalMux I__854 (
            .O(N__8972),
            .I(\transmit_module.Y_DELTA_PATTERN_20 ));
    InMux I__853 (
            .O(N__8969),
            .I(N__8966));
    LocalMux I__852 (
            .O(N__8966),
            .I(\transmit_module.Y_DELTA_PATTERN_21 ));
    InMux I__851 (
            .O(N__8963),
            .I(N__8960));
    LocalMux I__850 (
            .O(N__8960),
            .I(N__8957));
    Odrv4 I__849 (
            .O(N__8957),
            .I(\transmit_module.Y_DELTA_PATTERN_23 ));
    InMux I__848 (
            .O(N__8954),
            .I(N__8951));
    LocalMux I__847 (
            .O(N__8951),
            .I(\transmit_module.Y_DELTA_PATTERN_22 ));
    InMux I__846 (
            .O(N__8948),
            .I(N__8945));
    LocalMux I__845 (
            .O(N__8945),
            .I(N__8942));
    Odrv4 I__844 (
            .O(N__8942),
            .I(\transmit_module.Y_DELTA_PATTERN_5 ));
    InMux I__843 (
            .O(N__8939),
            .I(N__8936));
    LocalMux I__842 (
            .O(N__8936),
            .I(\transmit_module.Y_DELTA_PATTERN_1 ));
    InMux I__841 (
            .O(N__8933),
            .I(N__8930));
    LocalMux I__840 (
            .O(N__8930),
            .I(\transmit_module.Y_DELTA_PATTERN_4 ));
    InMux I__839 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__838 (
            .O(N__8924),
            .I(\transmit_module.Y_DELTA_PATTERN_69 ));
    InMux I__837 (
            .O(N__8921),
            .I(N__8918));
    LocalMux I__836 (
            .O(N__8918),
            .I(N__8915));
    Span4Mux_h I__835 (
            .O(N__8915),
            .I(N__8912));
    Odrv4 I__834 (
            .O(N__8912),
            .I(\transmit_module.Y_DELTA_PATTERN_56 ));
    InMux I__833 (
            .O(N__8909),
            .I(N__8906));
    LocalMux I__832 (
            .O(N__8906),
            .I(\transmit_module.Y_DELTA_PATTERN_58 ));
    InMux I__831 (
            .O(N__8903),
            .I(N__8900));
    LocalMux I__830 (
            .O(N__8900),
            .I(\transmit_module.Y_DELTA_PATTERN_57 ));
    InMux I__829 (
            .O(N__8897),
            .I(N__8894));
    LocalMux I__828 (
            .O(N__8894),
            .I(\transmit_module.Y_DELTA_PATTERN_61 ));
    InMux I__827 (
            .O(N__8891),
            .I(N__8888));
    LocalMux I__826 (
            .O(N__8888),
            .I(N__8885));
    Span4Mux_v I__825 (
            .O(N__8885),
            .I(N__8882));
    Odrv4 I__824 (
            .O(N__8882),
            .I(\line_buffer.n639 ));
    InMux I__823 (
            .O(N__8879),
            .I(N__8876));
    LocalMux I__822 (
            .O(N__8876),
            .I(N__8873));
    Odrv4 I__821 (
            .O(N__8873),
            .I(\line_buffer.n631 ));
    InMux I__820 (
            .O(N__8870),
            .I(N__8867));
    LocalMux I__819 (
            .O(N__8867),
            .I(\transmit_module.X_DELTA_PATTERN_11 ));
    InMux I__818 (
            .O(N__8864),
            .I(N__8861));
    LocalMux I__817 (
            .O(N__8861),
            .I(N__8858));
    Odrv4 I__816 (
            .O(N__8858),
            .I(\transmit_module.X_DELTA_PATTERN_10 ));
    InMux I__815 (
            .O(N__8855),
            .I(N__8852));
    LocalMux I__814 (
            .O(N__8852),
            .I(\transmit_module.Y_DELTA_PATTERN_24 ));
    InMux I__813 (
            .O(N__8849),
            .I(N__8846));
    LocalMux I__812 (
            .O(N__8846),
            .I(\transmit_module.Y_DELTA_PATTERN_71 ));
    InMux I__811 (
            .O(N__8843),
            .I(N__8840));
    LocalMux I__810 (
            .O(N__8840),
            .I(\transmit_module.Y_DELTA_PATTERN_70 ));
    InMux I__809 (
            .O(N__8837),
            .I(N__8834));
    LocalMux I__808 (
            .O(N__8834),
            .I(\transmit_module.Y_DELTA_PATTERN_60 ));
    InMux I__807 (
            .O(N__8831),
            .I(N__8828));
    LocalMux I__806 (
            .O(N__8828),
            .I(\transmit_module.Y_DELTA_PATTERN_59 ));
    InMux I__805 (
            .O(N__8825),
            .I(N__8822));
    LocalMux I__804 (
            .O(N__8822),
            .I(\transmit_module.Y_DELTA_PATTERN_42 ));
    InMux I__803 (
            .O(N__8819),
            .I(N__8816));
    LocalMux I__802 (
            .O(N__8816),
            .I(\transmit_module.Y_DELTA_PATTERN_41 ));
    InMux I__801 (
            .O(N__8813),
            .I(N__8810));
    LocalMux I__800 (
            .O(N__8810),
            .I(\transmit_module.Y_DELTA_PATTERN_14 ));
    InMux I__799 (
            .O(N__8807),
            .I(N__8804));
    LocalMux I__798 (
            .O(N__8804),
            .I(\transmit_module.Y_DELTA_PATTERN_15 ));
    InMux I__797 (
            .O(N__8801),
            .I(N__8798));
    LocalMux I__796 (
            .O(N__8798),
            .I(\transmit_module.Y_DELTA_PATTERN_16 ));
    InMux I__795 (
            .O(N__8795),
            .I(N__8792));
    LocalMux I__794 (
            .O(N__8792),
            .I(\transmit_module.Y_DELTA_PATTERN_17 ));
    InMux I__793 (
            .O(N__8789),
            .I(N__8786));
    LocalMux I__792 (
            .O(N__8786),
            .I(\transmit_module.Y_DELTA_PATTERN_19 ));
    InMux I__791 (
            .O(N__8783),
            .I(N__8780));
    LocalMux I__790 (
            .O(N__8780),
            .I(\transmit_module.Y_DELTA_PATTERN_18 ));
    InMux I__789 (
            .O(N__8777),
            .I(N__8774));
    LocalMux I__788 (
            .O(N__8774),
            .I(N__8771));
    Span4Mux_s2_v I__787 (
            .O(N__8771),
            .I(N__8767));
    InMux I__786 (
            .O(N__8770),
            .I(N__8764));
    Span4Mux_v I__785 (
            .O(N__8767),
            .I(N__8759));
    LocalMux I__784 (
            .O(N__8764),
            .I(N__8759));
    Span4Mux_v I__783 (
            .O(N__8759),
            .I(N__8755));
    InMux I__782 (
            .O(N__8758),
            .I(N__8752));
    Span4Mux_v I__781 (
            .O(N__8755),
            .I(N__8746));
    LocalMux I__780 (
            .O(N__8752),
            .I(N__8746));
    InMux I__779 (
            .O(N__8751),
            .I(N__8743));
    Span4Mux_v I__778 (
            .O(N__8746),
            .I(N__8738));
    LocalMux I__777 (
            .O(N__8743),
            .I(N__8738));
    Span4Mux_v I__776 (
            .O(N__8738),
            .I(N__8733));
    InMux I__775 (
            .O(N__8737),
            .I(N__8730));
    InMux I__774 (
            .O(N__8736),
            .I(N__8727));
    Span4Mux_v I__773 (
            .O(N__8733),
            .I(N__8722));
    LocalMux I__772 (
            .O(N__8730),
            .I(N__8722));
    LocalMux I__771 (
            .O(N__8727),
            .I(N__8719));
    Span4Mux_h I__770 (
            .O(N__8722),
            .I(N__8715));
    Span4Mux_h I__769 (
            .O(N__8719),
            .I(N__8712));
    InMux I__768 (
            .O(N__8718),
            .I(N__8709));
    Span4Mux_h I__767 (
            .O(N__8715),
            .I(N__8706));
    Span4Mux_v I__766 (
            .O(N__8712),
            .I(N__8702));
    LocalMux I__765 (
            .O(N__8709),
            .I(N__8699));
    Span4Mux_h I__764 (
            .O(N__8706),
            .I(N__8696));
    InMux I__763 (
            .O(N__8705),
            .I(N__8693));
    Span4Mux_v I__762 (
            .O(N__8702),
            .I(N__8688));
    Span4Mux_h I__761 (
            .O(N__8699),
            .I(N__8688));
    Span4Mux_h I__760 (
            .O(N__8696),
            .I(N__8683));
    LocalMux I__759 (
            .O(N__8693),
            .I(N__8683));
    Span4Mux_v I__758 (
            .O(N__8688),
            .I(N__8680));
    Span4Mux_h I__757 (
            .O(N__8683),
            .I(N__8677));
    Span4Mux_v I__756 (
            .O(N__8680),
            .I(N__8674));
    Span4Mux_v I__755 (
            .O(N__8677),
            .I(N__8671));
    Odrv4 I__754 (
            .O(N__8674),
            .I(TVP_VIDEO_c_2));
    Odrv4 I__753 (
            .O(N__8671),
            .I(TVP_VIDEO_c_2));
    InMux I__752 (
            .O(N__8666),
            .I(N__8663));
    LocalMux I__751 (
            .O(N__8663),
            .I(\transmit_module.Y_DELTA_PATTERN_55 ));
    InMux I__750 (
            .O(N__8660),
            .I(N__8657));
    LocalMux I__749 (
            .O(N__8657),
            .I(\transmit_module.Y_DELTA_PATTERN_54 ));
    InMux I__748 (
            .O(N__8654),
            .I(N__8651));
    LocalMux I__747 (
            .O(N__8651),
            .I(\transmit_module.Y_DELTA_PATTERN_53 ));
    InMux I__746 (
            .O(N__8648),
            .I(N__8645));
    LocalMux I__745 (
            .O(N__8645),
            .I(\transmit_module.Y_DELTA_PATTERN_52 ));
    InMux I__744 (
            .O(N__8642),
            .I(N__8639));
    LocalMux I__743 (
            .O(N__8639),
            .I(N__8633));
    InMux I__742 (
            .O(N__8638),
            .I(N__8630));
    InMux I__741 (
            .O(N__8637),
            .I(N__8627));
    InMux I__740 (
            .O(N__8636),
            .I(N__8623));
    Span4Mux_v I__739 (
            .O(N__8633),
            .I(N__8616));
    LocalMux I__738 (
            .O(N__8630),
            .I(N__8616));
    LocalMux I__737 (
            .O(N__8627),
            .I(N__8616));
    InMux I__736 (
            .O(N__8626),
            .I(N__8613));
    LocalMux I__735 (
            .O(N__8623),
            .I(N__8609));
    Span4Mux_v I__734 (
            .O(N__8616),
            .I(N__8604));
    LocalMux I__733 (
            .O(N__8613),
            .I(N__8604));
    InMux I__732 (
            .O(N__8612),
            .I(N__8601));
    Span4Mux_v I__731 (
            .O(N__8609),
            .I(N__8596));
    Span4Mux_v I__730 (
            .O(N__8604),
            .I(N__8591));
    LocalMux I__729 (
            .O(N__8601),
            .I(N__8591));
    InMux I__728 (
            .O(N__8600),
            .I(N__8588));
    InMux I__727 (
            .O(N__8599),
            .I(N__8585));
    Span4Mux_v I__726 (
            .O(N__8596),
            .I(N__8582));
    Span4Mux_v I__725 (
            .O(N__8591),
            .I(N__8579));
    LocalMux I__724 (
            .O(N__8588),
            .I(N__8576));
    LocalMux I__723 (
            .O(N__8585),
            .I(N__8573));
    Sp12to4 I__722 (
            .O(N__8582),
            .I(N__8570));
    Span4Mux_v I__721 (
            .O(N__8579),
            .I(N__8567));
    Span4Mux_h I__720 (
            .O(N__8576),
            .I(N__8564));
    Span4Mux_h I__719 (
            .O(N__8573),
            .I(N__8561));
    Span12Mux_h I__718 (
            .O(N__8570),
            .I(N__8558));
    Sp12to4 I__717 (
            .O(N__8567),
            .I(N__8555));
    IoSpan4Mux I__716 (
            .O(N__8564),
            .I(N__8552));
    Span4Mux_h I__715 (
            .O(N__8561),
            .I(N__8549));
    Span12Mux_v I__714 (
            .O(N__8558),
            .I(N__8546));
    Span12Mux_h I__713 (
            .O(N__8555),
            .I(N__8543));
    IoSpan4Mux I__712 (
            .O(N__8552),
            .I(N__8540));
    Span4Mux_h I__711 (
            .O(N__8549),
            .I(N__8537));
    Odrv12 I__710 (
            .O(N__8546),
            .I(TVP_VIDEO_c_8));
    Odrv12 I__709 (
            .O(N__8543),
            .I(TVP_VIDEO_c_8));
    Odrv4 I__708 (
            .O(N__8540),
            .I(TVP_VIDEO_c_8));
    Odrv4 I__707 (
            .O(N__8537),
            .I(TVP_VIDEO_c_8));
    InMux I__706 (
            .O(N__8528),
            .I(N__8524));
    InMux I__705 (
            .O(N__8527),
            .I(N__8521));
    LocalMux I__704 (
            .O(N__8524),
            .I(N__8515));
    LocalMux I__703 (
            .O(N__8521),
            .I(N__8515));
    InMux I__702 (
            .O(N__8520),
            .I(N__8512));
    Span4Mux_v I__701 (
            .O(N__8515),
            .I(N__8507));
    LocalMux I__700 (
            .O(N__8512),
            .I(N__8507));
    Span4Mux_v I__699 (
            .O(N__8507),
            .I(N__8503));
    InMux I__698 (
            .O(N__8506),
            .I(N__8500));
    Span4Mux_v I__697 (
            .O(N__8503),
            .I(N__8494));
    LocalMux I__696 (
            .O(N__8500),
            .I(N__8494));
    InMux I__695 (
            .O(N__8499),
            .I(N__8490));
    Span4Mux_h I__694 (
            .O(N__8494),
            .I(N__8487));
    InMux I__693 (
            .O(N__8493),
            .I(N__8484));
    LocalMux I__692 (
            .O(N__8490),
            .I(N__8481));
    Span4Mux_v I__691 (
            .O(N__8487),
            .I(N__8478));
    LocalMux I__690 (
            .O(N__8484),
            .I(N__8475));
    Span12Mux_s11_h I__689 (
            .O(N__8481),
            .I(N__8471));
    Sp12to4 I__688 (
            .O(N__8478),
            .I(N__8468));
    Span12Mux_s8_h I__687 (
            .O(N__8475),
            .I(N__8465));
    InMux I__686 (
            .O(N__8474),
            .I(N__8462));
    Span12Mux_v I__685 (
            .O(N__8471),
            .I(N__8459));
    Span12Mux_v I__684 (
            .O(N__8468),
            .I(N__8456));
    Span12Mux_v I__683 (
            .O(N__8465),
            .I(N__8453));
    LocalMux I__682 (
            .O(N__8462),
            .I(N__8450));
    Span12Mux_h I__681 (
            .O(N__8459),
            .I(N__8446));
    Span12Mux_h I__680 (
            .O(N__8456),
            .I(N__8441));
    Span12Mux_v I__679 (
            .O(N__8453),
            .I(N__8441));
    Span4Mux_h I__678 (
            .O(N__8450),
            .I(N__8438));
    InMux I__677 (
            .O(N__8449),
            .I(N__8435));
    Odrv12 I__676 (
            .O(N__8446),
            .I(TVP_VIDEO_c_9));
    Odrv12 I__675 (
            .O(N__8441),
            .I(TVP_VIDEO_c_9));
    Odrv4 I__674 (
            .O(N__8438),
            .I(TVP_VIDEO_c_9));
    LocalMux I__673 (
            .O(N__8435),
            .I(TVP_VIDEO_c_9));
    InMux I__672 (
            .O(N__8426),
            .I(N__8423));
    LocalMux I__671 (
            .O(N__8423),
            .I(N__8417));
    InMux I__670 (
            .O(N__8422),
            .I(N__8414));
    InMux I__669 (
            .O(N__8421),
            .I(N__8411));
    InMux I__668 (
            .O(N__8420),
            .I(N__8408));
    Span4Mux_h I__667 (
            .O(N__8417),
            .I(N__8405));
    LocalMux I__666 (
            .O(N__8414),
            .I(N__8401));
    LocalMux I__665 (
            .O(N__8411),
            .I(N__8398));
    LocalMux I__664 (
            .O(N__8408),
            .I(N__8394));
    Span4Mux_h I__663 (
            .O(N__8405),
            .I(N__8391));
    InMux I__662 (
            .O(N__8404),
            .I(N__8388));
    Span4Mux_h I__661 (
            .O(N__8401),
            .I(N__8385));
    Span4Mux_v I__660 (
            .O(N__8398),
            .I(N__8382));
    InMux I__659 (
            .O(N__8397),
            .I(N__8377));
    Span12Mux_h I__658 (
            .O(N__8394),
            .I(N__8374));
    Sp12to4 I__657 (
            .O(N__8391),
            .I(N__8371));
    LocalMux I__656 (
            .O(N__8388),
            .I(N__8368));
    Span4Mux_h I__655 (
            .O(N__8385),
            .I(N__8365));
    Span4Mux_v I__654 (
            .O(N__8382),
            .I(N__8362));
    InMux I__653 (
            .O(N__8381),
            .I(N__8359));
    InMux I__652 (
            .O(N__8380),
            .I(N__8356));
    LocalMux I__651 (
            .O(N__8377),
            .I(N__8353));
    Span12Mux_v I__650 (
            .O(N__8374),
            .I(N__8350));
    Span12Mux_v I__649 (
            .O(N__8371),
            .I(N__8343));
    Span12Mux_h I__648 (
            .O(N__8368),
            .I(N__8343));
    Sp12to4 I__647 (
            .O(N__8365),
            .I(N__8343));
    Sp12to4 I__646 (
            .O(N__8362),
            .I(N__8338));
    LocalMux I__645 (
            .O(N__8359),
            .I(N__8338));
    LocalMux I__644 (
            .O(N__8356),
            .I(N__8335));
    Span4Mux_h I__643 (
            .O(N__8353),
            .I(N__8332));
    Span12Mux_v I__642 (
            .O(N__8350),
            .I(N__8329));
    Span12Mux_v I__641 (
            .O(N__8343),
            .I(N__8322));
    Span12Mux_h I__640 (
            .O(N__8338),
            .I(N__8322));
    Span12Mux_h I__639 (
            .O(N__8335),
            .I(N__8322));
    Span4Mux_h I__638 (
            .O(N__8332),
            .I(N__8319));
    Odrv12 I__637 (
            .O(N__8329),
            .I(TVP_VIDEO_c_7));
    Odrv12 I__636 (
            .O(N__8322),
            .I(TVP_VIDEO_c_7));
    Odrv4 I__635 (
            .O(N__8319),
            .I(TVP_VIDEO_c_7));
    InMux I__634 (
            .O(N__8312),
            .I(N__8308));
    InMux I__633 (
            .O(N__8311),
            .I(N__8305));
    LocalMux I__632 (
            .O(N__8308),
            .I(N__8302));
    LocalMux I__631 (
            .O(N__8305),
            .I(N__8298));
    Span4Mux_v I__630 (
            .O(N__8302),
            .I(N__8295));
    InMux I__629 (
            .O(N__8301),
            .I(N__8292));
    Span4Mux_v I__628 (
            .O(N__8298),
            .I(N__8288));
    Span4Mux_v I__627 (
            .O(N__8295),
            .I(N__8283));
    LocalMux I__626 (
            .O(N__8292),
            .I(N__8283));
    InMux I__625 (
            .O(N__8291),
            .I(N__8280));
    Span4Mux_v I__624 (
            .O(N__8288),
            .I(N__8277));
    Span4Mux_v I__623 (
            .O(N__8283),
            .I(N__8271));
    LocalMux I__622 (
            .O(N__8280),
            .I(N__8271));
    Span4Mux_v I__621 (
            .O(N__8277),
            .I(N__8267));
    InMux I__620 (
            .O(N__8276),
            .I(N__8264));
    Span4Mux_v I__619 (
            .O(N__8271),
            .I(N__8260));
    InMux I__618 (
            .O(N__8270),
            .I(N__8257));
    Span4Mux_v I__617 (
            .O(N__8267),
            .I(N__8252));
    LocalMux I__616 (
            .O(N__8264),
            .I(N__8252));
    InMux I__615 (
            .O(N__8263),
            .I(N__8249));
    Span4Mux_v I__614 (
            .O(N__8260),
            .I(N__8244));
    LocalMux I__613 (
            .O(N__8257),
            .I(N__8244));
    Span4Mux_v I__612 (
            .O(N__8252),
            .I(N__8239));
    LocalMux I__611 (
            .O(N__8249),
            .I(N__8239));
    Span4Mux_v I__610 (
            .O(N__8244),
            .I(N__8235));
    Span4Mux_v I__609 (
            .O(N__8239),
            .I(N__8232));
    InMux I__608 (
            .O(N__8238),
            .I(N__8229));
    Sp12to4 I__607 (
            .O(N__8235),
            .I(N__8226));
    Span4Mux_v I__606 (
            .O(N__8232),
            .I(N__8221));
    LocalMux I__605 (
            .O(N__8229),
            .I(N__8221));
    Span12Mux_h I__604 (
            .O(N__8226),
            .I(N__8218));
    Span4Mux_h I__603 (
            .O(N__8221),
            .I(N__8215));
    Odrv12 I__602 (
            .O(N__8218),
            .I(TVP_VIDEO_c_6));
    Odrv4 I__601 (
            .O(N__8215),
            .I(TVP_VIDEO_c_6));
    InMux I__600 (
            .O(N__8210),
            .I(N__8206));
    InMux I__599 (
            .O(N__8209),
            .I(N__8203));
    LocalMux I__598 (
            .O(N__8206),
            .I(N__8200));
    LocalMux I__597 (
            .O(N__8203),
            .I(N__8196));
    Span4Mux_v I__596 (
            .O(N__8200),
            .I(N__8193));
    InMux I__595 (
            .O(N__8199),
            .I(N__8190));
    Span4Mux_v I__594 (
            .O(N__8196),
            .I(N__8187));
    Span4Mux_v I__593 (
            .O(N__8193),
            .I(N__8181));
    LocalMux I__592 (
            .O(N__8190),
            .I(N__8181));
    Span4Mux_v I__591 (
            .O(N__8187),
            .I(N__8177));
    InMux I__590 (
            .O(N__8186),
            .I(N__8174));
    Span4Mux_v I__589 (
            .O(N__8181),
            .I(N__8171));
    InMux I__588 (
            .O(N__8180),
            .I(N__8168));
    Span4Mux_v I__587 (
            .O(N__8177),
            .I(N__8162));
    LocalMux I__586 (
            .O(N__8174),
            .I(N__8162));
    Span4Mux_v I__585 (
            .O(N__8171),
            .I(N__8156));
    LocalMux I__584 (
            .O(N__8168),
            .I(N__8156));
    InMux I__583 (
            .O(N__8167),
            .I(N__8153));
    Span4Mux_v I__582 (
            .O(N__8162),
            .I(N__8150));
    InMux I__581 (
            .O(N__8161),
            .I(N__8147));
    Span4Mux_v I__580 (
            .O(N__8156),
            .I(N__8142));
    LocalMux I__579 (
            .O(N__8153),
            .I(N__8142));
    Span4Mux_v I__578 (
            .O(N__8150),
            .I(N__8137));
    LocalMux I__577 (
            .O(N__8147),
            .I(N__8137));
    Span4Mux_v I__576 (
            .O(N__8142),
            .I(N__8133));
    Span4Mux_v I__575 (
            .O(N__8137),
            .I(N__8130));
    InMux I__574 (
            .O(N__8136),
            .I(N__8127));
    Sp12to4 I__573 (
            .O(N__8133),
            .I(N__8124));
    Span4Mux_v I__572 (
            .O(N__8130),
            .I(N__8119));
    LocalMux I__571 (
            .O(N__8127),
            .I(N__8119));
    Span12Mux_h I__570 (
            .O(N__8124),
            .I(N__8116));
    Span4Mux_h I__569 (
            .O(N__8119),
            .I(N__8113));
    Odrv12 I__568 (
            .O(N__8116),
            .I(TVP_VIDEO_c_5));
    Odrv4 I__567 (
            .O(N__8113),
            .I(TVP_VIDEO_c_5));
    InMux I__566 (
            .O(N__8108),
            .I(N__8105));
    LocalMux I__565 (
            .O(N__8105),
            .I(N__8102));
    Span4Mux_v I__564 (
            .O(N__8102),
            .I(N__8096));
    InMux I__563 (
            .O(N__8101),
            .I(N__8093));
    InMux I__562 (
            .O(N__8100),
            .I(N__8089));
    InMux I__561 (
            .O(N__8099),
            .I(N__8085));
    Span4Mux_v I__560 (
            .O(N__8096),
            .I(N__8080));
    LocalMux I__559 (
            .O(N__8093),
            .I(N__8080));
    InMux I__558 (
            .O(N__8092),
            .I(N__8077));
    LocalMux I__557 (
            .O(N__8089),
            .I(N__8074));
    InMux I__556 (
            .O(N__8088),
            .I(N__8071));
    LocalMux I__555 (
            .O(N__8085),
            .I(N__8068));
    Span4Mux_v I__554 (
            .O(N__8080),
            .I(N__8063));
    LocalMux I__553 (
            .O(N__8077),
            .I(N__8063));
    Span4Mux_h I__552 (
            .O(N__8074),
            .I(N__8060));
    LocalMux I__551 (
            .O(N__8071),
            .I(N__8057));
    Span4Mux_s1_v I__550 (
            .O(N__8068),
            .I(N__8053));
    Span4Mux_v I__549 (
            .O(N__8063),
            .I(N__8050));
    Span4Mux_h I__548 (
            .O(N__8060),
            .I(N__8047));
    Span4Mux_h I__547 (
            .O(N__8057),
            .I(N__8044));
    InMux I__546 (
            .O(N__8056),
            .I(N__8041));
    Sp12to4 I__545 (
            .O(N__8053),
            .I(N__8038));
    Span4Mux_h I__544 (
            .O(N__8050),
            .I(N__8035));
    Span4Mux_h I__543 (
            .O(N__8047),
            .I(N__8032));
    Span4Mux_v I__542 (
            .O(N__8044),
            .I(N__8029));
    LocalMux I__541 (
            .O(N__8041),
            .I(N__8026));
    Span12Mux_s10_h I__540 (
            .O(N__8038),
            .I(N__8022));
    Sp12to4 I__539 (
            .O(N__8035),
            .I(N__8019));
    Span4Mux_h I__538 (
            .O(N__8032),
            .I(N__8012));
    Span4Mux_v I__537 (
            .O(N__8029),
            .I(N__8012));
    Span4Mux_h I__536 (
            .O(N__8026),
            .I(N__8012));
    InMux I__535 (
            .O(N__8025),
            .I(N__8009));
    Span12Mux_v I__534 (
            .O(N__8022),
            .I(N__8006));
    Span12Mux_h I__533 (
            .O(N__8019),
            .I(N__8003));
    Span4Mux_v I__532 (
            .O(N__8012),
            .I(N__8000));
    LocalMux I__531 (
            .O(N__8009),
            .I(N__7997));
    Span12Mux_v I__530 (
            .O(N__8006),
            .I(N__7994));
    Span12Mux_v I__529 (
            .O(N__8003),
            .I(N__7991));
    Span4Mux_v I__528 (
            .O(N__8000),
            .I(N__7988));
    Span4Mux_h I__527 (
            .O(N__7997),
            .I(N__7985));
    Odrv12 I__526 (
            .O(N__7994),
            .I(TVP_VIDEO_c_4));
    Odrv12 I__525 (
            .O(N__7991),
            .I(TVP_VIDEO_c_4));
    Odrv4 I__524 (
            .O(N__7988),
            .I(TVP_VIDEO_c_4));
    Odrv4 I__523 (
            .O(N__7985),
            .I(TVP_VIDEO_c_4));
    InMux I__522 (
            .O(N__7976),
            .I(N__7973));
    LocalMux I__521 (
            .O(N__7973),
            .I(N__7970));
    Span4Mux_v I__520 (
            .O(N__7970),
            .I(N__7966));
    InMux I__519 (
            .O(N__7969),
            .I(N__7963));
    Span4Mux_v I__518 (
            .O(N__7966),
            .I(N__7957));
    LocalMux I__517 (
            .O(N__7963),
            .I(N__7957));
    InMux I__516 (
            .O(N__7962),
            .I(N__7954));
    Span4Mux_v I__515 (
            .O(N__7957),
            .I(N__7951));
    LocalMux I__514 (
            .O(N__7954),
            .I(N__7948));
    Span4Mux_v I__513 (
            .O(N__7951),
            .I(N__7942));
    Span4Mux_v I__512 (
            .O(N__7948),
            .I(N__7942));
    InMux I__511 (
            .O(N__7947),
            .I(N__7939));
    Span4Mux_v I__510 (
            .O(N__7942),
            .I(N__7933));
    LocalMux I__509 (
            .O(N__7939),
            .I(N__7933));
    InMux I__508 (
            .O(N__7938),
            .I(N__7930));
    Span4Mux_v I__507 (
            .O(N__7933),
            .I(N__7924));
    LocalMux I__506 (
            .O(N__7930),
            .I(N__7924));
    InMux I__505 (
            .O(N__7929),
            .I(N__7921));
    Span4Mux_v I__504 (
            .O(N__7924),
            .I(N__7916));
    LocalMux I__503 (
            .O(N__7921),
            .I(N__7913));
    InMux I__502 (
            .O(N__7920),
            .I(N__7910));
    InMux I__501 (
            .O(N__7919),
            .I(N__7907));
    Sp12to4 I__500 (
            .O(N__7916),
            .I(N__7904));
    Span4Mux_h I__499 (
            .O(N__7913),
            .I(N__7901));
    LocalMux I__498 (
            .O(N__7910),
            .I(N__7898));
    LocalMux I__497 (
            .O(N__7907),
            .I(N__7895));
    Span12Mux_h I__496 (
            .O(N__7904),
            .I(N__7892));
    Sp12to4 I__495 (
            .O(N__7901),
            .I(N__7889));
    Span4Mux_h I__494 (
            .O(N__7898),
            .I(N__7886));
    Span12Mux_h I__493 (
            .O(N__7895),
            .I(N__7883));
    Span12Mux_h I__492 (
            .O(N__7892),
            .I(N__7876));
    Span12Mux_v I__491 (
            .O(N__7889),
            .I(N__7876));
    Sp12to4 I__490 (
            .O(N__7886),
            .I(N__7876));
    Odrv12 I__489 (
            .O(N__7883),
            .I(TVP_VIDEO_c_3));
    Odrv12 I__488 (
            .O(N__7876),
            .I(TVP_VIDEO_c_3));
    INV INVADV_R__i1C (
            .O(INVADV_R__i1C_net),
            .I(N__22090));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3373 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3384 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(\transmit_module.n3343 ),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3356 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3364 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\receive_module.n3330 ),
            .carryinitout(bfn_14_12_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_6_17_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_6_17_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_6_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i53_LC_6_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8660),
            .lcout(\transmit_module.Y_DELTA_PATTERN_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22149),
            .ce(N__17981),
            .sr(N__20660));
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_6_17_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_6_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_6_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i55_LC_6_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8921),
            .lcout(\transmit_module.Y_DELTA_PATTERN_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22149),
            .ce(N__17981),
            .sr(N__20660));
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_6_17_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_6_17_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_6_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i54_LC_6_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8666),
            .lcout(\transmit_module.Y_DELTA_PATTERN_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22149),
            .ce(N__17981),
            .sr(N__20660));
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_6_17_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_6_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_6_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i52_LC_6_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8654),
            .lcout(\transmit_module.Y_DELTA_PATTERN_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22149),
            .ce(N__17981),
            .sr(N__20660));
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_6_17_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_6_17_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_6_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i51_LC_6_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8648),
            .lcout(\transmit_module.Y_DELTA_PATTERN_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22149),
            .ce(N__17981),
            .sr(N__20660));
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_7_17_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_7_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i63_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9128),
            .lcout(\transmit_module.Y_DELTA_PATTERN_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22070),
            .ce(N__17980),
            .sr(N__20690));
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_7_19_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_7_19_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i9_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8864),
            .lcout(\transmit_module.X_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22087),
            .ce(N__12880),
            .sr(N__18724));
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_9_13_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_9_13_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_9_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i19_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8975),
            .lcout(\transmit_module.Y_DELTA_PATTERN_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21816),
            .ce(N__18713),
            .sr(N__20568));
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_9_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_9_13_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_9_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i13_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8813),
            .lcout(\transmit_module.Y_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21816),
            .ce(N__18713),
            .sr(N__20568));
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_9_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_9_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i14_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8807),
            .lcout(\transmit_module.Y_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21816),
            .ce(N__18713),
            .sr(N__20568));
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_9_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_9_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_9_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i15_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8801),
            .lcout(\transmit_module.Y_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21816),
            .ce(N__18713),
            .sr(N__20568));
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_9_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_9_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_9_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i16_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8795),
            .lcout(\transmit_module.Y_DELTA_PATTERN_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21816),
            .ce(N__18713),
            .sr(N__20568));
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_9_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_9_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i17_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8783),
            .lcout(\transmit_module.Y_DELTA_PATTERN_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21816),
            .ce(N__18713),
            .sr(N__20568));
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_9_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_9_13_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_9_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i18_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8789),
            .lcout(\transmit_module.Y_DELTA_PATTERN_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21816),
            .ce(N__18713),
            .sr(N__20568));
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_9_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_9_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_9_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i70_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8849),
            .lcout(\transmit_module.Y_DELTA_PATTERN_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22139),
            .ce(N__17939),
            .sr(N__20717));
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_9_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_9_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i71_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9383),
            .lcout(\transmit_module.Y_DELTA_PATTERN_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22139),
            .ce(N__17939),
            .sr(N__20717));
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9062),
            .lcout(\transmit_module.Y_DELTA_PATTERN_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22139),
            .ce(N__17939),
            .sr(N__20717));
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_9_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_9_15_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_9_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i69_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8843),
            .lcout(\transmit_module.Y_DELTA_PATTERN_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22139),
            .ce(N__17939),
            .sr(N__20717));
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_9_16_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_9_16_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_9_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i59_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8837),
            .lcout(\transmit_module.Y_DELTA_PATTERN_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22086),
            .ce(N__17984),
            .sr(N__20713));
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_9_16_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_9_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i60_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8897),
            .lcout(\transmit_module.Y_DELTA_PATTERN_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22086),
            .ce(N__17984),
            .sr(N__20713));
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_9_16_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_9_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i58_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8831),
            .lcout(\transmit_module.Y_DELTA_PATTERN_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22086),
            .ce(N__17984),
            .sr(N__20713));
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_9_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_9_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_9_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i40_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8819),
            .lcout(\transmit_module.Y_DELTA_PATTERN_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22086),
            .ce(N__17984),
            .sr(N__20713));
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_9_16_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_9_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i41_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8825),
            .lcout(\transmit_module.Y_DELTA_PATTERN_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22086),
            .ce(N__17984),
            .sr(N__20713));
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_16_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i68_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8927),
            .lcout(\transmit_module.Y_DELTA_PATTERN_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22086),
            .ce(N__17984),
            .sr(N__20713));
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_9_17_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_9_17_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_9_17_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i56_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__8903),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22088),
            .ce(N__17983),
            .sr(N__20691));
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_9_17_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_9_17_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_9_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i57_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8909),
            .lcout(\transmit_module.Y_DELTA_PATTERN_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22088),
            .ce(N__17983),
            .sr(N__20691));
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_9_17_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_9_17_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_9_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i61_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9158),
            .lcout(\transmit_module.Y_DELTA_PATTERN_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22088),
            .ce(N__17983),
            .sr(N__20691));
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_9_17_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_9_17_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_9_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i48_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9140),
            .lcout(\transmit_module.Y_DELTA_PATTERN_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22088),
            .ce(N__17983),
            .sr(N__20691));
    defparam \line_buffer.i2341_3_lut_LC_9_18_0 .C_ON=1'b0;
    defparam \line_buffer.i2341_3_lut_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2341_3_lut_LC_9_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2341_3_lut_LC_9_18_0  (
            .in0(N__8891),
            .in1(N__8879),
            .in2(_gnd_net_),
            .in3(N__23108),
            .lcout(\line_buffer.n3703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_9_19_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_9_19_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_9_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i11_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9119),
            .lcout(\transmit_module.X_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(N__12878),
            .sr(N__18703));
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_9_19_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_9_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i10_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8870),
            .lcout(\transmit_module.X_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(N__12878),
            .sr(N__18703));
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_10_10_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_10_10_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_10_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i23_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8855),
            .lcout(\transmit_module.Y_DELTA_PATTERN_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22145),
            .ce(N__18730),
            .sr(N__20698));
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_10_10_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_10_10_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_10_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i24_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9269),
            .lcout(\transmit_module.Y_DELTA_PATTERN_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22145),
            .ce(N__18730),
            .sr(N__20698));
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_10_11_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i6_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9263),
            .lcout(\transmit_module.Y_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22143),
            .ce(N__18731),
            .sr(N__20694));
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_10_11_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_10_11_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_10_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i5_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8981),
            .lcout(\transmit_module.Y_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22143),
            .ce(N__18731),
            .sr(N__20694));
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_10_12_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_10_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i20_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8969),
            .lcout(\transmit_module.Y_DELTA_PATTERN_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22104),
            .ce(N__18726),
            .sr(N__20697));
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_10_12_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_10_12_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i21_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8954),
            .lcout(\transmit_module.Y_DELTA_PATTERN_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22104),
            .ce(N__18726),
            .sr(N__20697));
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_10_12_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_10_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i22_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8963),
            .lcout(\transmit_module.Y_DELTA_PATTERN_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22104),
            .ce(N__18726),
            .sr(N__20697));
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_10_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_10_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i4_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8948),
            .lcout(\transmit_module.Y_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22142),
            .ce(N__18725),
            .sr(N__20695));
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_10_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_10_13_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_10_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i0_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8939),
            .lcout(\transmit_module.Y_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22142),
            .ce(N__18725),
            .sr(N__20695));
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_10_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_10_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i1_LC_10_13_5  (
            .in0(N__9005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22142),
            .ce(N__18725),
            .sr(N__20695));
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_10_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_10_13_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_10_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i3_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8933),
            .lcout(\transmit_module.Y_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22142),
            .ce(N__18725),
            .sr(N__20695));
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_10_14_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_10_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i44_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9023),
            .lcout(\transmit_module.Y_DELTA_PATTERN_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22103),
            .ce(N__17962),
            .sr(N__20517));
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9017),
            .lcout(\transmit_module.Y_DELTA_PATTERN_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22103),
            .ce(N__17962),
            .sr(N__20517));
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_10_14_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_10_14_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_10_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i45_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8999),
            .lcout(\transmit_module.Y_DELTA_PATTERN_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22103),
            .ce(N__17962),
            .sr(N__20517));
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8993),
            .lcout(\transmit_module.Y_DELTA_PATTERN_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22103),
            .ce(N__17962),
            .sr(N__20517));
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_10_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_10_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_10_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i2_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9011),
            .lcout(\transmit_module.Y_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22103),
            .ce(N__17962),
            .sr(N__20517));
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i46_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9086),
            .lcout(\transmit_module.Y_DELTA_PATTERN_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22103),
            .ce(N__17962),
            .sr(N__20517));
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_10_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_10_14_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_10_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i78_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9101),
            .lcout(\transmit_module.Y_DELTA_PATTERN_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22103),
            .ce(N__17962),
            .sr(N__20517));
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_10_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_10_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_10_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i67_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8987),
            .lcout(\transmit_module.Y_DELTA_PATTERN_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22138),
            .ce(N__17970),
            .sr(N__20649));
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_10_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_10_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_10_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i81_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9074),
            .lcout(\transmit_module.Y_DELTA_PATTERN_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22138),
            .ce(N__17970),
            .sr(N__20649));
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_10_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_10_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i79_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9050),
            .lcout(\transmit_module.Y_DELTA_PATTERN_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22138),
            .ce(N__17970),
            .sr(N__20649));
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9095),
            .lcout(\transmit_module.Y_DELTA_PATTERN_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22138),
            .ce(N__17970),
            .sr(N__20649));
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_10_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_10_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i66_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9080),
            .lcout(\transmit_module.Y_DELTA_PATTERN_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22138),
            .ce(N__17970),
            .sr(N__20649));
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i82_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9323),
            .lcout(\transmit_module.Y_DELTA_PATTERN_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22138),
            .ce(N__17970),
            .sr(N__20649));
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__9068),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22138),
            .ce(N__17970),
            .sr(N__20649));
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_10_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_10_15_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_10_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i80_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9056),
            .lcout(\transmit_module.Y_DELTA_PATTERN_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22138),
            .ce(N__17970),
            .sr(N__20649));
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_16_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i74_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9029),
            .lcout(\transmit_module.Y_DELTA_PATTERN_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22099),
            .ce(N__17969),
            .sr(N__20518));
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_16_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_16_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i65_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9044),
            .lcout(\transmit_module.Y_DELTA_PATTERN_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22099),
            .ce(N__17969),
            .sr(N__20518));
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i75_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9038),
            .lcout(\transmit_module.Y_DELTA_PATTERN_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22099),
            .ce(N__17969),
            .sr(N__20518));
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_17_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_17_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i50_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9176),
            .lcout(\transmit_module.Y_DELTA_PATTERN_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22118),
            .ce(N__17982),
            .sr(N__20656));
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_17_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_17_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i62_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9167),
            .lcout(\transmit_module.Y_DELTA_PATTERN_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22118),
            .ce(N__17982),
            .sr(N__20656));
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_17_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_17_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i73_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9152),
            .lcout(\transmit_module.Y_DELTA_PATTERN_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22118),
            .ce(N__17982),
            .sr(N__20656));
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_17_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i49_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9146),
            .lcout(\transmit_module.Y_DELTA_PATTERN_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22118),
            .ce(N__17982),
            .sr(N__20656));
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_17_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_17_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i64_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9134),
            .lcout(\transmit_module.Y_DELTA_PATTERN_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22118),
            .ce(N__17982),
            .sr(N__20656));
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_10_19_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_10_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i12_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9113),
            .lcout(\transmit_module.X_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21983),
            .ce(N__12881),
            .sr(N__18701));
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_10_19_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_10_19_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_10_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i13_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9593),
            .lcout(\transmit_module.X_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21983),
            .ce(N__12881),
            .sr(N__18701));
    defparam \receive_module.rx_counter.old_HS_50_LC_11_8_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_HS_50_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_HS_50_LC_11_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receive_module.rx_counter.old_HS_50_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19913),
            .lcout(old_HS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21009),
            .ce(),
            .sr(_gnd_net_));
    defparam i272_3_lut_3_lut_LC_11_8_6.C_ON=1'b0;
    defparam i272_3_lut_3_lut_LC_11_8_6.SEQ_MODE=4'b0000;
    defparam i272_3_lut_3_lut_LC_11_8_6.LUT_INIT=16'b0100010011111111;
    LogicCell40 i272_3_lut_3_lut_LC_11_8_6 (
            .in0(N__19912),
            .in1(N__9107),
            .in2(_gnd_net_),
            .in3(N__17770),
            .lcout(n2057),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.Y__i0_LC_11_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i0_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i0_LC_11_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i0_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__9968),
            .in2(_gnd_net_),
            .in3(N__9221),
            .lcout(\receive_module.rx_counter.Y_0 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\receive_module.rx_counter.n3349 ),
            .clk(N__21012),
            .ce(N__9190),
            .sr(N__17697));
    defparam \receive_module.rx_counter.Y__i1_LC_11_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i1_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i1_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i1_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__11074),
            .in2(_gnd_net_),
            .in3(N__9218),
            .lcout(\receive_module.rx_counter.Y_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3349 ),
            .carryout(\receive_module.rx_counter.n3350 ),
            .clk(N__21012),
            .ce(N__9190),
            .sr(N__17697));
    defparam \receive_module.rx_counter.Y__i2_LC_11_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i2_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i2_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i2_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__9940),
            .in2(_gnd_net_),
            .in3(N__9215),
            .lcout(\receive_module.rx_counter.Y_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3350 ),
            .carryout(\receive_module.rx_counter.n3351 ),
            .clk(N__21012),
            .ce(N__9190),
            .sr(N__17697));
    defparam \receive_module.rx_counter.Y__i3_LC_11_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i3_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i3_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i3_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__11104),
            .in2(_gnd_net_),
            .in3(N__9212),
            .lcout(\receive_module.rx_counter.Y_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3351 ),
            .carryout(\receive_module.rx_counter.n3352 ),
            .clk(N__21012),
            .ce(N__9190),
            .sr(N__17697));
    defparam \receive_module.rx_counter.Y__i4_LC_11_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i4_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i4_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i4_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__11134),
            .in2(_gnd_net_),
            .in3(N__9209),
            .lcout(\receive_module.rx_counter.Y_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3352 ),
            .carryout(\receive_module.rx_counter.n3353 ),
            .clk(N__21012),
            .ce(N__9190),
            .sr(N__17697));
    defparam \receive_module.rx_counter.Y__i5_LC_11_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i5_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i5_LC_11_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i5_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__9539),
            .in2(_gnd_net_),
            .in3(N__9206),
            .lcout(\receive_module.rx_counter.Y_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3353 ),
            .carryout(\receive_module.rx_counter.n3354 ),
            .clk(N__21012),
            .ce(N__9190),
            .sr(N__17697));
    defparam \receive_module.rx_counter.Y__i6_LC_11_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i6_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i6_LC_11_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i6_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__9554),
            .in2(_gnd_net_),
            .in3(N__9203),
            .lcout(\receive_module.rx_counter.Y_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3354 ),
            .carryout(\receive_module.rx_counter.n3355 ),
            .clk(N__21012),
            .ce(N__9190),
            .sr(N__17697));
    defparam \receive_module.rx_counter.Y__i7_LC_11_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i7_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i7_LC_11_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i7_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__9992),
            .in2(_gnd_net_),
            .in3(N__9200),
            .lcout(\receive_module.rx_counter.Y_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3355 ),
            .carryout(\receive_module.rx_counter.n3356 ),
            .clk(N__21012),
            .ce(N__9190),
            .sr(N__17697));
    defparam \receive_module.rx_counter.Y__i8_LC_11_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.Y__i8_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i8_LC_11_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i8_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__10009),
            .in2(_gnd_net_),
            .in3(N__9197),
            .lcout(\receive_module.rx_counter.Y_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21017),
            .ce(N__9194),
            .sr(N__17675));
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_11_11_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_11_11_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_11_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i26_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9257),
            .lcout(\transmit_module.Y_DELTA_PATTERN_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22117),
            .ce(N__18712),
            .sr(N__20692));
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_11_11_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_11_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i25_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9275),
            .lcout(\transmit_module.Y_DELTA_PATTERN_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22117),
            .ce(N__18712),
            .sr(N__20692));
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_11_11_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_11_11_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i7_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9227),
            .lcout(\transmit_module.Y_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22117),
            .ce(N__18712),
            .sr(N__20692));
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_11_12_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_11_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i10_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9329),
            .lcout(\transmit_module.Y_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22072),
            .ce(N__18720),
            .sr(N__20696));
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_11_12_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_11_12_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i27_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9416),
            .lcout(\transmit_module.Y_DELTA_PATTERN_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22072),
            .ce(N__18720),
            .sr(N__20696));
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_11_12_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_11_12_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i99_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19188),
            .lcout(\transmit_module.Y_DELTA_PATTERN_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22072),
            .ce(N__18720),
            .sr(N__20696));
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_12_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i9_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9251),
            .lcout(\transmit_module.Y_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22072),
            .ce(N__18720),
            .sr(N__20696));
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_11_12_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i12_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9245),
            .lcout(\transmit_module.Y_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22072),
            .ce(N__18720),
            .sr(N__20696));
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_11_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_11_12_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i8_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9233),
            .lcout(\transmit_module.Y_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22072),
            .ce(N__18720),
            .sr(N__20696));
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_11_12_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_11_12_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i11_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9335),
            .lcout(\transmit_module.Y_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22072),
            .ce(N__18720),
            .sr(N__20696));
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10130),
            .lcout(\transmit_module.Y_DELTA_PATTERN_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22141),
            .ce(N__10079),
            .sr(N__20693));
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_11_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_11_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_11_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i83_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9311),
            .lcout(\transmit_module.Y_DELTA_PATTERN_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22141),
            .ce(N__10079),
            .sr(N__20693));
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_11_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_11_13_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_11_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i84_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9287),
            .lcout(\transmit_module.Y_DELTA_PATTERN_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22141),
            .ce(N__10079),
            .sr(N__20693));
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_11_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i93_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9299),
            .lcout(\transmit_module.Y_DELTA_PATTERN_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22141),
            .ce(N__10079),
            .sr(N__20693));
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9305),
            .lcout(\transmit_module.Y_DELTA_PATTERN_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22141),
            .ce(N__10079),
            .sr(N__20693));
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_11_14_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_11_14_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_11_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i92_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9293),
            .lcout(\transmit_module.Y_DELTA_PATTERN_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22071),
            .ce(N__10067),
            .sr(N__20516));
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_11_14_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_11_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i90_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9365),
            .lcout(\transmit_module.Y_DELTA_PATTERN_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22071),
            .ce(N__10067),
            .sr(N__20516));
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_11_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_11_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i85_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9281),
            .lcout(\transmit_module.Y_DELTA_PATTERN_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22071),
            .ce(N__10067),
            .sr(N__20516));
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_11_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_11_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_11_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i86_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10031),
            .lcout(\transmit_module.Y_DELTA_PATTERN_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22071),
            .ce(N__10067),
            .sr(N__20516));
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_11_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_11_14_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i91_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9371),
            .lcout(\transmit_module.Y_DELTA_PATTERN_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22071),
            .ce(N__10067),
            .sr(N__20516));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i1_LC_11_15_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i1_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i1_LC_11_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i1_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__10100),
            .in2(_gnd_net_),
            .in3(N__9359),
            .lcout(\transmit_module.video_signal_controller.VGA_X_0 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\transmit_module.video_signal_controller.n3377 ),
            .clk(N__22095),
            .ce(),
            .sr(N__17644));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i2_LC_11_15_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i2_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i2_LC_11_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i2_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__10124),
            .in2(_gnd_net_),
            .in3(N__9356),
            .lcout(\transmit_module.video_signal_controller.VGA_X_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3377 ),
            .carryout(\transmit_module.video_signal_controller.n3378 ),
            .clk(N__22095),
            .ce(),
            .sr(N__17644));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i3_LC_11_15_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i3_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i3_LC_11_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i3_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__10112),
            .in2(_gnd_net_),
            .in3(N__9353),
            .lcout(\transmit_module.video_signal_controller.VGA_X_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3378 ),
            .carryout(\transmit_module.video_signal_controller.n3379 ),
            .clk(N__22095),
            .ce(),
            .sr(N__17644));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i4_LC_11_15_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i4_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i4_LC_11_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i4_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__11199),
            .in2(_gnd_net_),
            .in3(N__9350),
            .lcout(\transmit_module.video_signal_controller.VGA_X_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3379 ),
            .carryout(\transmit_module.video_signal_controller.n3380 ),
            .clk(N__22095),
            .ce(),
            .sr(N__17644));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i5_LC_11_15_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i5_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i5_LC_11_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i5_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__11230),
            .in2(_gnd_net_),
            .in3(N__9347),
            .lcout(\transmit_module.video_signal_controller.VGA_X_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3380 ),
            .carryout(\transmit_module.video_signal_controller.n3381 ),
            .clk(N__22095),
            .ce(),
            .sr(N__17644));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i6_LC_11_15_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i6_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i6_LC_11_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i6_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__11173),
            .in2(_gnd_net_),
            .in3(N__9344),
            .lcout(\transmit_module.video_signal_controller.VGA_X_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3381 ),
            .carryout(\transmit_module.video_signal_controller.n3382 ),
            .clk(N__22095),
            .ce(),
            .sr(N__17644));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i7_LC_11_15_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i7_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i7_LC_11_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i7_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__10162),
            .in2(_gnd_net_),
            .in3(N__9341),
            .lcout(\transmit_module.video_signal_controller.VGA_X_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3382 ),
            .carryout(\transmit_module.video_signal_controller.n3383 ),
            .clk(N__22095),
            .ce(),
            .sr(N__17644));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i8_LC_11_15_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i8_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i8_LC_11_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i8_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__10183),
            .in2(_gnd_net_),
            .in3(N__9338),
            .lcout(\transmit_module.video_signal_controller.VGA_X_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3383 ),
            .carryout(\transmit_module.video_signal_controller.n3384 ),
            .clk(N__22095),
            .ce(),
            .sr(N__17644));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i9_LC_11_16_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i9_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i9_LC_11_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i9_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__12016),
            .in2(_gnd_net_),
            .in3(N__9425),
            .lcout(\transmit_module.video_signal_controller.VGA_X_8 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\transmit_module.video_signal_controller.n3385 ),
            .clk(N__21949),
            .ce(),
            .sr(N__17645));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i10_LC_11_16_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i10_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i10_LC_11_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i10_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__10698),
            .in2(_gnd_net_),
            .in3(N__9422),
            .lcout(\transmit_module.video_signal_controller.VGA_X_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3385 ),
            .carryout(\transmit_module.video_signal_controller.n3386 ),
            .clk(N__21949),
            .ce(),
            .sr(N__17645));
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i11_LC_11_16_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i11_LC_11_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_266_267__i11_LC_11_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_266_267__i11_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__10732),
            .in2(_gnd_net_),
            .in3(N__9419),
            .lcout(\transmit_module.video_signal_controller.VGA_X_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21949),
            .ce(),
            .sr(N__17645));
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_11_17_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i28_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9407),
            .lcout(\transmit_module.Y_DELTA_PATTERN_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__18707),
            .sr(N__20630));
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_11_17_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_11_17_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_11_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i29_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9401),
            .lcout(\transmit_module.Y_DELTA_PATTERN_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__18707),
            .sr(N__20630));
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_11_17_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_11_17_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_11_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i30_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9395),
            .lcout(\transmit_module.Y_DELTA_PATTERN_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__18707),
            .sr(N__20630));
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_11_17_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i31_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18743),
            .lcout(\transmit_module.Y_DELTA_PATTERN_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__18707),
            .sr(N__20630));
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_17_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_17_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i72_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9389),
            .lcout(\transmit_module.Y_DELTA_PATTERN_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__18707),
            .sr(N__20630));
    defparam \transmit_module.i2_4_lut_LC_11_18_4 .C_ON=1'b0;
    defparam \transmit_module.i2_4_lut_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_4_lut_LC_11_18_4 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \transmit_module.i2_4_lut_LC_11_18_4  (
            .in0(N__16575),
            .in1(N__19708),
            .in2(N__20684),
            .in3(N__19605),
            .lcout(\transmit_module.n2099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1681_4_lut_LC_11_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1681_4_lut_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1681_4_lut_LC_11_19_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1681_4_lut_LC_11_19_0  (
            .in0(N__10660),
            .in1(N__10667),
            .in2(N__20712),
            .in3(N__20252),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_11_20_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_11_20_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_11_20_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i15_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__12931),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22042),
            .ce(N__12867),
            .sr(N__18694));
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_11_20_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_11_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i14_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9599),
            .lcout(\transmit_module.X_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22042),
            .ce(N__12867),
            .sr(N__18694));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2435_LC_11_21_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2435_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2435_LC_11_21_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2435_LC_11_21_2  (
            .in0(N__9587),
            .in1(N__22929),
            .in2(N__9572),
            .in3(N__23132),
            .lcout(\line_buffer.n3785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_rep_25_LC_12_9_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_rep_25_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_rep_25_LC_12_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_rep_25_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__9537),
            .in2(_gnd_net_),
            .in3(N__9552),
            .lcout(\receive_module.rx_counter.n3861 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_4_lut_LC_12_9_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_4_lut_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_4_lut_LC_12_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_4_lut_LC_12_9_1  (
            .in0(N__9553),
            .in1(N__9991),
            .in2(N__10010),
            .in3(N__9538),
            .lcout(\receive_module.rx_counter.n3619 ),
            .ltout(\receive_module.rx_counter.n3619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i4_4_lut_LC_12_9_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i4_4_lut_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i4_4_lut_LC_12_9_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \receive_module.rx_counter.i4_4_lut_LC_12_9_2  (
            .in0(N__11070),
            .in1(N__11100),
            .in2(N__9521),
            .in3(N__11130),
            .lcout(\receive_module.rx_counter.n10_adj_570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_9_3 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_9_3  (
            .in0(N__15912),
            .in1(N__15752),
            .in2(N__15860),
            .in3(N__11302),
            .lcout(\line_buffer.n642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_9_LC_12_9_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_9_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_9_LC_12_9_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_9_LC_12_9_4  (
            .in0(N__11303),
            .in1(N__15913),
            .in2(N__15765),
            .in3(N__15859),
            .lcout(\line_buffer.n578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_LC_12_9_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_LC_12_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__9965),
            .in2(_gnd_net_),
            .in3(N__11069),
            .lcout(),
            .ltout(\receive_module.rx_counter.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_4_lut_LC_12_9_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_4_lut_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_4_lut_LC_12_9_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \receive_module.rx_counter.i1_4_lut_LC_12_9_6  (
            .in0(N__11093),
            .in1(N__11129),
            .in2(N__10013),
            .in3(N__9939),
            .lcout(),
            .ltout(\receive_module.rx_counter.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_LC_12_9_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_LC_12_9_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_LC_12_9_7  (
            .in0(N__10005),
            .in1(N__9990),
            .in2(N__9977),
            .in3(N__9974),
            .lcout(\receive_module.rx_counter.n3657 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_16_LC_12_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_16_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_16_LC_12_10_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_16_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__9938),
            .in2(_gnd_net_),
            .in3(N__9966),
            .lcout(\receive_module.rx_counter.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.SYNC_45_LC_12_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.SYNC_45_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.SYNC_45_LC_12_10_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \receive_module.rx_counter.SYNC_45_LC_12_10_2  (
            .in0(N__9967),
            .in1(N__9947),
            .in2(_gnd_net_),
            .in3(N__9941),
            .lcout(DEBUG_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21013),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_12_10_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_12_10_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_12_10_4  (
            .in0(N__15853),
            .in1(N__15911),
            .in2(N__15760),
            .in3(N__11304),
            .lcout(\line_buffer.n610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2390_2_lut_3_lut_4_lut_LC_12_11_0 .C_ON=1'b0;
    defparam \line_buffer.i2390_2_lut_3_lut_4_lut_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2390_2_lut_3_lut_4_lut_LC_12_11_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \line_buffer.i2390_2_lut_3_lut_4_lut_LC_12_11_0  (
            .in0(N__15847),
            .in1(N__15910),
            .in2(N__15759),
            .in3(N__11308),
            .lcout(\line_buffer.n512 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i13_LC_12_11_1 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i13_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i13_LC_12_11_1 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \receive_module.BRAM_ADDR__i13_LC_12_11_1  (
            .in0(N__11310),
            .in1(N__15739),
            .in2(N__17838),
            .in3(N__15689),
            .lcout(DEBUG_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21018),
            .ce(),
            .sr(N__17690));
    defparam \receive_module.BRAM_ADDR__i3_LC_12_11_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i3_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i3_LC_12_11_2 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \receive_module.BRAM_ADDR__i3_LC_12_11_2  (
            .in0(N__15089),
            .in1(N__15113),
            .in2(N__17836),
            .in3(N__11314),
            .lcout(RX_ADDR_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21018),
            .ce(),
            .sr(N__17690));
    defparam \receive_module.BRAM_ADDR__i2_LC_12_11_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i2_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i2_LC_12_11_3 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \receive_module.BRAM_ADDR__i2_LC_12_11_3  (
            .in0(N__11311),
            .in1(N__15353),
            .in2(N__17840),
            .in3(N__15377),
            .lcout(RX_ADDR_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21018),
            .ce(),
            .sr(N__17690));
    defparam \receive_module.BRAM_ADDR__i1_LC_12_11_4 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i1_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i1_LC_12_11_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \receive_module.BRAM_ADDR__i1_LC_12_11_4  (
            .in0(N__17813),
            .in1(N__12980),
            .in2(N__13035),
            .in3(N__11313),
            .lcout(RX_ADDR_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21018),
            .ce(),
            .sr(N__17690));
    defparam \receive_module.BRAM_ADDR__i10_LC_12_11_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i10_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i10_LC_12_11_5 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \receive_module.BRAM_ADDR__i10_LC_12_11_5  (
            .in0(N__11309),
            .in1(N__15956),
            .in2(N__17837),
            .in3(N__15932),
            .lcout(RX_ADDR_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21018),
            .ce(),
            .sr(N__17690));
    defparam \receive_module.BRAM_ADDR__i9_LC_12_11_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i9_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i9_LC_12_11_6 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \receive_module.BRAM_ADDR__i9_LC_12_11_6  (
            .in0(N__13619),
            .in1(N__13598),
            .in2(N__17835),
            .in3(N__11315),
            .lcout(RX_ADDR_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21018),
            .ce(),
            .sr(N__17690));
    defparam \receive_module.BRAM_ADDR__i8_LC_12_11_7 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i8_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i8_LC_12_11_7 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \receive_module.BRAM_ADDR__i8_LC_12_11_7  (
            .in0(N__11312),
            .in1(N__13880),
            .in2(N__17839),
            .in3(N__13853),
            .lcout(RX_ADDR_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21018),
            .ce(),
            .sr(N__17690));
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_12_12_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_12_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i98_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10043),
            .lcout(\transmit_module.Y_DELTA_PATTERN_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22085),
            .ce(N__10075),
            .sr(N__20367));
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10037),
            .lcout(\transmit_module.Y_DELTA_PATTERN_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22140),
            .ce(N__10074),
            .sr(N__20368));
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10019),
            .lcout(\transmit_module.Y_DELTA_PATTERN_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22140),
            .ce(N__10074),
            .sr(N__20368));
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10025),
            .lcout(\transmit_module.Y_DELTA_PATTERN_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22140),
            .ce(N__10074),
            .sr(N__20368));
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_12_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_12_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i97_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10142),
            .lcout(\transmit_module.Y_DELTA_PATTERN_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22140),
            .ce(N__10074),
            .sr(N__20368));
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_12_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_12_13_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_12_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i96_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10136),
            .lcout(\transmit_module.Y_DELTA_PATTERN_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22140),
            .ce(N__10074),
            .sr(N__20368));
    defparam \transmit_module.video_signal_controller.i3_3_lut_LC_12_14_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i3_3_lut_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i3_3_lut_LC_12_14_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \transmit_module.video_signal_controller.i3_3_lut_LC_12_14_1  (
            .in0(N__10123),
            .in1(_gnd_net_),
            .in2(N__11200),
            .in3(N__10111),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n8_adj_569_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1759_4_lut_LC_12_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1759_4_lut_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1759_4_lut_LC_12_14_2 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \transmit_module.video_signal_controller.i1759_4_lut_LC_12_14_2  (
            .in0(N__11225),
            .in1(N__10099),
            .in2(N__10088),
            .in3(N__12045),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3029_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1777_4_lut_LC_12_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1777_4_lut_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1777_4_lut_LC_12_14_3 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \transmit_module.video_signal_controller.i1777_4_lut_LC_12_14_3  (
            .in0(N__10739),
            .in1(N__10700),
            .in2(N__10085),
            .in3(N__12019),
            .lcout(\transmit_module.video_signal_controller.n2030 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_21_LC_12_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_21_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_21_LC_12_14_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_rep_21_LC_12_14_6  (
            .in0(N__10182),
            .in1(N__11168),
            .in2(_gnd_net_),
            .in3(N__10161),
            .lcout(\transmit_module.video_signal_controller.n3857 ),
            .ltout(\transmit_module.video_signal_controller.n3857_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2242_3_lut_4_lut_LC_12_14_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2242_3_lut_4_lut_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2242_3_lut_4_lut_LC_12_14_7 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \transmit_module.video_signal_controller.i2242_3_lut_4_lut_LC_12_14_7  (
            .in0(N__10738),
            .in1(N__10699),
            .in2(N__10082),
            .in3(N__12018),
            .lcout(\transmit_module.video_signal_controller.n3603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_12_15_0 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_12_15_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i0_LC_12_15_0  (
            .in0(N__16568),
            .in1(N__12755),
            .in2(N__16511),
            .in3(N__19545),
            .lcout(TX_ADDR_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__17497),
            .sr(N__20609));
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_LC_12_15_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_LC_12_15_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_LC_12_15_3  (
            .in0(N__19544),
            .in1(N__16261),
            .in2(N__20572),
            .in3(N__16213),
            .lcout(\transmit_module.n2125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_28_LC_12_15_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_28_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_28_LC_12_15_4 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_28_LC_12_15_4  (
            .in0(N__16260),
            .in1(N__20452),
            .in2(N__16221),
            .in3(N__19543),
            .lcout(\transmit_module.n3864 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1133_1_lut_2_lut_3_lut_4_lut_LC_12_15_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1133_1_lut_2_lut_3_lut_4_lut_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1133_1_lut_2_lut_3_lut_4_lut_LC_12_15_6 .LUT_INIT=16'b0000011111111111;
    LogicCell40 \transmit_module.video_signal_controller.i1133_1_lut_2_lut_3_lut_4_lut_LC_12_15_6  (
            .in0(N__12044),
            .in1(N__12011),
            .in2(N__11974),
            .in3(N__19542),
            .lcout(n2404),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_16_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_16_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__16259),
            .in2(_gnd_net_),
            .in3(N__16208),
            .lcout(\transmit_module.n3859 ),
            .ltout(\transmit_module.n3859_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1076_3_lut_4_lut_LC_12_16_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1076_3_lut_4_lut_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1076_3_lut_4_lut_LC_12_16_1 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \transmit_module.video_signal_controller.i1076_3_lut_4_lut_LC_12_16_1  (
            .in0(N__16481),
            .in1(N__12965),
            .in2(N__10187),
            .in3(N__19589),
            .lcout(\transmit_module.BRAM_ADDR_13_N_256_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_20_LC_12_16_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_20_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_20_LC_12_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_20_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__10730),
            .in2(_gnd_net_),
            .in3(N__10696),
            .lcout(\transmit_module.video_signal_controller.n3856 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.old_VGA_HS_39_LC_12_16_4 .C_ON=1'b0;
    defparam \transmit_module.old_VGA_HS_39_LC_12_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.old_VGA_HS_39_LC_12_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.old_VGA_HS_39_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16209),
            .lcout(\transmit_module.old_VGA_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21948),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_14_LC_12_16_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_14_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_14_LC_12_16_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_adj_14_LC_12_16_5  (
            .in0(N__11226),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11172),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i37_4_lut_LC_12_16_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i37_4_lut_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i37_4_lut_LC_12_16_6 .LUT_INIT=16'b0011001100101110;
    LogicCell40 \transmit_module.video_signal_controller.i37_4_lut_LC_12_16_6  (
            .in0(N__11147),
            .in1(N__10184),
            .in2(N__10166),
            .in3(N__10163),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_HS_54_LC_12_16_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_HS_54_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_HS_54_LC_12_16_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \transmit_module.video_signal_controller.VGA_HS_54_LC_12_16_7  (
            .in0(N__10731),
            .in1(N__12017),
            .in2(N__10145),
            .in3(N__10697),
            .lcout(ADV_HSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21948),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i6_3_lut_LC_12_17_0 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i6_3_lut_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i6_3_lut_LC_12_17_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i6_3_lut_LC_12_17_0  (
            .in0(N__19249),
            .in1(N__16406),
            .in2(_gnd_net_),
            .in3(N__16435),
            .lcout(\transmit_module.n183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_3_lut_4_lut_LC_12_17_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_3_lut_4_lut_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_3_lut_4_lut_LC_12_17_3 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_19_3_lut_4_lut_LC_12_17_3  (
            .in0(N__10729),
            .in1(N__10695),
            .in2(N__12053),
            .in3(N__12012),
            .lcout(\transmit_module.n3855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i7_3_lut_LC_12_18_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i7_3_lut_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i7_3_lut_LC_12_18_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i7_3_lut_LC_12_18_2  (
            .in0(N__19253),
            .in1(N__16682),
            .in2(_gnd_net_),
            .in3(N__16701),
            .lcout(\transmit_module.n182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i7_3_lut_4_lut_LC_12_18_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i7_3_lut_4_lut_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i7_3_lut_4_lut_LC_12_18_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i7_3_lut_4_lut_LC_12_18_3  (
            .in0(N__16702),
            .in1(N__12785),
            .in2(N__19727),
            .in3(N__19607),
            .lcout(\transmit_module.n214 ),
            .ltout(\transmit_module.n214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i6_LC_12_18_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i6_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i6_LC_12_18_4 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i6_LC_12_18_4  (
            .in0(N__20573),
            .in1(N__10661),
            .in2(N__10649),
            .in3(N__20206),
            .lcout(\transmit_module.TX_ADDR_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21947),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1683_4_lut_LC_12_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1683_4_lut_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1683_4_lut_LC_12_19_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1683_4_lut_LC_12_19_0  (
            .in0(N__10918),
            .in1(N__10925),
            .in2(N__20681),
            .in3(N__20234),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i9_3_lut_LC_12_19_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i9_3_lut_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i9_3_lut_LC_12_19_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i9_3_lut_LC_12_19_1  (
            .in0(N__19257),
            .in1(N__12938),
            .in2(_gnd_net_),
            .in3(N__12955),
            .lcout(\transmit_module.n180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i6_3_lut_4_lut_LC_12_19_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i6_3_lut_4_lut_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i6_3_lut_4_lut_LC_12_19_2 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i6_3_lut_4_lut_LC_12_19_2  (
            .in0(N__19616),
            .in1(N__12794),
            .in2(N__19737),
            .in3(N__16431),
            .lcout(\transmit_module.n215 ),
            .ltout(\transmit_module.n215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1680_4_lut_LC_12_19_3 .C_ON=1'b0;
    defparam \transmit_module.i1680_4_lut_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1680_4_lut_LC_12_19_3 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.i1680_4_lut_LC_12_19_3  (
            .in0(N__20233),
            .in1(N__20605),
            .in2(N__10424),
            .in3(N__10204),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i5_LC_12_19_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i5_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i5_LC_12_19_4 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.BRAM_ADDR__i5_LC_12_19_4  (
            .in0(N__10205),
            .in1(N__10193),
            .in2(N__20682),
            .in3(N__20235),
            .lcout(\transmit_module.TX_ADDR_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i9_3_lut_4_lut_LC_12_19_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i9_3_lut_4_lut_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i9_3_lut_4_lut_LC_12_19_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i9_3_lut_4_lut_LC_12_19_5  (
            .in0(N__19723),
            .in1(N__12956),
            .in2(N__12773),
            .in3(N__19615),
            .lcout(\transmit_module.n212 ),
            .ltout(\transmit_module.n212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i8_LC_12_19_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i8_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i8_LC_12_19_6 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \transmit_module.BRAM_ADDR__i8_LC_12_19_6  (
            .in0(N__10919),
            .in1(N__20508),
            .in2(N__10910),
            .in3(N__20236),
            .lcout(\transmit_module.TX_ADDR_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_12_20_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i8_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10907),
            .lcout(\transmit_module.X_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21786),
            .ce(N__12879),
            .sr(N__18693));
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_12_20_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_12_20_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_12_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i7_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10892),
            .lcout(\transmit_module.X_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21786),
            .ce(N__12879),
            .sr(N__18693));
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_12_20_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_12_20_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_12_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i6_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10886),
            .lcout(\transmit_module.X_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21786),
            .ce(N__12879),
            .sr(N__18693));
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_12_20_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_12_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i5_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10880),
            .lcout(\transmit_module.X_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21786),
            .ce(N__12879),
            .sr(N__18693));
    defparam \line_buffer.n3785_bdd_4_lut_LC_12_21_4 .C_ON=1'b0;
    defparam \line_buffer.n3785_bdd_4_lut_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3785_bdd_4_lut_LC_12_21_4 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n3785_bdd_4_lut_LC_12_21_4  (
            .in0(N__10874),
            .in1(N__10862),
            .in2(N__10856),
            .in3(N__22930),
            .lcout(\line_buffer.n3788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_9_0 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_9_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_9_0  (
            .in0(N__15917),
            .in1(N__15751),
            .in2(N__15855),
            .in3(N__11300),
            .lcout(\line_buffer.n577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_10_LC_13_9_1 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_10_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_10_LC_13_9_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_10_LC_13_9_1  (
            .in0(N__11298),
            .in1(N__15840),
            .in2(N__15764),
            .in3(N__15915),
            .lcout(\line_buffer.n513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i2393_2_lut_rep_18_LC_13_9_2 .C_ON=1'b0;
    defparam \receive_module.i2393_2_lut_rep_18_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.i2393_2_lut_rep_18_LC_13_9_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \receive_module.i2393_2_lut_rep_18_LC_13_9_2  (
            .in0(N__17758),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11301),
            .lcout(\receive_module.n3854 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_adj_17_LC_13_9_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_adj_17_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_adj_17_LC_13_9_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_adj_17_LC_13_9_3  (
            .in0(N__11135),
            .in1(N__11111),
            .in2(N__11105),
            .in3(N__11075),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3648_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2397_4_lut_LC_13_9_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2397_4_lut_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2397_4_lut_LC_13_9_4 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \receive_module.rx_counter.i2397_4_lut_LC_13_9_4  (
            .in0(N__11051),
            .in1(N__11045),
            .in2(N__11039),
            .in3(N__18845),
            .lcout(DEBUG_c_5),
            .ltout(DEBUG_c_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_7_LC_13_9_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_7_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_7_LC_13_9_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_7_LC_13_9_5  (
            .in0(N__15746),
            .in1(N__15839),
            .in2(N__11036),
            .in3(N__15916),
            .lcout(\line_buffer.n641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_8_LC_13_9_6 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_8_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_8_LC_13_9_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_8_LC_13_9_6  (
            .in0(N__15914),
            .in1(N__15747),
            .in2(N__15854),
            .in3(N__11299),
            .lcout(\line_buffer.n609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i0_LC_13_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i0_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i0_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_264__i0_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__13535),
            .in2(_gnd_net_),
            .in3(N__10937),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_0 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\receive_module.rx_counter.n3387 ),
            .clk(N__21010),
            .ce(N__16720),
            .sr(N__13487));
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i1_LC_13_10_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i1_LC_13_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i1_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_264__i1_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__13547),
            .in2(_gnd_net_),
            .in3(N__10934),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3387 ),
            .carryout(\receive_module.rx_counter.n3388 ),
            .clk(N__21010),
            .ce(N__16720),
            .sr(N__13487));
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i2_LC_13_10_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i2_LC_13_10_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i2_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_264__i2_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__13571),
            .in2(_gnd_net_),
            .in3(N__10931),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3388 ),
            .carryout(\receive_module.rx_counter.n3389 ),
            .clk(N__21010),
            .ce(N__16720),
            .sr(N__13487));
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i3_LC_13_10_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i3_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i3_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_264__i3_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__13523),
            .in2(_gnd_net_),
            .in3(N__10928),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3389 ),
            .carryout(\receive_module.rx_counter.n3390 ),
            .clk(N__21010),
            .ce(N__16720),
            .sr(N__13487));
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i4_LC_13_10_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i4_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i4_LC_13_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_264__i4_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__13583),
            .in2(_gnd_net_),
            .in3(N__11339),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3390 ),
            .carryout(\receive_module.rx_counter.n3391 ),
            .clk(N__21010),
            .ce(N__16720),
            .sr(N__13487));
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i5_LC_13_10_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i5_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_264__i5_LC_13_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_264__i5_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__13559),
            .in2(_gnd_net_),
            .in3(N__11336),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21010),
            .ce(N__16720),
            .sr(N__13487));
    defparam \receive_module.BRAM_ADDR__i7_LC_13_11_0 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i7_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i7_LC_13_11_0 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \receive_module.BRAM_ADDR__i7_LC_13_11_0  (
            .in0(N__14129),
            .in1(N__14105),
            .in2(N__17833),
            .in3(N__11320),
            .lcout(RX_ADDR_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21014),
            .ce(),
            .sr(N__17702));
    defparam \receive_module.BRAM_ADDR__i6_LC_13_11_1 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i6_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i6_LC_13_11_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \receive_module.BRAM_ADDR__i6_LC_13_11_1  (
            .in0(N__11317),
            .in1(N__17812),
            .in2(N__14357),
            .in3(N__14381),
            .lcout(RX_ADDR_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21014),
            .ce(),
            .sr(N__17702));
    defparam \receive_module.BRAM_ADDR__i5_LC_13_11_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i5_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i5_LC_13_11_2 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \receive_module.BRAM_ADDR__i5_LC_13_11_2  (
            .in0(N__14591),
            .in1(N__14611),
            .in2(N__17834),
            .in3(N__11319),
            .lcout(RX_ADDR_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21014),
            .ce(),
            .sr(N__17702));
    defparam \receive_module.BRAM_ADDR__i4_LC_13_11_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i4_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i4_LC_13_11_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \receive_module.BRAM_ADDR__i4_LC_13_11_3  (
            .in0(N__11316),
            .in1(N__17811),
            .in2(N__14846),
            .in3(N__14870),
            .lcout(RX_ADDR_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21014),
            .ce(),
            .sr(N__17702));
    defparam \receive_module.BRAM_ADDR__i0_LC_13_11_4 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i0_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i0_LC_13_11_4 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \receive_module.BRAM_ADDR__i0_LC_13_11_4  (
            .in0(N__13241),
            .in1(N__13268),
            .in2(N__17832),
            .in3(N__11318),
            .lcout(RX_ADDR_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21014),
            .ce(),
            .sr(N__17702));
    defparam \transmit_module.video_signal_controller.i1_3_lut_LC_13_11_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_3_lut_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_3_lut_LC_13_11_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_3_lut_LC_13_11_7  (
            .in0(N__11234),
            .in1(N__11204),
            .in2(_gnd_net_),
            .in3(N__11177),
            .lcout(\transmit_module.video_signal_controller.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1753_4_lut_LC_13_13_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1753_4_lut_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1753_4_lut_LC_13_13_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \transmit_module.video_signal_controller.i1753_4_lut_LC_13_13_0  (
            .in0(N__15660),
            .in1(N__16388),
            .in2(N__15620),
            .in3(N__15639),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3023_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_1 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_1  (
            .in0(N__16366),
            .in1(N__16345),
            .in2(N__11393),
            .in3(N__11363),
            .lcout(\transmit_module.video_signal_controller.n3577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_13_13_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_13_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__16324),
            .in2(_gnd_net_),
            .in3(N__16309),
            .lcout(\transmit_module.video_signal_controller.n3575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i487_3_lut_LC_13_13_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i487_3_lut_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i487_3_lut_LC_13_13_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \transmit_module.video_signal_controller.i487_3_lut_LC_13_13_3  (
            .in0(N__15638),
            .in1(N__15614),
            .in2(_gnd_net_),
            .in3(N__15659),
            .lcout(\transmit_module.video_signal_controller.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2335_3_lut_LC_13_13_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2335_3_lut_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2335_3_lut_LC_13_13_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2335_3_lut_LC_13_13_4  (
            .in0(N__15618),
            .in1(N__16389),
            .in2(_gnd_net_),
            .in3(N__11351),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3697_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VS_55_LC_13_13_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VS_55_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VS_55_LC_13_13_5 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VS_55_LC_13_13_5  (
            .in0(N__15640),
            .in1(N__15677),
            .in2(N__11390),
            .in3(N__15661),
            .lcout(ADV_VSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21667),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_1 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_1  (
            .in0(N__17330),
            .in1(N__11387),
            .in2(N__16397),
            .in3(N__11350),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n6_adj_568_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_13_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_13_14_2 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \transmit_module.video_signal_controller.i3_4_lut_LC_13_14_2  (
            .in0(N__16294),
            .in1(N__11381),
            .in2(N__11375),
            .in3(N__11372),
            .lcout(\transmit_module.n3549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3  (
            .in0(N__17369),
            .in1(N__17347),
            .in2(_gnd_net_),
            .in3(N__16344),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_13_14_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_13_14_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i4_4_lut_LC_13_14_4  (
            .in0(N__16293),
            .in1(N__16365),
            .in2(N__11366),
            .in3(N__11362),
            .lcout(\transmit_module.video_signal_controller.n2015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i12_LC_13_14_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i12_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i12_LC_13_14_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \transmit_module.BRAM_ADDR__i12_LC_13_14_5  (
            .in0(N__12740),
            .in1(N__16577),
            .in2(N__16496),
            .in3(N__19590),
            .lcout(TX_ADDR_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22084),
            .ce(N__17498),
            .sr(N__20366));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_16_3_lut_4_lut_LC_13_15_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_16_3_lut_4_lut_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_16_3_lut_4_lut_LC_13_15_0 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_16_3_lut_4_lut_LC_13_15_0  (
            .in0(N__12049),
            .in1(N__12023),
            .in2(N__11975),
            .in3(N__19549),
            .lcout(n3852),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i1_3_lut_4_lut_LC_13_15_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i1_3_lut_4_lut_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i1_3_lut_4_lut_LC_13_15_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i1_3_lut_4_lut_LC_13_15_1  (
            .in0(N__19548),
            .in1(N__19722),
            .in2(N__12686),
            .in3(N__16472),
            .lcout(\transmit_module.n220 ),
            .ltout(\transmit_module.n220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1670_4_lut_LC_13_15_2 .C_ON=1'b0;
    defparam \transmit_module.i1670_4_lut_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1670_4_lut_LC_13_15_2 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \transmit_module.i1670_4_lut_LC_13_15_2  (
            .in0(N__20384),
            .in1(N__16588),
            .in2(N__11957),
            .in3(N__20178),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i13_LC_13_15_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i13_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i13_LC_13_15_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \transmit_module.BRAM_ADDR__i13_LC_13_15_4  (
            .in0(N__21214),
            .in1(N__11735),
            .in2(_gnd_net_),
            .in3(N__17490),
            .lcout(DEBUG_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22077),
            .ce(),
            .sr(N__20613));
    defparam \transmit_module.video_signal_controller.mux_15_i2_3_lut_4_lut_LC_13_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i2_3_lut_4_lut_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i2_3_lut_4_lut_LC_13_15_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i2_3_lut_4_lut_LC_13_15_5  (
            .in0(N__19547),
            .in1(N__19721),
            .in2(N__12674),
            .in3(N__16544),
            .lcout(\transmit_module.n219 ),
            .ltout(\transmit_module.n219_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1676_4_lut_LC_13_15_6 .C_ON=1'b0;
    defparam \transmit_module.i1676_4_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1676_4_lut_LC_13_15_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \transmit_module.i1676_4_lut_LC_13_15_6  (
            .in0(N__20383),
            .in1(N__12728),
            .in2(N__11729),
            .in3(N__20179),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_3_lut_LC_13_15_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_3_lut_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_3_lut_LC_13_15_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_17_3_lut_LC_13_15_7  (
            .in0(N__19546),
            .in1(N__16258),
            .in2(_gnd_net_),
            .in3(N__16220),
            .lcout(\transmit_module.n3853 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ADV_R__i1_LC_13_16_0.C_ON=1'b0;
    defparam ADV_R__i1_LC_13_16_0.SEQ_MODE=4'b1000;
    defparam ADV_R__i1_LC_13_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i1_LC_13_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22169),
            .lcout(n1850),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__12290));
    defparam ADV_R__i2_LC_13_16_1.C_ON=1'b0;
    defparam ADV_R__i2_LC_13_16_1.SEQ_MODE=4'b1000;
    defparam ADV_R__i2_LC_13_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i2_LC_13_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17381),
            .lcout(n1849),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__12290));
    defparam ADV_R__i3_LC_13_16_2.C_ON=1'b0;
    defparam ADV_R__i3_LC_13_16_2.SEQ_MODE=4'b1000;
    defparam ADV_R__i3_LC_13_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i3_LC_13_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18143),
            .lcout(n1848),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__12290));
    defparam ADV_R__i4_LC_13_16_3.C_ON=1'b0;
    defparam ADV_R__i4_LC_13_16_3.SEQ_MODE=4'b1000;
    defparam ADV_R__i4_LC_13_16_3.LUT_INIT=16'b1100110011001100;
    LogicCell40 ADV_R__i4_LC_13_16_3 (
            .in0(_gnd_net_),
            .in1(N__18236),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n1847),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__12290));
    defparam ADV_R__i5_LC_13_16_4.C_ON=1'b0;
    defparam ADV_R__i5_LC_13_16_4.SEQ_MODE=4'b1000;
    defparam ADV_R__i5_LC_13_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i5_LC_13_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20759),
            .lcout(n1846),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__12290));
    defparam ADV_R__i6_LC_13_16_5.C_ON=1'b0;
    defparam ADV_R__i6_LC_13_16_5.SEQ_MODE=4'b1000;
    defparam ADV_R__i6_LC_13_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i6_LC_13_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18761),
            .lcout(n1845),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__12290));
    defparam ADV_R__i7_LC_13_16_6.C_ON=1'b0;
    defparam ADV_R__i7_LC_13_16_6.SEQ_MODE=4'b1000;
    defparam ADV_R__i7_LC_13_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i7_LC_13_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12809),
            .lcout(n1844),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__12290));
    defparam ADV_R__i8_LC_13_16_7.C_ON=1'b0;
    defparam ADV_R__i8_LC_13_16_7.SEQ_MODE=4'b1000;
    defparam ADV_R__i8_LC_13_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i8_LC_13_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18047),
            .lcout(ADV_B_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__12290));
    defparam \transmit_module.BRAM_ADDR__i0_LC_13_17_0 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i0_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i0_LC_13_17_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.BRAM_ADDR__i0_LC_13_17_0  (
            .in0(N__16595),
            .in1(N__12278),
            .in2(N__20601),
            .in3(N__20194),
            .lcout(\transmit_module.TX_ADDR_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22091),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i3_3_lut_4_lut_LC_13_17_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i3_3_lut_4_lut_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i3_3_lut_4_lut_LC_13_17_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i3_3_lut_4_lut_LC_13_17_1  (
            .in0(N__19707),
            .in1(N__16669),
            .in2(N__12656),
            .in3(N__19606),
            .lcout(\transmit_module.n218 ),
            .ltout(\transmit_module.n218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1677_4_lut_LC_13_17_2 .C_ON=1'b0;
    defparam \transmit_module.i1677_4_lut_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1677_4_lut_LC_13_17_2 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \transmit_module.i1677_4_lut_LC_13_17_2  (
            .in0(N__20490),
            .in1(N__12694),
            .in2(N__12269),
            .in3(N__20193),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i2_3_lut_LC_13_17_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i2_3_lut_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i2_3_lut_LC_13_17_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i2_3_lut_LC_13_17_3  (
            .in0(N__19226),
            .in1(N__16517),
            .in2(_gnd_net_),
            .in3(N__16539),
            .lcout(\transmit_module.n187 ),
            .ltout(\transmit_module.n187_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i1_LC_13_17_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i1_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i1_LC_13_17_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \transmit_module.BRAM_ADDR__i1_LC_13_17_4  (
            .in0(N__12716),
            .in1(N__20512),
            .in2(N__12707),
            .in3(N__20195),
            .lcout(\transmit_module.TX_ADDR_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22091),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_17_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_17_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i2_LC_13_17_5  (
            .in0(N__20196),
            .in1(N__20491),
            .in2(N__12698),
            .in3(N__12704),
            .lcout(\transmit_module.TX_ADDR_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22091),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_17_7 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i3_3_lut_LC_13_17_7  (
            .in0(N__19227),
            .in1(N__16649),
            .in2(_gnd_net_),
            .in3(N__16668),
            .lcout(\transmit_module.n186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_2_lut_LC_13_18_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_2_lut_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_2_lut_LC_13_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_2_lut_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__16463),
            .in2(N__12932),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n204 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\transmit_module.n3336 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_3_lut_LC_13_18_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_3_lut_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_3_lut_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_3_lut_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__16538),
            .in2(_gnd_net_),
            .in3(N__12659),
            .lcout(\transmit_module.n203 ),
            .ltout(),
            .carryin(\transmit_module.n3336 ),
            .carryout(\transmit_module.n3337 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_4_lut_LC_13_18_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_4_lut_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_4_lut_LC_13_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_4_lut_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__16667),
            .in2(_gnd_net_),
            .in3(N__12644),
            .lcout(\transmit_module.n202 ),
            .ltout(),
            .carryin(\transmit_module.n3337 ),
            .carryout(\transmit_module.n3338 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_5_lut_LC_13_18_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_5_lut_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_5_lut_LC_13_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_5_lut_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__19768),
            .in2(_gnd_net_),
            .in3(N__12641),
            .lcout(\transmit_module.n201 ),
            .ltout(),
            .carryin(\transmit_module.n3338 ),
            .carryout(\transmit_module.n3339 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_6_lut_LC_13_18_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_6_lut_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_6_lut_LC_13_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_6_lut_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__16619),
            .in2(_gnd_net_),
            .in3(N__12797),
            .lcout(\transmit_module.n200 ),
            .ltout(),
            .carryin(\transmit_module.n3339 ),
            .carryout(\transmit_module.n3340 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_7_lut_LC_13_18_5 .C_ON=1'b1;
    defparam \transmit_module.add_13_7_lut_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_7_lut_LC_13_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_7_lut_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__16427),
            .in2(_gnd_net_),
            .in3(N__12788),
            .lcout(\transmit_module.n199 ),
            .ltout(),
            .carryin(\transmit_module.n3340 ),
            .carryout(\transmit_module.n3341 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_8_lut_LC_13_18_6 .C_ON=1'b1;
    defparam \transmit_module.add_13_8_lut_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_8_lut_LC_13_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_8_lut_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__16700),
            .in2(_gnd_net_),
            .in3(N__12779),
            .lcout(\transmit_module.n198 ),
            .ltout(),
            .carryin(\transmit_module.n3341 ),
            .carryout(\transmit_module.n3342 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_9_lut_LC_13_18_7 .C_ON=1'b1;
    defparam \transmit_module.add_13_9_lut_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_9_lut_LC_13_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_9_lut_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__17315),
            .in2(_gnd_net_),
            .in3(N__12776),
            .lcout(\transmit_module.n197 ),
            .ltout(),
            .carryin(\transmit_module.n3342 ),
            .carryout(\transmit_module.n3343 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_10_lut_LC_13_19_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_10_lut_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_10_lut_LC_13_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_10_lut_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__12953),
            .in2(_gnd_net_),
            .in3(N__12764),
            .lcout(\transmit_module.n196 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\transmit_module.n3344 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_11_lut_LC_13_19_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_11_lut_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_11_lut_LC_13_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_11_lut_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__19634),
            .in2(_gnd_net_),
            .in3(N__12761),
            .lcout(\transmit_module.n195 ),
            .ltout(),
            .carryin(\transmit_module.n3344 ),
            .carryout(\transmit_module.n3345 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_12_lut_LC_13_19_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_12_lut_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_12_lut_LC_13_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_12_lut_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__19133),
            .in2(_gnd_net_),
            .in3(N__12758),
            .lcout(\transmit_module.n194 ),
            .ltout(),
            .carryin(\transmit_module.n3345 ),
            .carryout(\transmit_module.n3346 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_13_lut_LC_13_19_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_13_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_13_lut_LC_13_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_13_lut_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__23133),
            .in2(_gnd_net_),
            .in3(N__12743),
            .lcout(\transmit_module.n193 ),
            .ltout(),
            .carryin(\transmit_module.n3346 ),
            .carryout(\transmit_module.n3347 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_14_lut_LC_13_19_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_14_lut_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_14_lut_LC_13_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_14_lut_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__22832),
            .in2(_gnd_net_),
            .in3(N__12731),
            .lcout(\transmit_module.n192 ),
            .ltout(),
            .carryin(\transmit_module.n3347 ),
            .carryout(\transmit_module.n3348 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_15_lut_LC_13_19_5 .C_ON=1'b0;
    defparam \transmit_module.add_13_15_lut_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_15_lut_LC_13_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_15_lut_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__21257),
            .in2(_gnd_net_),
            .in3(N__12968),
            .lcout(\transmit_module.n191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_13_19_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_13_19_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i9_LC_13_19_6  (
            .in0(N__19635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21828),
            .ce(N__18466),
            .sr(N__20661));
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_13_19_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_13_19_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_13_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i8_LC_13_19_7  (
            .in0(N__12954),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21828),
            .ce(N__18466),
            .sr(N__20661));
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_13_20_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_13_20_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_13_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i0_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12911),
            .lcout(\transmit_module.X_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(N__12874),
            .sr(N__18702));
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_13_20_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_13_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i1_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12905),
            .lcout(\transmit_module.X_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(N__12874),
            .sr(N__18702));
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_13_20_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_13_20_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_13_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i2_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12887),
            .lcout(\transmit_module.X_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(N__12874),
            .sr(N__18702));
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_13_20_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_13_20_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_13_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i4_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12899),
            .lcout(\transmit_module.X_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(N__12874),
            .sr(N__18702));
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_13_20_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_13_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i3_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12893),
            .lcout(\transmit_module.X_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(N__12874),
            .sr(N__18702));
    defparam \line_buffer.dout_i6_LC_13_21_0 .C_ON=1'b0;
    defparam \line_buffer.dout_i6_LC_13_21_0 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i6_LC_13_21_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i6_LC_13_21_0  (
            .in0(N__21284),
            .in1(N__12815),
            .in2(_gnd_net_),
            .in3(N__16790),
            .lcout(TX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21686),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_VS_51_LC_14_9_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_VS_51_LC_14_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_VS_51_LC_14_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receive_module.rx_counter.old_VS_51_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17801),
            .lcout(\receive_module.rx_counter.PULSE_1HZ_N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21005),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_18_LC_14_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_18_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_18_LC_14_10_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_18_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__13582),
            .in2(_gnd_net_),
            .in3(N__13570),
            .lcout(\receive_module.rx_counter.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i140_2_lut_rep_26_LC_14_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i140_2_lut_rep_26_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i140_2_lut_rep_26_LC_14_10_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \receive_module.rx_counter.i140_2_lut_rep_26_LC_14_10_2  (
            .in0(N__13499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17773),
            .lcout(\receive_module.rx_counter.n3862 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2331_2_lut_LC_14_10_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2331_2_lut_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2331_2_lut_LC_14_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i2331_2_lut_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__13558),
            .in2(_gnd_net_),
            .in3(N__13546),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3693_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_4_lut_LC_14_10_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_4_lut_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_4_lut_LC_14_10_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \receive_module.rx_counter.i5_4_lut_LC_14_10_6  (
            .in0(N__13534),
            .in1(N__13522),
            .in2(N__13511),
            .in3(N__13508),
            .lcout(\receive_module.rx_counter.n11 ),
            .ltout(\receive_module.rx_counter.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1294_2_lut_3_lut_LC_14_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1294_2_lut_3_lut_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1294_2_lut_3_lut_LC_14_10_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \receive_module.rx_counter.i1294_2_lut_3_lut_LC_14_10_7  (
            .in0(N__17772),
            .in1(_gnd_net_),
            .in2(N__13502),
            .in3(N__13498),
            .lcout(\receive_module.rx_counter.n2562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_2_lut_LC_14_11_0 .C_ON=1'b1;
    defparam \receive_module.add_12_2_lut_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_2_lut_LC_14_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_2_lut_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__13269),
            .in2(_gnd_net_),
            .in3(N__13235),
            .lcout(\receive_module.n136 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\receive_module.n3323 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_3_lut_LC_14_11_1 .C_ON=1'b1;
    defparam \receive_module.add_12_3_lut_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_3_lut_LC_14_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_3_lut_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__13010),
            .in2(_gnd_net_),
            .in3(N__12971),
            .lcout(\receive_module.n135 ),
            .ltout(),
            .carryin(\receive_module.n3323 ),
            .carryout(\receive_module.n3324 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_4_lut_LC_14_11_2 .C_ON=1'b1;
    defparam \receive_module.add_12_4_lut_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_4_lut_LC_14_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_4_lut_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(N__15387),
            .in2(_gnd_net_),
            .in3(N__15341),
            .lcout(\receive_module.n134 ),
            .ltout(),
            .carryin(\receive_module.n3324 ),
            .carryout(\receive_module.n3325 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_5_lut_LC_14_11_3 .C_ON=1'b1;
    defparam \receive_module.add_12_5_lut_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_5_lut_LC_14_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_5_lut_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__15120),
            .in2(_gnd_net_),
            .in3(N__15080),
            .lcout(\receive_module.n133 ),
            .ltout(),
            .carryin(\receive_module.n3325 ),
            .carryout(\receive_module.n3326 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_6_lut_LC_14_11_4 .C_ON=1'b1;
    defparam \receive_module.add_12_6_lut_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_6_lut_LC_14_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_6_lut_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__14871),
            .in2(_gnd_net_),
            .in3(N__14837),
            .lcout(\receive_module.n132 ),
            .ltout(),
            .carryin(\receive_module.n3326 ),
            .carryout(\receive_module.n3327 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_7_lut_LC_14_11_5 .C_ON=1'b1;
    defparam \receive_module.add_12_7_lut_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_7_lut_LC_14_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_7_lut_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__14610),
            .in2(_gnd_net_),
            .in3(N__14585),
            .lcout(\receive_module.n131 ),
            .ltout(),
            .carryin(\receive_module.n3327 ),
            .carryout(\receive_module.n3328 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_8_lut_LC_14_11_6 .C_ON=1'b1;
    defparam \receive_module.add_12_8_lut_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_8_lut_LC_14_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_8_lut_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(N__14382),
            .in2(_gnd_net_),
            .in3(N__14348),
            .lcout(\receive_module.n130 ),
            .ltout(),
            .carryin(\receive_module.n3328 ),
            .carryout(\receive_module.n3329 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_9_lut_LC_14_11_7 .C_ON=1'b1;
    defparam \receive_module.add_12_9_lut_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_9_lut_LC_14_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_9_lut_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__14130),
            .in2(_gnd_net_),
            .in3(N__14099),
            .lcout(\receive_module.n129 ),
            .ltout(),
            .carryin(\receive_module.n3329 ),
            .carryout(\receive_module.n3330 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_10_lut_LC_14_12_0 .C_ON=1'b1;
    defparam \receive_module.add_12_10_lut_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_10_lut_LC_14_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_10_lut_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__13899),
            .in2(_gnd_net_),
            .in3(N__13841),
            .lcout(\receive_module.n128 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\receive_module.n3331 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_11_lut_LC_14_12_1 .C_ON=1'b1;
    defparam \receive_module.add_12_11_lut_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_11_lut_LC_14_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_11_lut_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__13638),
            .in2(_gnd_net_),
            .in3(N__13586),
            .lcout(\receive_module.n127 ),
            .ltout(),
            .carryin(\receive_module.n3331 ),
            .carryout(\receive_module.n3332 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_12_lut_LC_14_12_2 .C_ON=1'b1;
    defparam \receive_module.add_12_12_lut_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_12_lut_LC_14_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_12_lut_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__15975),
            .in2(_gnd_net_),
            .in3(N__15920),
            .lcout(\receive_module.n126 ),
            .ltout(),
            .carryin(\receive_module.n3332 ),
            .carryout(\receive_module.n3333 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i11_LC_14_12_3 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i11_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i11_LC_14_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i11_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__15909),
            .in2(_gnd_net_),
            .in3(N__15863),
            .lcout(RX_ADDR_11),
            .ltout(),
            .carryin(\receive_module.n3333 ),
            .carryout(\receive_module.n3334 ),
            .clk(N__21015),
            .ce(N__15785),
            .sr(N__17698));
    defparam \receive_module.BRAM_ADDR__i12_LC_14_12_4 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i12_LC_14_12_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i12_LC_14_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i12_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__15829),
            .in2(_gnd_net_),
            .in3(N__15788),
            .lcout(RX_ADDR_12),
            .ltout(),
            .carryin(\receive_module.n3334 ),
            .carryout(\receive_module.n3335 ),
            .clk(N__21015),
            .ce(N__15785),
            .sr(N__17698));
    defparam \receive_module.add_12_15_lut_LC_14_12_5 .C_ON=1'b0;
    defparam \receive_module.add_12_15_lut_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_15_lut_LC_14_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_15_lut_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(N__15766),
            .in2(_gnd_net_),
            .in3(N__15692),
            .lcout(\receive_module.n123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i0_LC_14_13_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i0_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i0_LC_14_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i0_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__15676),
            .in2(_gnd_net_),
            .in3(N__15665),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_0 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\transmit_module.video_signal_controller.n3366 ),
            .clk(N__22037),
            .ce(N__17643),
            .sr(N__17594));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i1_LC_14_13_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i1_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i1_LC_14_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i1_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__15662),
            .in2(_gnd_net_),
            .in3(N__15644),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3366 ),
            .carryout(\transmit_module.video_signal_controller.n3367 ),
            .clk(N__22037),
            .ce(N__17643),
            .sr(N__17594));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i2_LC_14_13_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i2_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i2_LC_14_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i2_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__15641),
            .in2(_gnd_net_),
            .in3(N__15623),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3367 ),
            .carryout(\transmit_module.video_signal_controller.n3368 ),
            .clk(N__22037),
            .ce(N__17643),
            .sr(N__17594));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i3_LC_14_13_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i3_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i3_LC_14_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i3_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__15619),
            .in2(_gnd_net_),
            .in3(N__15599),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3368 ),
            .carryout(\transmit_module.video_signal_controller.n3369 ),
            .clk(N__22037),
            .ce(N__17643),
            .sr(N__17594));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i4_LC_14_13_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i4_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i4_LC_14_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i4_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__16393),
            .in2(_gnd_net_),
            .in3(N__16370),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3369 ),
            .carryout(\transmit_module.video_signal_controller.n3370 ),
            .clk(N__22037),
            .ce(N__17643),
            .sr(N__17594));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i5_LC_14_13_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i5_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i5_LC_14_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i5_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__16367),
            .in2(_gnd_net_),
            .in3(N__16349),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3370 ),
            .carryout(\transmit_module.video_signal_controller.n3371 ),
            .clk(N__22037),
            .ce(N__17643),
            .sr(N__17594));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i6_LC_14_13_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i6_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i6_LC_14_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i6_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__16346),
            .in2(_gnd_net_),
            .in3(N__16328),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3371 ),
            .carryout(\transmit_module.video_signal_controller.n3372 ),
            .clk(N__22037),
            .ce(N__17643),
            .sr(N__17594));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i7_LC_14_13_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i7_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i7_LC_14_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i7_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__16325),
            .in2(_gnd_net_),
            .in3(N__16313),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3372 ),
            .carryout(\transmit_module.video_signal_controller.n3373 ),
            .clk(N__22037),
            .ce(N__17643),
            .sr(N__17594));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i8_LC_14_14_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i8_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i8_LC_14_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i8_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__16310),
            .in2(_gnd_net_),
            .in3(N__16298),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_8 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\transmit_module.video_signal_controller.n3374 ),
            .clk(N__22041),
            .ce(N__17638),
            .sr(N__17593));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i9_LC_14_14_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i9_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i9_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i9_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__16295),
            .in2(_gnd_net_),
            .in3(N__16280),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3374 ),
            .carryout(\transmit_module.video_signal_controller.n3375 ),
            .clk(N__22041),
            .ce(N__17638),
            .sr(N__17593));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i10_LC_14_14_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i10_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i10_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i10_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__17348),
            .in2(_gnd_net_),
            .in3(N__16277),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3375 ),
            .carryout(\transmit_module.video_signal_controller.n3376 ),
            .clk(N__22041),
            .ce(N__17638),
            .sr(N__17593));
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i11_LC_14_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i11_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_265__i11_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_265__i11_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__17368),
            .in2(_gnd_net_),
            .in3(N__16274),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22041),
            .ce(N__17638),
            .sr(N__17593));
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_29_LC_14_15_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_29_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_29_LC_14_15_2 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_29_LC_14_15_2  (
            .in0(N__19568),
            .in1(N__20489),
            .in2(N__16271),
            .in3(N__16228),
            .lcout(\transmit_module.n3865 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_15_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i1_3_lut_LC_14_15_3  (
            .in0(N__19221),
            .in1(N__16445),
            .in2(_gnd_net_),
            .in3(N__16471),
            .lcout(\transmit_module.n188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_14_15_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_14_15_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_14_15_7  (
            .in0(N__19222),
            .in1(N__16576),
            .in2(N__20600),
            .in3(N__19567),
            .lcout(\transmit_module.n2321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_16_1 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16543),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__18458),
            .sr(N__20686));
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_14_16_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_14_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i11_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23094),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__18458),
            .sr(N__20686));
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_16_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22926),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__18458),
            .sr(N__20686));
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_16_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21253),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__18458),
            .sr(N__20686));
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16470),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21876),
            .ce(N__18458),
            .sr(N__20686));
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16622),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(N__18459),
            .sr(N__20711));
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_1 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16439),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(N__18459),
            .sr(N__20711));
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_17_2 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16709),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(N__18459),
            .sr(N__20711));
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_17_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17318),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(N__18459),
            .sr(N__20711));
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_14_17_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_14_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i3_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19772),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(N__18459),
            .sr(N__20711));
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16670),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21908),
            .ce(N__18459),
            .sr(N__20711));
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_18_0 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_18_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_12_i8_3_lut_LC_14_18_0  (
            .in0(N__16643),
            .in1(N__19251),
            .in2(_gnd_net_),
            .in3(N__17316),
            .lcout(\transmit_module.n181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_18_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_18_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i5_3_lut_LC_14_18_1  (
            .in0(N__19250),
            .in1(N__16637),
            .in2(_gnd_net_),
            .in3(N__16620),
            .lcout(\transmit_module.n184 ),
            .ltout(\transmit_module.n184_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i4_LC_14_18_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i4_LC_14_18_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i4_LC_14_18_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i4_LC_14_18_2  (
            .in0(N__20249),
            .in1(N__20619),
            .in2(N__16631),
            .in3(N__17291),
            .lcout(\transmit_module.TX_ADDR_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21875),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i5_3_lut_4_lut_LC_14_18_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i5_3_lut_4_lut_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i5_3_lut_4_lut_LC_14_18_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i5_3_lut_4_lut_LC_14_18_3  (
            .in0(N__16628),
            .in1(N__16621),
            .in2(N__19739),
            .in3(N__19609),
            .lcout(\transmit_module.n216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i8_3_lut_4_lut_LC_14_18_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i8_3_lut_4_lut_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i8_3_lut_4_lut_LC_14_18_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i8_3_lut_4_lut_LC_14_18_5  (
            .in0(N__17317),
            .in1(N__16601),
            .in2(N__19738),
            .in3(N__19608),
            .lcout(\transmit_module.n213 ),
            .ltout(\transmit_module.n213_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_6 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i7_LC_14_18_6  (
            .in0(N__20250),
            .in1(N__20620),
            .in2(N__17321),
            .in3(N__17060),
            .lcout(\transmit_module.TX_ADDR_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21875),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_18_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_18_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.BRAM_ADDR__i9_LC_14_18_7  (
            .in0(N__20746),
            .in1(N__20732),
            .in2(N__20685),
            .in3(N__20251),
            .lcout(\transmit_module.TX_ADDR_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21875),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1679_4_lut_LC_14_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1679_4_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1679_4_lut_LC_14_19_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1679_4_lut_LC_14_19_0  (
            .in0(N__17297),
            .in1(N__17290),
            .in2(N__20701),
            .in3(N__20239),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_19_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_19_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i10_3_lut_LC_14_19_5  (
            .in0(N__19252),
            .in1(N__17066),
            .in2(_gnd_net_),
            .in3(N__19636),
            .lcout(\transmit_module.n179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1682_4_lut_LC_14_19_6 .C_ON=1'b0;
    defparam \transmit_module.i1682_4_lut_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1682_4_lut_LC_14_19_6 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1682_4_lut_LC_14_19_6  (
            .in0(N__17059),
            .in1(N__17048),
            .in2(N__20700),
            .in3(N__20240),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3767_bdd_4_lut_LC_14_21_5 .C_ON=1'b0;
    defparam \line_buffer.n3767_bdd_4_lut_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3767_bdd_4_lut_LC_14_21_5 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n3767_bdd_4_lut_LC_14_21_5  (
            .in0(N__16832),
            .in1(N__18338),
            .in2(N__16811),
            .in3(N__22907),
            .lcout(\line_buffer.n3770 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2343_3_lut_LC_15_9_0 .C_ON=1'b0;
    defparam \line_buffer.i2343_3_lut_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2343_3_lut_LC_15_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2343_3_lut_LC_15_9_0  (
            .in0(N__16784),
            .in1(N__16766),
            .in2(_gnd_net_),
            .in3(N__23125),
            .lcout(\line_buffer.n3705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__16732),
            .in2(_gnd_net_),
            .in3(N__16754),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21006),
            .ce(N__16721),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i23_1_lut_LC_15_11_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i23_1_lut_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i23_1_lut_LC_15_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \receive_module.rx_counter.i23_1_lut_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17771),
            .lcout(\receive_module.BRAM_ADDR_13__N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1289_2_lut_LC_15_13_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1289_2_lut_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1289_2_lut_LC_15_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1289_2_lut_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__17534),
            .in2(_gnd_net_),
            .in3(N__17639),
            .lcout(\transmit_module.video_signal_controller.n2551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.SYNC_BUFF1_51_LC_15_13_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.SYNC_BUFF1_51_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.SYNC_BUFF1_51_LC_15_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.video_signal_controller.SYNC_BUFF1_51_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17560),
            .lcout(\transmit_module.video_signal_controller.SYNC_BUFF1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21685),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.SYNC_BUFF2_52_LC_15_13_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.SYNC_BUFF2_52_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.SYNC_BUFF2_52_LC_15_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.video_signal_controller.SYNC_BUFF2_52_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17540),
            .lcout(\transmit_module.video_signal_controller.SYNC_BUFF2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21685),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1716_4_lut_LC_15_14_0 .C_ON=1'b0;
    defparam \transmit_module.i1716_4_lut_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1716_4_lut_LC_15_14_0 .LUT_INIT=16'b1111011111110100;
    LogicCell40 \transmit_module.i1716_4_lut_LC_15_14_0  (
            .in0(N__19258),
            .in1(N__20232),
            .in2(N__20617),
            .in3(N__17518),
            .lcout(\transmit_module.n2039 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2353_3_lut_LC_15_14_3 .C_ON=1'b0;
    defparam \line_buffer.i2353_3_lut_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2353_3_lut_LC_15_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2353_3_lut_LC_15_14_3  (
            .in0(N__17459),
            .in1(N__17441),
            .in2(_gnd_net_),
            .in3(N__23107),
            .lcout(\line_buffer.n3715 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3827_bdd_4_lut_LC_15_14_4 .C_ON=1'b0;
    defparam \line_buffer.n3827_bdd_4_lut_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3827_bdd_4_lut_LC_15_14_4 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n3827_bdd_4_lut_LC_15_14_4  (
            .in0(N__17426),
            .in1(N__18389),
            .in2(N__17405),
            .in3(N__22872),
            .lcout(),
            .ltout(\line_buffer.n3830_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i1_LC_15_14_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i1_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i1_LC_15_14_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \line_buffer.dout_i1_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__21277),
            .in2(N__17384),
            .in3(N__22703),
            .lcout(TX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21684),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_15_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_15_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__17364),
            .in2(_gnd_net_),
            .in3(N__17346),
            .lcout(\transmit_module.video_signal_controller.n3858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_15_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_15_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_15_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i38_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17996),
            .lcout(\transmit_module.Y_DELTA_PATTERN_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(N__17913),
            .sr(N__20683));
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_15_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_15_15_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_15_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i37_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18035),
            .lcout(\transmit_module.Y_DELTA_PATTERN_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(N__17913),
            .sr(N__20683));
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_15_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_15_15_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_15_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i35_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18017),
            .lcout(\transmit_module.Y_DELTA_PATTERN_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(N__17913),
            .sr(N__20683));
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_15_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_15_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_15_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i34_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18029),
            .lcout(\transmit_module.Y_DELTA_PATTERN_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(N__17913),
            .sr(N__20683));
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_15_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_15_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i36_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18023),
            .lcout(\transmit_module.Y_DELTA_PATTERN_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(N__17913),
            .sr(N__20683));
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_15_15_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_15_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i39_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18011),
            .lcout(\transmit_module.Y_DELTA_PATTERN_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(N__17913),
            .sr(N__20683));
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_15_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_15_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_15_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i33_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17990),
            .lcout(\transmit_module.Y_DELTA_PATTERN_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(N__17913),
            .sr(N__20683));
    defparam \line_buffer.n3779_bdd_4_lut_LC_15_16_2 .C_ON=1'b0;
    defparam \line_buffer.n3779_bdd_4_lut_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3779_bdd_4_lut_LC_15_16_2 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.n3779_bdd_4_lut_LC_15_16_2  (
            .in0(N__22921),
            .in1(N__17885),
            .in2(N__17870),
            .in3(N__18065),
            .lcout(\line_buffer.n3782 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2425_LC_15_16_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2425_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2425_LC_15_16_3 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2425_LC_15_16_3  (
            .in0(N__18110),
            .in1(N__17849),
            .in2(N__21289),
            .in3(N__22919),
            .lcout(),
            .ltout(\line_buffer.n3773_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i3_LC_15_16_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i3_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i3_LC_15_16_4 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.dout_i3_LC_15_16_4  (
            .in0(N__18299),
            .in1(N__18248),
            .in2(N__18239),
            .in3(N__21272),
            .lcout(TX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21559),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2440_LC_15_16_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2440_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2440_LC_15_16_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2440_LC_15_16_5  (
            .in0(N__18227),
            .in1(N__22918),
            .in2(N__18215),
            .in3(N__23093),
            .lcout(),
            .ltout(\line_buffer.n3803_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3803_bdd_4_lut_LC_15_16_6 .C_ON=1'b0;
    defparam \line_buffer.n3803_bdd_4_lut_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3803_bdd_4_lut_LC_15_16_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.n3803_bdd_4_lut_LC_15_16_6  (
            .in0(N__22920),
            .in1(N__18194),
            .in2(N__18173),
            .in3(N__18170),
            .lcout(),
            .ltout(\line_buffer.n3806_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i2_LC_15_16_7 .C_ON=1'b0;
    defparam \line_buffer.dout_i2_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i2_LC_15_16_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \line_buffer.dout_i2_LC_15_16_7  (
            .in0(N__21271),
            .in1(_gnd_net_),
            .in2(N__18152),
            .in3(N__18149),
            .lcout(TX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21559),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2344_3_lut_LC_15_17_1 .C_ON=1'b0;
    defparam \line_buffer.i2344_3_lut_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2344_3_lut_LC_15_17_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2344_3_lut_LC_15_17_1  (
            .in0(N__18134),
            .in1(N__18125),
            .in2(_gnd_net_),
            .in3(N__23091),
            .lcout(\line_buffer.n3706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2420_LC_15_17_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2420_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2420_LC_15_17_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2420_LC_15_17_5  (
            .in0(N__18104),
            .in1(N__22908),
            .in2(N__18083),
            .in3(N__23090),
            .lcout(\line_buffer.n3779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2430_LC_15_18_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2430_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2430_LC_15_18_0 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2430_LC_15_18_0  (
            .in0(N__18059),
            .in1(N__18479),
            .in2(N__21290),
            .in3(N__22925),
            .lcout(),
            .ltout(\line_buffer.n3791_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i7_LC_15_18_1 .C_ON=1'b0;
    defparam \line_buffer.dout_i7_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i7_LC_15_18_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \line_buffer.dout_i7_LC_15_18_1  (
            .in0(N__18533),
            .in1(N__21276),
            .in2(N__18050),
            .in3(N__18260),
            .lcout(TX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21558),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2340_3_lut_LC_15_18_2 .C_ON=1'b0;
    defparam \line_buffer.i2340_3_lut_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2340_3_lut_LC_15_18_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2340_3_lut_LC_15_18_2  (
            .in0(N__18515),
            .in1(N__18500),
            .in2(_gnd_net_),
            .in3(N__23092),
            .lcout(\line_buffer.n3702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_18_7 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i4_3_lut_LC_15_18_7  (
            .in0(N__19259),
            .in1(N__18473),
            .in2(_gnd_net_),
            .in3(N__19763),
            .lcout(\transmit_module.n185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_15_19_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_15_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i10_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19128),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21827),
            .ce(N__18467),
            .sr(N__20618));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2460_LC_15_20_7 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2460_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2460_LC_15_20_7 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2460_LC_15_20_7  (
            .in0(N__18428),
            .in1(N__22934),
            .in2(N__18407),
            .in3(N__23130),
            .lcout(\line_buffer.n3827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2415_LC_15_21_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2415_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2415_LC_15_21_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2415_LC_15_21_6  (
            .in0(N__18377),
            .in1(N__22928),
            .in2(N__18356),
            .in3(N__23131),
            .lcout(\line_buffer.n3767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2352_3_lut_LC_15_22_3 .C_ON=1'b0;
    defparam \line_buffer.i2352_3_lut_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2352_3_lut_LC_15_22_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2352_3_lut_LC_15_22_3  (
            .in0(N__18332),
            .in1(N__18317),
            .in2(_gnd_net_),
            .in3(N__23129),
            .lcout(\line_buffer.n3714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2355_3_lut_LC_15_25_4 .C_ON=1'b0;
    defparam \line_buffer.i2355_3_lut_LC_15_25_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2355_3_lut_LC_15_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2355_3_lut_LC_15_25_4  (
            .in0(N__18287),
            .in1(N__18275),
            .in2(_gnd_net_),
            .in3(N__23143),
            .lcout(\line_buffer.n3717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_LC_16_9_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_LC_16_9_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_LC_16_9_0  (
            .in0(N__19852),
            .in1(N__19822),
            .in2(_gnd_net_),
            .in3(N__19837),
            .lcout(\receive_module.rx_counter.n3547 ),
            .ltout(\receive_module.rx_counter.n3547_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2251_3_lut_LC_16_9_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2251_3_lut_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2251_3_lut_LC_16_9_1 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \receive_module.rx_counter.i2251_3_lut_LC_16_9_1  (
            .in0(N__19807),
            .in1(_gnd_net_),
            .in2(N__18863),
            .in3(N__21097),
            .lcout(\receive_module.rx_counter.n3613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_adj_15_LC_16_9_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_adj_15_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_adj_15_LC_16_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_adj_15_LC_16_9_4  (
            .in0(N__21096),
            .in1(N__19806),
            .in2(_gnd_net_),
            .in3(N__18860),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3646_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i35_4_lut_LC_16_9_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i35_4_lut_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i35_4_lut_LC_16_9_5 .LUT_INIT=16'b1010100010111001;
    LogicCell40 \receive_module.rx_counter.i35_4_lut_LC_16_9_5  (
            .in0(N__21061),
            .in1(N__21079),
            .in2(N__18854),
            .in3(N__18851),
            .lcout(\receive_module.rx_counter.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2406_LC_16_13_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2406_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2406_LC_16_13_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2406_LC_16_13_6  (
            .in0(N__18836),
            .in1(N__22896),
            .in2(N__18818),
            .in3(N__23118),
            .lcout(),
            .ltout(\line_buffer.n3761_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3761_bdd_4_lut_LC_16_13_7 .C_ON=1'b0;
    defparam \line_buffer.n3761_bdd_4_lut_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3761_bdd_4_lut_LC_16_13_7 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.n3761_bdd_4_lut_LC_16_13_7  (
            .in0(N__22897),
            .in1(N__18806),
            .in2(N__18788),
            .in3(N__18785),
            .lcout(\line_buffer.n3764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i5_LC_16_14_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i5_LC_16_14_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i5_LC_16_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i5_LC_16_14_4  (
            .in0(N__21261),
            .in1(N__18767),
            .in2(_gnd_net_),
            .in3(N__20774),
            .lcout(TX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21683),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_16_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_16_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_16_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i32_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18749),
            .lcout(\transmit_module.Y_DELTA_PATTERN_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21479),
            .ce(N__18708),
            .sr(N__20577));
    defparam \line_buffer.i2356_3_lut_LC_16_17_4 .C_ON=1'b0;
    defparam \line_buffer.i2356_3_lut_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2356_3_lut_LC_16_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2356_3_lut_LC_16_17_4  (
            .in0(N__18569),
            .in1(N__18551),
            .in2(_gnd_net_),
            .in3(N__23117),
            .lcout(\line_buffer.n3718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i11_3_lut_4_lut_LC_16_18_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i11_3_lut_4_lut_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i11_3_lut_4_lut_LC_16_18_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i11_3_lut_4_lut_LC_16_18_3  (
            .in0(N__19730),
            .in1(N__18527),
            .in2(N__19132),
            .in3(N__19593),
            .lcout(\transmit_module.n210 ),
            .ltout(\transmit_module.n210_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i10_LC_16_18_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i10_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i10_LC_16_18_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \transmit_module.BRAM_ADDR__i10_LC_16_18_4  (
            .in0(N__19100),
            .in1(N__20598),
            .in2(N__19790),
            .in3(N__20237),
            .lcout(\transmit_module.TX_ADDR_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21557),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i4_3_lut_4_lut_LC_16_18_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i4_3_lut_4_lut_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i4_3_lut_4_lut_LC_16_18_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i4_3_lut_4_lut_LC_16_18_5  (
            .in0(N__19728),
            .in1(N__19764),
            .in2(N__19787),
            .in3(N__19591),
            .lcout(\transmit_module.n217 ),
            .ltout(\transmit_module.n217_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i3_LC_16_18_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i3_LC_16_18_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i3_LC_16_18_6 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \transmit_module.BRAM_ADDR__i3_LC_16_18_6  (
            .in0(N__19490),
            .in1(N__20599),
            .in2(N__19775),
            .in3(N__20238),
            .lcout(\transmit_module.TX_ADDR_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21557),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_15_i10_3_lut_4_lut_LC_16_18_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_15_i10_3_lut_4_lut_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_15_i10_3_lut_4_lut_LC_16_18_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \transmit_module.video_signal_controller.mux_15_i10_3_lut_4_lut_LC_16_18_7  (
            .in0(N__19729),
            .in1(N__19658),
            .in2(N__19646),
            .in3(N__19592),
            .lcout(\transmit_module.n211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1678_4_lut_LC_16_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1678_4_lut_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1678_4_lut_LC_16_19_0 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \transmit_module.i1678_4_lut_LC_16_19_0  (
            .in0(N__19496),
            .in1(N__19489),
            .in2(N__20666),
            .in3(N__20253),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i11_3_lut_LC_16_19_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i11_3_lut_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i11_3_lut_LC_16_19_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i11_3_lut_LC_16_19_3  (
            .in0(N__19245),
            .in1(N__19139),
            .in2(_gnd_net_),
            .in3(N__19127),
            .lcout(\transmit_module.n178 ),
            .ltout(\transmit_module.n178_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1685_4_lut_LC_16_19_4 .C_ON=1'b0;
    defparam \transmit_module.i1685_4_lut_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1685_4_lut_LC_16_19_4 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \transmit_module.i1685_4_lut_LC_16_19_4  (
            .in0(N__20587),
            .in1(N__19094),
            .in2(N__19088),
            .in3(N__20254),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_6.C_ON=1'b0;
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_6 (
            .in0(N__21050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_TVP_CLK_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i26_1_lut_rep_24_LC_17_8_3.C_ON=1'b0;
    defparam i26_1_lut_rep_24_LC_17_8_3.SEQ_MODE=4'b0000;
    defparam i26_1_lut_rep_24_LC_17_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 i26_1_lut_rep_24_LC_17_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19906),
            .lcout(n3860),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.X_263__i0_LC_17_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i0_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i0_LC_17_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i0_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__19880),
            .in2(_gnd_net_),
            .in3(N__19874),
            .lcout(\receive_module.rx_counter.n10 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\receive_module.rx_counter.n3357 ),
            .clk(N__21000),
            .ce(),
            .sr(N__20899));
    defparam \receive_module.rx_counter.X_263__i1_LC_17_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i1_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i1_LC_17_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i1_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__19871),
            .in2(_gnd_net_),
            .in3(N__19865),
            .lcout(\receive_module.rx_counter.n9 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3357 ),
            .carryout(\receive_module.rx_counter.n3358 ),
            .clk(N__21000),
            .ce(),
            .sr(N__20899));
    defparam \receive_module.rx_counter.X_263__i2_LC_17_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i2_LC_17_9_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i2_LC_17_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i2_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__19862),
            .in2(_gnd_net_),
            .in3(N__19856),
            .lcout(\receive_module.rx_counter.n8 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3358 ),
            .carryout(\receive_module.rx_counter.n3359 ),
            .clk(N__21000),
            .ce(),
            .sr(N__20899));
    defparam \receive_module.rx_counter.X_263__i3_LC_17_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i3_LC_17_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i3_LC_17_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i3_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__19853),
            .in2(_gnd_net_),
            .in3(N__19841),
            .lcout(\receive_module.rx_counter.X_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3359 ),
            .carryout(\receive_module.rx_counter.n3360 ),
            .clk(N__21000),
            .ce(),
            .sr(N__20899));
    defparam \receive_module.rx_counter.X_263__i4_LC_17_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i4_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i4_LC_17_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i4_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__19838),
            .in2(_gnd_net_),
            .in3(N__19826),
            .lcout(\receive_module.rx_counter.X_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3360 ),
            .carryout(\receive_module.rx_counter.n3361 ),
            .clk(N__21000),
            .ce(),
            .sr(N__20899));
    defparam \receive_module.rx_counter.X_263__i5_LC_17_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i5_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i5_LC_17_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i5_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(N__19823),
            .in2(_gnd_net_),
            .in3(N__19811),
            .lcout(\receive_module.rx_counter.X_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3361 ),
            .carryout(\receive_module.rx_counter.n3362 ),
            .clk(N__21000),
            .ce(),
            .sr(N__20899));
    defparam \receive_module.rx_counter.X_263__i6_LC_17_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i6_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i6_LC_17_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i6_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__19808),
            .in2(_gnd_net_),
            .in3(N__19793),
            .lcout(\receive_module.rx_counter.X_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3362 ),
            .carryout(\receive_module.rx_counter.n3363 ),
            .clk(N__21000),
            .ce(),
            .sr(N__20899));
    defparam \receive_module.rx_counter.X_263__i7_LC_17_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i7_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i7_LC_17_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i7_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(N__21098),
            .in2(_gnd_net_),
            .in3(N__21083),
            .lcout(\receive_module.rx_counter.X_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3363 ),
            .carryout(\receive_module.rx_counter.n3364 ),
            .clk(N__21000),
            .ce(),
            .sr(N__20899));
    defparam \receive_module.rx_counter.X_263__i8_LC_17_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_263__i8_LC_17_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i8_LC_17_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i8_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__21080),
            .in2(_gnd_net_),
            .in3(N__21068),
            .lcout(\receive_module.rx_counter.X_8 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\receive_module.rx_counter.n3365 ),
            .clk(N__21002),
            .ce(),
            .sr(N__20903));
    defparam \receive_module.rx_counter.X_263__i9_LC_17_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.X_263__i9_LC_17_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_263__i9_LC_17_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_263__i9_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__21062),
            .in2(_gnd_net_),
            .in3(N__21065),
            .lcout(\receive_module.rx_counter.X_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21002),
            .ce(),
            .sr(N__20903));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_13_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_13_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_13_1  (
            .in0(N__20882),
            .in1(N__22892),
            .in2(N__20873),
            .in3(N__23136),
            .lcout(\line_buffer.n3833 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2359_3_lut_LC_17_13_7 .C_ON=1'b0;
    defparam \line_buffer.i2359_3_lut_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2359_3_lut_LC_17_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2359_3_lut_LC_17_13_7  (
            .in0(N__20852),
            .in1(N__20834),
            .in2(_gnd_net_),
            .in3(N__23137),
            .lcout(\line_buffer.n3721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3833_bdd_4_lut_LC_17_14_7 .C_ON=1'b0;
    defparam \line_buffer.n3833_bdd_4_lut_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3833_bdd_4_lut_LC_17_14_7 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n3833_bdd_4_lut_LC_17_14_7  (
            .in0(N__20822),
            .in1(N__20804),
            .in2(N__20798),
            .in3(N__22866),
            .lcout(\line_buffer.n3836 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i4_LC_17_17_2 .C_ON=1'b0;
    defparam \line_buffer.dout_i4_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i4_LC_17_17_2 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.dout_i4_LC_17_17_2  (
            .in0(N__20768),
            .in1(N__21288),
            .in2(N__22340),
            .in3(N__21155),
            .lcout(TX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21966),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1684_4_lut_LC_17_19_4 .C_ON=1'b0;
    defparam \transmit_module.i1684_4_lut_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1684_4_lut_LC_17_19_4 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1684_4_lut_LC_17_19_4  (
            .in0(N__20747),
            .in1(N__20728),
            .in2(N__20665),
            .in3(N__20255),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2358_3_lut_LC_17_20_4 .C_ON=1'b0;
    defparam \line_buffer.i2358_3_lut_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2358_3_lut_LC_17_20_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2358_3_lut_LC_17_20_4  (
            .in0(N__22367),
            .in1(N__22358),
            .in2(_gnd_net_),
            .in3(N__23144),
            .lcout(\line_buffer.n3720 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2450_LC_18_15_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2450_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2450_LC_18_15_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2450_LC_18_15_2  (
            .in0(N__22328),
            .in1(N__22927),
            .in2(N__22313),
            .in3(N__23106),
            .lcout(\line_buffer.n3815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2337_3_lut_LC_19_9_5 .C_ON=1'b0;
    defparam \line_buffer.i2337_3_lut_LC_19_9_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2337_3_lut_LC_19_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2337_3_lut_LC_19_9_5  (
            .in0(N__22292),
            .in1(N__22277),
            .in2(_gnd_net_),
            .in3(N__23141),
            .lcout(\line_buffer.n3699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3815_bdd_4_lut_LC_19_15_1 .C_ON=1'b0;
    defparam \line_buffer.n3815_bdd_4_lut_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3815_bdd_4_lut_LC_19_15_1 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n3815_bdd_4_lut_LC_19_15_1  (
            .in0(N__22262),
            .in1(N__22241),
            .in2(N__22235),
            .in3(N__22932),
            .lcout(\line_buffer.n3818 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3821_bdd_4_lut_LC_19_16_4 .C_ON=1'b0;
    defparam \line_buffer.n3821_bdd_4_lut_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3821_bdd_4_lut_LC_19_16_4 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n3821_bdd_4_lut_LC_19_16_4  (
            .in0(N__22211),
            .in1(N__23183),
            .in2(N__22196),
            .in3(N__22933),
            .lcout(),
            .ltout(\line_buffer.n3824_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i0_LC_19_16_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i0_LC_19_16_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i0_LC_19_16_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \line_buffer.dout_i0_LC_19_16_5  (
            .in0(_gnd_net_),
            .in1(N__21291),
            .in2(N__22178),
            .in3(N__22175),
            .lcout(TX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21924),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_19_17_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_19_17_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_LC_19_17_1  (
            .in0(N__21107),
            .in1(N__21308),
            .in2(N__21295),
            .in3(N__22931),
            .lcout(\line_buffer.n3797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2338_3_lut_LC_19_19_1 .C_ON=1'b0;
    defparam \line_buffer.i2338_3_lut_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2338_3_lut_LC_19_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2338_3_lut_LC_19_19_1  (
            .in0(N__21146),
            .in1(N__21128),
            .in2(_gnd_net_),
            .in3(N__23134),
            .lcout(\line_buffer.n3700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2455_LC_19_19_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2455_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2455_LC_19_19_4 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2455_LC_19_19_4  (
            .in0(N__23135),
            .in1(N__23222),
            .in2(N__23201),
            .in3(N__22891),
            .lcout(\line_buffer.n3821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2445_LC_20_14_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2445_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2445_LC_20_14_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2445_LC_20_14_0  (
            .in0(N__23174),
            .in1(N__22864),
            .in2(N__23159),
            .in3(N__23142),
            .lcout(),
            .ltout(\line_buffer.n3809_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3809_bdd_4_lut_LC_20_14_1 .C_ON=1'b0;
    defparam \line_buffer.n3809_bdd_4_lut_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3809_bdd_4_lut_LC_20_14_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.n3809_bdd_4_lut_LC_20_14_1  (
            .in0(N__22865),
            .in1(N__22742),
            .in2(N__22724),
            .in3(N__22721),
            .lcout(\line_buffer.n3812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_24_31_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_24_31_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_24_31_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_24_31_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // main
