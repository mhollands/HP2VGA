// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 9 2018 04:44:33

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "RAM" view "INTERFACE"

module RAM (
    raddr,
    waddr,
    dout,
    din,
    rclk,
    wclk,
    write_en);

    input [13:0] raddr;
    input [13:0] waddr;
    output [7:0] dout;
    input [7:0] din;
    input rclk;
    input wclk;
    input write_en;

    wire N__13191;
    wire N__13190;
    wire N__13189;
    wire N__13181;
    wire N__13180;
    wire N__13179;
    wire N__13170;
    wire N__13169;
    wire N__13168;
    wire N__13161;
    wire N__13160;
    wire N__13159;
    wire N__13152;
    wire N__13151;
    wire N__13150;
    wire N__13143;
    wire N__13142;
    wire N__13141;
    wire N__13134;
    wire N__13133;
    wire N__13132;
    wire N__13125;
    wire N__13124;
    wire N__13123;
    wire N__13116;
    wire N__13115;
    wire N__13114;
    wire N__13107;
    wire N__13106;
    wire N__13105;
    wire N__13098;
    wire N__13097;
    wire N__13096;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13080;
    wire N__13079;
    wire N__13078;
    wire N__13071;
    wire N__13070;
    wire N__13069;
    wire N__13062;
    wire N__13061;
    wire N__13060;
    wire N__13053;
    wire N__13052;
    wire N__13051;
    wire N__13044;
    wire N__13043;
    wire N__13042;
    wire N__13035;
    wire N__13034;
    wire N__13033;
    wire N__13026;
    wire N__13025;
    wire N__13024;
    wire N__13017;
    wire N__13016;
    wire N__13015;
    wire N__13008;
    wire N__13007;
    wire N__13006;
    wire N__12999;
    wire N__12998;
    wire N__12997;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12981;
    wire N__12980;
    wire N__12979;
    wire N__12972;
    wire N__12971;
    wire N__12970;
    wire N__12963;
    wire N__12962;
    wire N__12961;
    wire N__12954;
    wire N__12953;
    wire N__12952;
    wire N__12945;
    wire N__12944;
    wire N__12943;
    wire N__12936;
    wire N__12935;
    wire N__12934;
    wire N__12927;
    wire N__12926;
    wire N__12925;
    wire N__12918;
    wire N__12917;
    wire N__12916;
    wire N__12909;
    wire N__12908;
    wire N__12907;
    wire N__12900;
    wire N__12899;
    wire N__12898;
    wire N__12891;
    wire N__12890;
    wire N__12889;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12873;
    wire N__12872;
    wire N__12871;
    wire N__12864;
    wire N__12863;
    wire N__12862;
    wire N__12855;
    wire N__12854;
    wire N__12853;
    wire N__12846;
    wire N__12845;
    wire N__12844;
    wire N__12837;
    wire N__12836;
    wire N__12835;
    wire N__12828;
    wire N__12827;
    wire N__12826;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12810;
    wire N__12809;
    wire N__12808;
    wire N__12801;
    wire N__12800;
    wire N__12799;
    wire N__12792;
    wire N__12791;
    wire N__12790;
    wire N__12783;
    wire N__12782;
    wire N__12781;
    wire N__12774;
    wire N__12773;
    wire N__12772;
    wire N__12755;
    wire N__12752;
    wire N__12751;
    wire N__12750;
    wire N__12749;
    wire N__12748;
    wire N__12747;
    wire N__12744;
    wire N__12739;
    wire N__12736;
    wire N__12731;
    wire N__12730;
    wire N__12729;
    wire N__12728;
    wire N__12719;
    wire N__12716;
    wire N__12715;
    wire N__12714;
    wire N__12713;
    wire N__12712;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12684;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12667;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12651;
    wire N__12648;
    wire N__12645;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12598;
    wire N__12593;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12580;
    wire N__12579;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12567;
    wire N__12566;
    wire N__12561;
    wire N__12560;
    wire N__12559;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12546;
    wire N__12543;
    wire N__12540;
    wire N__12535;
    wire N__12532;
    wire N__12529;
    wire N__12524;
    wire N__12521;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12493;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12430;
    wire N__12425;
    wire N__12424;
    wire N__12423;
    wire N__12420;
    wire N__12415;
    wire N__12414;
    wire N__12413;
    wire N__12408;
    wire N__12403;
    wire N__12402;
    wire N__12401;
    wire N__12400;
    wire N__12399;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12384;
    wire N__12381;
    wire N__12376;
    wire N__12369;
    wire N__12366;
    wire N__12365;
    wire N__12364;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12350;
    wire N__12349;
    wire N__12346;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12335;
    wire N__12330;
    wire N__12329;
    wire N__12328;
    wire N__12327;
    wire N__12322;
    wire N__12321;
    wire N__12320;
    wire N__12315;
    wire N__12314;
    wire N__12313;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12290;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12280;
    wire N__12279;
    wire N__12278;
    wire N__12275;
    wire N__12270;
    wire N__12265;
    wire N__12264;
    wire N__12263;
    wire N__12258;
    wire N__12253;
    wire N__12248;
    wire N__12245;
    wire N__12240;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12192;
    wire N__12189;
    wire N__12186;
    wire N__12183;
    wire N__12178;
    wire N__12175;
    wire N__12170;
    wire N__12165;
    wire N__12160;
    wire N__12155;
    wire N__12150;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11864;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11714;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11690;
    wire N__11687;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11423;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10999;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10991;
    wire N__10990;
    wire N__10987;
    wire N__10986;
    wire N__10985;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10964;
    wire N__10963;
    wire N__10962;
    wire N__10961;
    wire N__10960;
    wire N__10953;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10933;
    wire N__10932;
    wire N__10931;
    wire N__10928;
    wire N__10927;
    wire N__10926;
    wire N__10925;
    wire N__10924;
    wire N__10923;
    wire N__10922;
    wire N__10921;
    wire N__10920;
    wire N__10911;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10899;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10878;
    wire N__10877;
    wire N__10876;
    wire N__10873;
    wire N__10870;
    wire N__10869;
    wire N__10868;
    wire N__10865;
    wire N__10864;
    wire N__10863;
    wire N__10862;
    wire N__10859;
    wire N__10858;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10842;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10828;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10816;
    wire N__10813;
    wire N__10812;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10786;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10770;
    wire N__10767;
    wire N__10760;
    wire N__10757;
    wire N__10750;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10740;
    wire N__10737;
    wire N__10736;
    wire N__10727;
    wire N__10724;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10710;
    wire N__10709;
    wire N__10706;
    wire N__10705;
    wire N__10704;
    wire N__10703;
    wire N__10696;
    wire N__10687;
    wire N__10678;
    wire N__10675;
    wire N__10672;
    wire N__10669;
    wire N__10664;
    wire N__10657;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10641;
    wire N__10640;
    wire N__10639;
    wire N__10638;
    wire N__10637;
    wire N__10636;
    wire N__10633;
    wire N__10632;
    wire N__10631;
    wire N__10624;
    wire N__10617;
    wire N__10608;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10594;
    wire N__10591;
    wire N__10590;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10480;
    wire N__10475;
    wire N__10472;
    wire N__10465;
    wire N__10460;
    wire N__10455;
    wire N__10452;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10301;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10289;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10281;
    wire N__10276;
    wire N__10273;
    wire N__10272;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10247;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10239;
    wire N__10238;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10198;
    wire N__10197;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10173;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10148;
    wire N__10145;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10137;
    wire N__10136;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10099;
    wire N__10098;
    wire N__10097;
    wire N__10096;
    wire N__10095;
    wire N__10094;
    wire N__10093;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10063;
    wire N__10062;
    wire N__10061;
    wire N__10060;
    wire N__10059;
    wire N__10058;
    wire N__10057;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10027;
    wire N__10026;
    wire N__10025;
    wire N__10022;
    wire N__10021;
    wire N__10018;
    wire N__10017;
    wire N__10014;
    wire N__10013;
    wire N__10010;
    wire N__10009;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9977;
    wire N__9976;
    wire N__9973;
    wire N__9972;
    wire N__9969;
    wire N__9968;
    wire N__9965;
    wire N__9964;
    wire N__9961;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9918;
    wire N__9913;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9598;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9587;
    wire N__9580;
    wire N__9577;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9542;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9517;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9487;
    wire N__9484;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9431;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8771;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8764;
    wire N__8763;
    wire N__8762;
    wire N__8761;
    wire N__8760;
    wire N__8759;
    wire N__8758;
    wire N__8757;
    wire N__8756;
    wire N__8755;
    wire N__8754;
    wire N__8753;
    wire N__8752;
    wire N__8751;
    wire N__8750;
    wire N__8749;
    wire N__8748;
    wire N__8747;
    wire N__8746;
    wire N__8745;
    wire N__8744;
    wire N__8743;
    wire N__8742;
    wire N__8741;
    wire N__8740;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8638;
    wire N__8635;
    wire N__8632;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8491;
    wire N__8488;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8015;
    wire N__8014;
    wire N__8013;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8005;
    wire N__8004;
    wire N__8003;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7987;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7972;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7941;
    wire N__7936;
    wire N__7933;
    wire N__7930;
    wire N__7927;
    wire N__7924;
    wire N__7917;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7882;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7831;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7756;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7741;
    wire N__7738;
    wire N__7735;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7708;
    wire N__7705;
    wire N__7702;
    wire N__7699;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7660;
    wire N__7657;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7618;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7519;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7462;
    wire N__7459;
    wire N__7456;
    wire N__7453;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7253;
    wire N__7250;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6982;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6799;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6736;
    wire N__6733;
    wire N__6730;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5948;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5040;
    wire N__5037;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5019;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5000;
    wire N__4997;
    wire N__4992;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4973;
    wire N__4970;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4951;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4934;
    wire N__4933;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4929;
    wire N__4928;
    wire N__4927;
    wire N__4926;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4921;
    wire N__4920;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4913;
    wire N__4912;
    wire N__4911;
    wire N__4910;
    wire N__4909;
    wire N__4908;
    wire N__4907;
    wire N__4906;
    wire N__4905;
    wire N__4904;
    wire N__4903;
    wire N__4902;
    wire N__4901;
    wire N__4900;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4372;
    wire N__4369;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4355;
    wire N__4350;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4330;
    wire N__4325;
    wire N__4324;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4303;
    wire N__4298;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4262;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4251;
    wire N__4248;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4229;
    wire N__4228;
    wire N__4225;
    wire N__4220;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4199;
    wire N__4196;
    wire N__4191;
    wire N__4190;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4147;
    wire N__4146;
    wire N__4145;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4131;
    wire N__4128;
    wire N__4123;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4103;
    wire N__4100;
    wire N__4095;
    wire N__4092;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4059;
    wire N__4054;
    wire N__4051;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4028;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4016;
    wire N__4015;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4007;
    wire N__4004;
    wire N__3999;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3964;
    wire N__3961;
    wire N__3958;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3925;
    wire N__3922;
    wire N__3919;
    wire N__3914;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3906;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3891;
    wire N__3890;
    wire N__3885;
    wire N__3882;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3844;
    wire GNDG0;
    wire din_c_3;
    wire din_c_2;
    wire VCCG0;
    wire din_c_6;
    wire din_c_7;
    wire din_c_4;
    wire din_c_5;
    wire raddr_c_5;
    wire waddr_c_3;
    wire waddr_c_6;
    wire wclk_c_g;
    wire raddr_c_2;
    wire raddr_c_7;
    wire waddr_c_5;
    wire din_c_1;
    wire raddr_c_8;
    wire waddr_c_4;
    wire raddr_c_10;
    wire raddr_c_4;
    wire waddr_c_9;
    wire raddr_c_9;
    wire waddr_c_7;
    wire raddr_c_0;
    wire waddr_c_10;
    wire waddr_c_8;
    wire raddr_c_1;
    wire raddr_c_6;
    wire waddr_c_2;
    wire din_c_0;
    wire rclk_c_g;
    wire raddr_c_3;
    wire waddr_c_1;
    wire waddr_c_0;
    wire mem_WE_4;
    wire mem_WE_0;
    wire mem_WE_8;
    wire mem_WE_12;
    wire mem_WE_16;
    wire mem_WE_20;
    wire mem_WE_24;
    wire write_en_c;
    wire waddr_c_13;
    wire waddr_c_11;
    wire waddr_c_12;
    wire mem_WE_28;
    wire mem_out_bus0_0;
    wire mem_out_bus4_0;
    wire mem_out_bus0_1;
    wire mem_out_bus4_1;
    wire mem_out_bus4_7;
    wire mem_out_bus0_7;
    wire mem_out_bus0_6;
    wire mem_out_bus4_6;
    wire CONSTANT_ONE_NET;
    wire mem_out_bus5_1;
    wire mem_out_bus1_1;
    wire mem_out_bus5_0;
    wire mem_out_bus1_0;
    wire dout_obuf_RNO_4Z0Z_1;
    wire mem_N_162_cascade_;
    wire dout_c_1;
    wire dout_obuf_RNO_4Z0Z_0;
    wire mem_N_156_cascade_;
    wire dout_c_0;
    wire dout_obuf_RNO_2Z0Z_1;
    wire mem_N_160;
    wire dout_obuf_RNO_2Z0Z_0;
    wire mem_N_154;
    wire mem_out_bus5_2;
    wire mem_out_bus1_2;
    wire dout_obuf_RNO_2Z0Z_2;
    wire mem_N_166_cascade_;
    wire dout_c_2;
    wire dout_obuf_RNO_4Z0Z_7;
    wire mem_out_bus5_7;
    wire mem_out_bus1_7;
    wire dout_obuf_RNO_2Z0Z_7_cascade_;
    wire mem_N_150;
    wire mem_N_149_cascade_;
    wire dout_c_7;
    wire mem_out_bus2_1;
    wire mem_out_bus6_1;
    wire dout_obuf_RNO_5Z0Z_1;
    wire mem_out_bus6_0;
    wire mem_out_bus2_0;
    wire dout_obuf_RNO_5Z0Z_0;
    wire mem_out_bus6_3;
    wire mem_out_bus2_3;
    wire mem_out_bus7_0;
    wire mem_out_bus3_0;
    wire dout_obuf_RNO_3Z0Z_0;
    wire mem_out_bus7_2;
    wire mem_out_bus3_2;
    wire dout_obuf_RNO_3Z0Z_2;
    wire mem_out_bus7_3;
    wire mem_out_bus3_3;
    wire mem_out_bus4_2;
    wire mem_out_bus0_2;
    wire mem_out_bus4_3;
    wire mem_out_bus0_3;
    wire mem_out_bus4_5;
    wire mem_out_bus0_5;
    wire mem_out_bus0_4;
    wire mem_out_bus4_4;
    wire dout_obuf_RNO_4Z0Z_4;
    wire mem_N_180_cascade_;
    wire dout_c_4;
    wire dout_obuf_RNO_4Z0Z_6;
    wire mem_N_145_cascade_;
    wire dout_c_6;
    wire dout_obuf_RNO_4Z0Z_3;
    wire dout_obuf_RNO_5Z0Z_3;
    wire mem_out_bus5_3;
    wire mem_out_bus1_3;
    wire dout_obuf_RNO_3Z0Z_3;
    wire dout_obuf_RNO_2Z0Z_3_cascade_;
    wire mem_N_174;
    wire mem_N_172_cascade_;
    wire dout_c_3;
    wire dout_obuf_RNO_4Z0Z_2;
    wire mem_N_168;
    wire mem_out_bus1_4;
    wire mem_out_bus5_4;
    wire dout_obuf_RNO_2Z0Z_4_cascade_;
    wire mem_N_178;
    wire mem_out_bus1_6;
    wire mem_out_bus5_6;
    wire dout_obuf_RNO_2Z0Z_6_cascade_;
    wire mem_N_144;
    wire mem_out_bus6_4;
    wire mem_out_bus2_4;
    wire dout_obuf_RNO_5Z0Z_4;
    wire mem_out_bus2_2;
    wire mem_out_bus6_2;
    wire dout_obuf_RNO_5Z0Z_2;
    wire mem_out_bus6_6;
    wire mem_out_bus2_6;
    wire dout_obuf_RNO_5Z0Z_6;
    wire mem_out_bus6_7;
    wire mem_out_bus2_7;
    wire dout_obuf_RNO_5Z0Z_7;
    wire mem_out_bus7_1;
    wire mem_out_bus3_1;
    wire dout_obuf_RNO_3Z0Z_1;
    wire mem_out_bus7_4;
    wire mem_out_bus3_4;
    wire dout_obuf_RNO_3Z0Z_4;
    wire mem_out_bus7_7;
    wire mem_out_bus3_7;
    wire dout_obuf_RNO_3Z0Z_7;
    wire mem_out_bus7_6;
    wire mem_out_bus3_6;
    wire dout_obuf_RNO_3Z0Z_6;
    wire dout_obuf_RNO_4Z0Z_5;
    wire mem_out_bus1_5;
    wire mem_out_bus5_5;
    wire mem_radregZ0Z_12;
    wire dout_obuf_RNO_2Z0Z_5_cascade_;
    wire mem_N_140;
    wire mem_radregZ0Z_11;
    wire mem_N_139;
    wire dout_c_5;
    wire mem_out_bus6_5;
    wire mem_out_bus2_5;
    wire dout_obuf_RNO_5Z0Z_5;
    wire mem_radregZ0Z_13;
    wire mem_out_bus7_5;
    wire mem_out_bus3_5;
    wire dout_obuf_RNO_3Z0Z_5;
    wire _gnd_net_;

    defparam mem_mem_3_0_physical.WRITE_MODE=3;
    defparam mem_mem_3_0_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_3_0_physical (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,mem_out_bus3_1,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,mem_out_bus3_0,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__7339,N__6676,N__7774,N__8308,N__5356,N__9289,N__7114,N__4693,N__8533,N__5584,N__6244}),
            .WADDR({N__6028,N__6892,N__5806,N__6460,N__8857,N__8101,N__7558,N__9070,N__5140,N__4468,N__9685}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__8012,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__4991,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__4923),
            .RE(N__10964),
            .WCLKE(N__10238),
            .WCLK(N__8764),
            .WE(N__10985));
    defparam mem_mem_5_2_physical.WRITE_MODE=3;
    defparam mem_mem_5_2_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_5_2_physical (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,mem_out_bus5_5,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,mem_out_bus5_4,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__7390,N__6727,N__7831,N__8365,N__5419,N__9340,N__7177,N__4738,N__8590,N__5647,N__6295}),
            .WADDR({N__6073,N__6943,N__5857,N__6511,N__8896,N__8140,N__7609,N__9121,N__5185,N__4513,N__9742}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__9524,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__4368,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__4903),
            .RE(N__10636),
            .WCLKE(N__10317),
            .WCLK(N__8742),
            .WE(N__10632));
    defparam mem_mem_2_0_physical.WRITE_MODE=3;
    defparam mem_mem_2_0_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_2_0_physical (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,mem_out_bus2_1,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,mem_out_bus2_0,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__7387,N__6724,N__7822,N__8356,N__5404,N__9337,N__7162,N__4741,N__8581,N__5632,N__6292}),
            .WADDR({N__6076,N__6940,N__5854,N__6508,N__8905,N__8149,N__7606,N__9118,N__5188,N__4516,N__9733}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__8004,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__5018,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__4916),
            .RE(N__10899),
            .WCLKE(N__10196),
            .WCLK(N__8757),
            .WE(N__10924));
    defparam mem_mem_1_3_physical.WRITE_MODE=3;
    defparam mem_mem_1_3_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_1_3_physical (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,mem_out_bus1_7,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,mem_out_bus1_6,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__7399,N__6736,N__7834,N__8368,N__5416,N__9349,N__7174,N__4753,N__8593,N__5644,N__6304}),
            .WADDR({N__6088,N__6952,N__5866,N__6520,N__8917,N__8161,N__7618,N__9130,N__5200,N__4528,N__9745}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__4147,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__4247,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__4917),
            .RE(N__10898),
            .WCLKE(N__10136),
            .WCLK(N__8756),
            .WE(N__10878));
    defparam mem_mem_4_2_physical.WRITE_MODE=3;
    defparam mem_mem_4_2_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_4_2_physical (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,mem_out_bus4_5,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,mem_out_bus4_4,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__7438,N__6775,N__7879,N__8413,N__5467,N__9388,N__7225,N__4786,N__8638,N__5695,N__6343}),
            .WADDR({N__6121,N__6991,N__5905,N__6559,N__8944,N__8188,N__7657,N__9169,N__5233,N__4561,N__9790}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__9522,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__4376,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__4912),
            .RE(N__10594),
            .WCLKE(N__10281),
            .WCLK(N__8751),
            .WE(N__10703));
    defparam mem_mem_7_2_physical.WRITE_MODE=3;
    defparam mem_mem_7_2_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_7_2_physical (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,mem_out_bus7_5,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,mem_out_bus7_4,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__7294,N__6631,N__7735,N__8269,N__5323,N__9244,N__7081,N__4642,N__8494,N__5551,N__6199}),
            .WADDR({N__5977,N__6847,N__5761,N__6415,N__8800,N__8044,N__7513,N__9025,N__5089,N__4417,N__9646}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__9523,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__4324,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__4911),
            .RE(N__10869),
            .WCLKE(N__9565),
            .WCLK(N__8752),
            .WE(N__10921));
    defparam mem_mem_0_0_physical.WRITE_MODE=3;
    defparam mem_mem_0_0_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_0_0_physical (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,mem_out_bus0_1,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,mem_out_bus0_0,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__7472,N__6809,N__7910,N__8444,N__5495,N__9422,N__7253,N__4823,N__8669,N__5723,N__6377}),
            .WADDR({N__6158,N__7025,N__5939,N__6593,N__8984,N__8228,N__7691,N__9203,N__5270,N__4598,N__9821}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__8014,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__5051,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__4931),
            .RE(N__10960),
            .WCLKE(N__9938),
            .WCLK(N__8770),
            .WE(N__10931));
    defparam mem_mem_3_3_physical.WRITE_MODE=3;
    defparam mem_mem_3_3_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_3_3_physical (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,mem_out_bus3_7,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,mem_out_bus3_6,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__7303,N__6640,N__7738,N__8272,N__5320,N__9253,N__7078,N__4657,N__8497,N__5548,N__6208}),
            .WADDR({N__5992,N__6856,N__5770,N__6424,N__8821,N__8065,N__7522,N__9034,N__5104,N__4432,N__9649}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__4103,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__4190,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__4929),
            .RE(N__10998),
            .WCLKE(N__10247),
            .WCLK(N__8771),
            .WE(N__11000));
    defparam mem_mem_6_2_physical.WRITE_MODE=3;
    defparam mem_mem_6_2_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_6_2_physical (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,mem_out_bus6_5,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,mem_out_bus6_4,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__7342,N__6679,N__7783,N__8317,N__5371,N__9292,N__7129,N__4690,N__8542,N__5599,N__6247}),
            .WADDR({N__6025,N__6895,N__5809,N__6463,N__8848,N__8092,N__7561,N__9073,N__5137,N__4465,N__9694}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__9516,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__4349,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__4904),
            .RE(N__10710),
            .WCLKE(N__9598),
            .WCLK(N__8745),
            .WE(N__10787));
    defparam mem_mem_5_1_physical.WRITE_MODE=3;
    defparam mem_mem_5_1_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_5_1_physical (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,mem_out_bus5_3,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,mem_out_bus5_2,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__7402,N__6739,N__7843,N__8377,N__5431,N__9352,N__7189,N__4750,N__8602,N__5659,N__6307}),
            .WADDR({N__6085,N__6955,N__5869,N__6523,N__8908,N__8152,N__7621,N__9133,N__5197,N__4525,N__9754}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__4039,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__3925,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__4905),
            .RE(N__10582),
            .WCLKE(N__10324),
            .WCLK(N__8744),
            .WE(N__10589));
    defparam mem_mem_2_1_physical.WRITE_MODE=3;
    defparam mem_mem_2_1_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_2_1_physical (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,mem_out_bus2_3,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,mem_out_bus2_2,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__7375,N__6712,N__7810,N__8344,N__5392,N__9325,N__7150,N__4729,N__8569,N__5620,N__6280}),
            .WADDR({N__6064,N__6928,N__5842,N__6496,N__8893,N__8137,N__7594,N__9106,N__5176,N__4504,N__9721}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__4007,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__3881,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__4918),
            .RE(N__10932),
            .WCLKE(N__10197),
            .WCLK(N__8759),
            .WE(N__10925));
    defparam mem_mem_1_2_physical.WRITE_MODE=3;
    defparam mem_mem_1_2_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_1_2_physical (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,mem_out_bus1_5,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,mem_out_bus1_4,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__7411,N__6748,N__7846,N__8380,N__5428,N__9361,N__7186,N__4765,N__8605,N__5656,N__6316}),
            .WADDR({N__6100,N__6964,N__5878,N__6532,N__8929,N__8173,N__7630,N__9142,N__5212,N__4540,N__9757}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__9520,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__4355,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__4919),
            .RE(N__10842),
            .WCLKE(N__10137),
            .WCLK(N__8758),
            .WE(N__10877));
    defparam mem_mem_4_3_physical.WRITE_MODE=3;
    defparam mem_mem_4_3_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_4_3_physical (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,mem_out_bus4_7,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,mem_out_bus4_6,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__7426,N__6763,N__7867,N__8401,N__5455,N__9376,N__7213,N__4774,N__8626,N__5683,N__6331}),
            .WADDR({N__6109,N__6979,N__5893,N__6547,N__8932,N__8176,N__7645,N__9157,N__5221,N__4549,N__9778}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__4146,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__4262,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__4910),
            .RE(N__10637),
            .WCLKE(N__10272),
            .WCLK(N__8749),
            .WE(N__10590));
    defparam mem_mem_0_1_physical.WRITE_MODE=3;
    defparam mem_mem_0_1_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_0_1_physical (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,mem_out_bus0_3,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,mem_out_bus0_2,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__7466,N__6803,N__7904,N__8438,N__5488,N__9416,N__7246,N__4817,N__8663,N__5716,N__6371}),
            .WADDR({N__6152,N__7019,N__5933,N__6587,N__8978,N__8222,N__7685,N__9197,N__5264,N__4592,N__9815}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__4014,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__3891,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__4930),
            .RE(N__10926),
            .WCLKE(N__9937),
            .WCLK(N__8769),
            .WE(N__10927));
    defparam mem_mem_3_2_physical.WRITE_MODE=3;
    defparam mem_mem_3_2_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_3_2_physical (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,mem_out_bus3_5,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,mem_out_bus3_4,dangling_wire_627,dangling_wire_628,dangling_wire_629}),
            .RADDR({N__7315,N__6652,N__7750,N__8284,N__5332,N__9265,N__7090,N__4669,N__8509,N__5560,N__6220}),
            .WADDR({N__6004,N__6868,N__5782,N__6436,N__8833,N__8077,N__7534,N__9046,N__5116,N__4444,N__9661}),
            .MASK({dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645}),
            .WDATA({dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,N__9487,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,N__4303,dangling_wire_657,dangling_wire_658,dangling_wire_659}),
            .RCLKE(),
            .RCLK(N__4927),
            .RE(N__10991),
            .WCLKE(N__10246),
            .WCLK(N__8768),
            .WE(N__10999));
    defparam mem_mem_6_3_physical.WRITE_MODE=3;
    defparam mem_mem_6_3_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_6_3_physical (
            .RDATA({dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,mem_out_bus6_7,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,mem_out_bus6_6,dangling_wire_671,dangling_wire_672,dangling_wire_673}),
            .RADDR({N__7330,N__6667,N__7771,N__8305,N__5359,N__9280,N__7117,N__4678,N__8530,N__5587,N__6235}),
            .WADDR({N__6013,N__6883,N__5797,N__6451,N__8836,N__8080,N__7549,N__9061,N__5125,N__4453,N__9682}),
            .MASK({dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689}),
            .WDATA({dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,N__4131,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,N__4228,dangling_wire_701,dangling_wire_702,dangling_wire_703}),
            .RCLKE(),
            .RCLK(N__4906),
            .RE(N__10786),
            .WCLKE(N__9602),
            .WCLK(N__8747),
            .WE(N__10788));
    defparam mem_mem_5_0_physical.WRITE_MODE=3;
    defparam mem_mem_5_0_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_5_0_physical (
            .RDATA({dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,mem_out_bus5_1,dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,dangling_wire_714,mem_out_bus5_0,dangling_wire_715,dangling_wire_716,dangling_wire_717}),
            .RADDR({N__7414,N__6751,N__7855,N__8389,N__5443,N__9364,N__7201,N__4762,N__8614,N__5671,N__6319}),
            .WADDR({N__6097,N__6967,N__5881,N__6535,N__8920,N__8164,N__7633,N__9145,N__5209,N__4537,N__9766}),
            .MASK({dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,dangling_wire_723,dangling_wire_724,dangling_wire_725,dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733}),
            .WDATA({dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,N__8003,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,N__5036,dangling_wire_745,dangling_wire_746,dangling_wire_747}),
            .RCLKE(),
            .RCLK(N__4908),
            .RE(N__10530),
            .WCLKE(N__10325),
            .WCLK(N__8746),
            .WE(N__10631));
    defparam mem_mem_2_2_physical.WRITE_MODE=3;
    defparam mem_mem_2_2_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_2_2_physical (
            .RDATA({dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,mem_out_bus2_5,dangling_wire_752,dangling_wire_753,dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757,dangling_wire_758,mem_out_bus2_4,dangling_wire_759,dangling_wire_760,dangling_wire_761}),
            .RADDR({N__7363,N__6700,N__7798,N__8332,N__5380,N__9313,N__7138,N__4717,N__8557,N__5608,N__6268}),
            .WADDR({N__6052,N__6916,N__5830,N__6484,N__8881,N__8125,N__7582,N__9094,N__5164,N__4492,N__9709}),
            .MASK({dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,dangling_wire_767,dangling_wire_768,dangling_wire_769,dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777}),
            .WDATA({dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,N__9497,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785,dangling_wire_786,dangling_wire_787,dangling_wire_788,N__4330,dangling_wire_789,dangling_wire_790,dangling_wire_791}),
            .RCLKE(),
            .RCLK(N__4920),
            .RE(N__10933),
            .WCLKE(N__10198),
            .WCLK(N__8761),
            .WE(N__10961));
    defparam mem_mem_7_1_physical.WRITE_MODE=3;
    defparam mem_mem_7_1_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_7_1_physical (
            .RDATA({dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,mem_out_bus7_3,dangling_wire_796,dangling_wire_797,dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801,dangling_wire_802,mem_out_bus7_2,dangling_wire_803,dangling_wire_804,dangling_wire_805}),
            .RADDR({N__7306,N__6643,N__7747,N__8281,N__5335,N__9256,N__7093,N__4654,N__8506,N__5563,N__6211}),
            .WADDR({N__5989,N__6859,N__5773,N__6427,N__8812,N__8056,N__7525,N__9037,N__5101,N__4429,N__9658}),
            .MASK({dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,dangling_wire_811,dangling_wire_812,dangling_wire_813,dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821}),
            .WDATA({dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,N__4015,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829,dangling_wire_830,dangling_wire_831,dangling_wire_832,N__3906,dangling_wire_833,dangling_wire_834,dangling_wire_835}),
            .RCLKE(),
            .RCLK(N__4909),
            .RE(N__10868),
            .WCLKE(N__9558),
            .WCLK(N__8750),
            .WE(N__10864));
    defparam mem_mem_1_1_physical.WRITE_MODE=3;
    defparam mem_mem_1_1_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_1_1_physical (
            .RDATA({dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,mem_out_bus1_3,dangling_wire_840,dangling_wire_841,dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845,dangling_wire_846,mem_out_bus1_2,dangling_wire_847,dangling_wire_848,dangling_wire_849}),
            .RADDR({N__7423,N__6760,N__7858,N__8392,N__5440,N__9373,N__7198,N__4777,N__8617,N__5668,N__6328}),
            .WADDR({N__6112,N__6976,N__5890,N__6544,N__8941,N__8185,N__7642,N__9154,N__5224,N__4552,N__9769}),
            .MASK({dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,dangling_wire_855,dangling_wire_856,dangling_wire_857,dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865}),
            .WDATA({dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,N__3998,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873,dangling_wire_874,dangling_wire_875,dangling_wire_876,N__3890,dangling_wire_877,dangling_wire_878,dangling_wire_879}),
            .RCLKE(),
            .RCLK(N__4921),
            .RE(N__10828),
            .WCLKE(N__10144),
            .WCLK(N__8760),
            .WE(N__10816));
    defparam mem_mem_4_0_physical.WRITE_MODE=3;
    defparam mem_mem_4_0_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_4_0_physical (
            .RDATA({dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,mem_out_bus4_1,dangling_wire_884,dangling_wire_885,dangling_wire_886,dangling_wire_887,dangling_wire_888,dangling_wire_889,dangling_wire_890,mem_out_bus4_0,dangling_wire_891,dangling_wire_892,dangling_wire_893}),
            .RADDR({N__7462,N__6799,N__7903,N__8437,N__5491,N__9412,N__7249,N__4810,N__8662,N__5719,N__6367}),
            .WADDR({N__6145,N__7015,N__5929,N__6583,N__8968,N__8212,N__7681,N__9193,N__5257,N__4585,N__9814}),
            .MASK({dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,dangling_wire_899,dangling_wire_900,dangling_wire_901,dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909}),
            .WDATA({dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,N__8015,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917,dangling_wire_918,dangling_wire_919,dangling_wire_920,N__5050,dangling_wire_921,dangling_wire_922,dangling_wire_923}),
            .RCLKE(),
            .RCLK(N__4915),
            .RE(N__10811),
            .WCLKE(N__10289),
            .WCLK(N__8754),
            .WE(N__10740));
    defparam mem_mem_2_3_physical.WRITE_MODE=3;
    defparam mem_mem_2_3_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_2_3_physical (
            .RDATA({dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,mem_out_bus2_7,dangling_wire_928,dangling_wire_929,dangling_wire_930,dangling_wire_931,dangling_wire_932,dangling_wire_933,dangling_wire_934,mem_out_bus2_6,dangling_wire_935,dangling_wire_936,dangling_wire_937}),
            .RADDR({N__7351,N__6688,N__7786,N__8320,N__5368,N__9301,N__7126,N__4705,N__8545,N__5596,N__6256}),
            .WADDR({N__6040,N__6904,N__5818,N__6472,N__8869,N__8113,N__7570,N__9082,N__5152,N__4480,N__9697}),
            .MASK({dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,dangling_wire_943,dangling_wire_944,dangling_wire_945,dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953}),
            .WDATA({dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,N__4122,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961,dangling_wire_962,dangling_wire_963,dangling_wire_964,N__4219,dangling_wire_965,dangling_wire_966,dangling_wire_967}),
            .RCLKE(),
            .RCLK(N__4922),
            .RE(N__10963),
            .WCLKE(N__10202),
            .WCLK(N__8763),
            .WE(N__10962));
    defparam mem_mem_7_0_physical.WRITE_MODE=3;
    defparam mem_mem_7_0_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_7_0_physical (
            .RDATA({dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,mem_out_bus7_1,dangling_wire_972,dangling_wire_973,dangling_wire_974,dangling_wire_975,dangling_wire_976,dangling_wire_977,dangling_wire_978,mem_out_bus7_0,dangling_wire_979,dangling_wire_980,dangling_wire_981}),
            .RADDR({N__7318,N__6655,N__7759,N__8293,N__5347,N__9268,N__7105,N__4666,N__8518,N__5575,N__6223}),
            .WADDR({N__6001,N__6871,N__5785,N__6439,N__8824,N__8068,N__7537,N__9049,N__5113,N__4441,N__9670}),
            .MASK({dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,dangling_wire_987,dangling_wire_988,dangling_wire_989,dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997}),
            .WDATA({dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,N__8013,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005,dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,N__4984,dangling_wire_1009,dangling_wire_1010,dangling_wire_1011}),
            .RCLKE(),
            .RCLK(N__4907),
            .RE(N__10798),
            .WCLKE(N__9541),
            .WCLK(N__8748),
            .WE(N__10863));
    defparam mem_mem_1_0_physical.WRITE_MODE=3;
    defparam mem_mem_1_0_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_1_0_physical (
            .RDATA({dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,mem_out_bus1_1,dangling_wire_1016,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019,dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,mem_out_bus1_0,dangling_wire_1023,dangling_wire_1024,dangling_wire_1025}),
            .RADDR({N__7435,N__6772,N__7870,N__8404,N__5452,N__9385,N__7210,N__4789,N__8629,N__5680,N__6340}),
            .WADDR({N__6124,N__6988,N__5902,N__6556,N__8953,N__8197,N__7654,N__9166,N__5236,N__4564,N__9781}),
            .MASK({dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033,dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041}),
            .WDATA({dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,N__8002,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049,dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,N__5040,dangling_wire_1053,dangling_wire_1054,dangling_wire_1055}),
            .RCLKE(),
            .RCLK(N__4924),
            .RE(N__10876),
            .WCLKE(N__10145),
            .WCLK(N__8762),
            .WE(N__10812));
    defparam mem_mem_4_1_physical.WRITE_MODE=3;
    defparam mem_mem_4_1_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_4_1_physical (
            .RDATA({dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,mem_out_bus4_3,dangling_wire_1060,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063,dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,mem_out_bus4_2,dangling_wire_1067,dangling_wire_1068,dangling_wire_1069}),
            .RADDR({N__7450,N__6787,N__7891,N__8425,N__5479,N__9400,N__7237,N__4798,N__8650,N__5707,N__6355}),
            .WADDR({N__6133,N__7003,N__5917,N__6571,N__8956,N__8200,N__7669,N__9181,N__5245,N__4573,N__9802}),
            .MASK({dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077,dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085}),
            .WDATA({dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,N__4046,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093,dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,N__3932,dangling_wire_1097,dangling_wire_1098,dangling_wire_1099}),
            .RCLKE(),
            .RCLK(N__4914),
            .RE(N__10638),
            .WCLKE(N__10288),
            .WCLK(N__8753),
            .WE(N__10736));
    defparam mem_mem_0_2_physical.WRITE_MODE=3;
    defparam mem_mem_0_2_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_0_2_physical (
            .RDATA({dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,mem_out_bus0_5,dangling_wire_1104,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107,dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,mem_out_bus0_4,dangling_wire_1111,dangling_wire_1112,dangling_wire_1113}),
            .RADDR({N__7459,N__6796,N__7894,N__8428,N__5476,N__9409,N__7234,N__4811,N__8653,N__5704,N__6364}),
            .WADDR({N__6146,N__7012,N__5926,N__6580,N__8972,N__8216,N__7678,N__9190,N__5258,N__4586,N__9805}),
            .MASK({dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121,dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129}),
            .WDATA({dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,N__9521,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137,dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,N__4372,dangling_wire_1141,dangling_wire_1142,dangling_wire_1143}),
            .RCLKE(),
            .RCLK(N__4928),
            .RE(N__10920),
            .WCLKE(N__9936),
            .WCLK(N__8767),
            .WE(N__10862));
    defparam mem_mem_3_1_physical.WRITE_MODE=3;
    defparam mem_mem_3_1_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_3_1_physical (
            .RDATA({dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,mem_out_bus3_3,dangling_wire_1148,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151,dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,mem_out_bus3_2,dangling_wire_1155,dangling_wire_1156,dangling_wire_1157}),
            .RADDR({N__7327,N__6664,N__7762,N__8296,N__5344,N__9277,N__7102,N__4681,N__8521,N__5572,N__6232}),
            .WADDR({N__6016,N__6880,N__5794,N__6448,N__8845,N__8089,N__7546,N__9058,N__5128,N__4456,N__9673}),
            .MASK({dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165,dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173}),
            .WDATA({dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,N__3982,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181,dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,N__3868,dangling_wire_1185,dangling_wire_1186,dangling_wire_1187}),
            .RCLKE(),
            .RCLK(N__4925),
            .RE(N__10990),
            .WCLKE(N__10239),
            .WCLK(N__8766),
            .WE(N__10986));
    defparam mem_mem_6_0_physical.WRITE_MODE=3;
    defparam mem_mem_6_0_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_6_0_physical (
            .RDATA({dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,mem_out_bus6_1,dangling_wire_1192,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195,dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,mem_out_bus6_0,dangling_wire_1199,dangling_wire_1200,dangling_wire_1201}),
            .RADDR({N__7366,N__6703,N__7807,N__8341,N__5395,N__9316,N__7153,N__4714,N__8566,N__5623,N__6271}),
            .WADDR({N__6049,N__6919,N__5833,N__6487,N__8872,N__8116,N__7585,N__9097,N__5161,N__4489,N__9718}),
            .MASK({dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209,dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217}),
            .WDATA({dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,N__8005,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225,dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,N__5011,dangling_wire_1229,dangling_wire_1230,dangling_wire_1231}),
            .RCLKE(),
            .RCLK(N__4900),
            .RE(N__10641),
            .WCLKE(N__9587),
            .WCLK(N__8741),
            .WE(N__10704));
    defparam mem_mem_5_3_physical.WRITE_MODE=3;
    defparam mem_mem_5_3_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_5_3_physical (
            .RDATA({dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,mem_out_bus5_7,dangling_wire_1236,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239,dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,mem_out_bus5_6,dangling_wire_1243,dangling_wire_1244,dangling_wire_1245}),
            .RADDR({N__7378,N__6715,N__7819,N__8353,N__5407,N__9328,N__7165,N__4726,N__8578,N__5635,N__6283}),
            .WADDR({N__6061,N__6931,N__5845,N__6499,N__8884,N__8128,N__7597,N__9109,N__5173,N__4501,N__9730}),
            .MASK({dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253,dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261}),
            .WDATA({dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,N__4145,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269,dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,N__4251,dangling_wire_1273,dangling_wire_1274,dangling_wire_1275}),
            .RCLKE(),
            .RCLK(N__4901),
            .RE(N__10640),
            .WCLKE(N__10300),
            .WCLK(N__8740),
            .WE(N__10639));
    defparam mem_mem_7_3_physical.WRITE_MODE=3;
    defparam mem_mem_7_3_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_7_3_physical (
            .RDATA({dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,mem_out_bus7_7,dangling_wire_1280,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283,dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,mem_out_bus7_6,dangling_wire_1287,dangling_wire_1288,dangling_wire_1289}),
            .RADDR({N__7282,N__6619,N__7723,N__8257,N__5311,N__9232,N__7069,N__4630,N__8482,N__5539,N__6187}),
            .WADDR({N__5965,N__6835,N__5749,N__6403,N__8788,N__8032,N__7501,N__9013,N__5077,N__4405,N__9634}),
            .MASK({dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297,dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305}),
            .WDATA({dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,N__4144,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313,dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,N__4240,dangling_wire_1317,dangling_wire_1318,dangling_wire_1319}),
            .RCLKE(),
            .RCLK(N__4913),
            .RE(N__10922),
            .WCLKE(N__9566),
            .WCLK(N__8755),
            .WE(N__10923));
    defparam mem_mem_0_3_physical.WRITE_MODE=3;
    defparam mem_mem_0_3_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_0_3_physical (
            .RDATA({dangling_wire_1320,dangling_wire_1321,dangling_wire_1322,dangling_wire_1323,mem_out_bus0_7,dangling_wire_1324,dangling_wire_1325,dangling_wire_1326,dangling_wire_1327,dangling_wire_1328,dangling_wire_1329,dangling_wire_1330,mem_out_bus0_6,dangling_wire_1331,dangling_wire_1332,dangling_wire_1333}),
            .RADDR({N__7447,N__6784,N__7882,N__8416,N__5464,N__9397,N__7222,N__4801,N__8641,N__5692,N__6352}),
            .WADDR({N__6136,N__7000,N__5914,N__6568,N__8965,N__8209,N__7666,N__9178,N__5248,N__4576,N__9793}),
            .MASK({dangling_wire_1334,dangling_wire_1335,dangling_wire_1336,dangling_wire_1337,dangling_wire_1338,dangling_wire_1339,dangling_wire_1340,dangling_wire_1341,dangling_wire_1342,dangling_wire_1343,dangling_wire_1344,dangling_wire_1345,dangling_wire_1346,dangling_wire_1347,dangling_wire_1348,dangling_wire_1349}),
            .WDATA({dangling_wire_1350,dangling_wire_1351,dangling_wire_1352,dangling_wire_1353,N__4154,dangling_wire_1354,dangling_wire_1355,dangling_wire_1356,dangling_wire_1357,dangling_wire_1358,dangling_wire_1359,dangling_wire_1360,N__4261,dangling_wire_1361,dangling_wire_1362,dangling_wire_1363}),
            .RCLKE(),
            .RCLK(N__4926),
            .RE(N__10885),
            .WCLKE(N__9935),
            .WCLK(N__8765),
            .WE(N__10858));
    defparam mem_mem_6_1_physical.WRITE_MODE=3;
    defparam mem_mem_6_1_physical.READ_MODE=3;
    SB_RAM40_4K mem_mem_6_1_physical (
            .RDATA({dangling_wire_1364,dangling_wire_1365,dangling_wire_1366,dangling_wire_1367,mem_out_bus6_3,dangling_wire_1368,dangling_wire_1369,dangling_wire_1370,dangling_wire_1371,dangling_wire_1372,dangling_wire_1373,dangling_wire_1374,mem_out_bus6_2,dangling_wire_1375,dangling_wire_1376,dangling_wire_1377}),
            .RADDR({N__7354,N__6691,N__7795,N__8329,N__5383,N__9304,N__7141,N__4702,N__8554,N__5611,N__6259}),
            .WADDR({N__6037,N__6907,N__5821,N__6475,N__8860,N__8104,N__7573,N__9085,N__5149,N__4477,N__9706}),
            .MASK({dangling_wire_1378,dangling_wire_1379,dangling_wire_1380,dangling_wire_1381,dangling_wire_1382,dangling_wire_1383,dangling_wire_1384,dangling_wire_1385,dangling_wire_1386,dangling_wire_1387,dangling_wire_1388,dangling_wire_1389,dangling_wire_1390,dangling_wire_1391,dangling_wire_1392,dangling_wire_1393}),
            .WDATA({dangling_wire_1394,dangling_wire_1395,dangling_wire_1396,dangling_wire_1397,N__4027,dangling_wire_1398,dangling_wire_1399,dangling_wire_1400,dangling_wire_1401,dangling_wire_1402,dangling_wire_1403,dangling_wire_1404,N__3913,dangling_wire_1405,dangling_wire_1406,dangling_wire_1407}),
            .RCLKE(),
            .RCLK(N__4902),
            .RE(N__10709),
            .WCLKE(N__9597),
            .WCLK(N__8743),
            .WE(N__10705));
    PRE_IO_GBUF wclk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__13189),
            .GLOBALBUFFEROUTPUT(wclk_c_g));
    IO_PAD wclk_ibuf_gb_io_iopad (
            .OE(N__13191),
            .DIN(N__13190),
            .DOUT(N__13189),
            .PACKAGEPIN(wclk));
    defparam wclk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam wclk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO wclk_ibuf_gb_io_preio (
            .PADOEN(N__13191),
            .PADOUT(N__13190),
            .PADIN(N__13189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF rclk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__13179),
            .GLOBALBUFFEROUTPUT(rclk_c_g));
    IO_PAD rclk_ibuf_gb_io_iopad (
            .OE(N__13181),
            .DIN(N__13180),
            .DOUT(N__13179),
            .PACKAGEPIN(rclk));
    defparam rclk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam rclk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO rclk_ibuf_gb_io_preio (
            .PADOEN(N__13181),
            .PADOUT(N__13180),
            .PADIN(N__13179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_0_iopad (
            .OE(N__13170),
            .DIN(N__13169),
            .DOUT(N__13168),
            .PACKAGEPIN(waddr[0]));
    defparam waddr_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_0_preio (
            .PADOEN(N__13170),
            .PADOUT(N__13169),
            .PADIN(N__13168),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout_obuf_3_iopad (
            .OE(N__13161),
            .DIN(N__13160),
            .DOUT(N__13159),
            .PACKAGEPIN(dout[3]));
    defparam dout_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam dout_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO dout_obuf_3_preio (
            .PADOEN(N__13161),
            .PADOUT(N__13160),
            .PADIN(N__13159),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11819),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_12_iopad (
            .OE(N__13152),
            .DIN(N__13151),
            .DOUT(N__13150),
            .PACKAGEPIN(waddr[12]));
    defparam waddr_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_12_preio (
            .PADOEN(N__13152),
            .PADOUT(N__13151),
            .PADIN(N__13150),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_4_iopad (
            .OE(N__13143),
            .DIN(N__13142),
            .DOUT(N__13141),
            .PACKAGEPIN(waddr[4]));
    defparam waddr_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_4_preio (
            .PADOEN(N__13143),
            .PADOUT(N__13142),
            .PADIN(N__13141),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout_obuf_6_iopad (
            .OE(N__13134),
            .DIN(N__13133),
            .DOUT(N__13132),
            .PACKAGEPIN(dout[6]));
    defparam dout_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam dout_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO dout_obuf_6_preio (
            .PADOEN(N__13134),
            .PADOUT(N__13133),
            .PADIN(N__13132),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11522),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_3_iopad (
            .OE(N__13125),
            .DIN(N__13124),
            .DOUT(N__13123),
            .PACKAGEPIN(raddr[3]));
    defparam raddr_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_3_preio (
            .PADOEN(N__13125),
            .PADOUT(N__13124),
            .PADIN(N__13123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD din_ibuf_0_iopad (
            .OE(N__13116),
            .DIN(N__13115),
            .DOUT(N__13114),
            .PACKAGEPIN(din[0]));
    defparam din_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam din_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO din_ibuf_0_preio (
            .PADOEN(N__13116),
            .PADOUT(N__13115),
            .PADIN(N__13114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(din_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_3_iopad (
            .OE(N__13107),
            .DIN(N__13106),
            .DOUT(N__13105),
            .PACKAGEPIN(waddr[3]));
    defparam waddr_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_3_preio (
            .PADOEN(N__13107),
            .PADOUT(N__13106),
            .PADIN(N__13105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_11_iopad (
            .OE(N__13098),
            .DIN(N__13097),
            .DOUT(N__13096),
            .PACKAGEPIN(raddr[11]));
    defparam raddr_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_11_preio.PIN_TYPE=6'b000000;
    PRE_IO raddr_ibuf_11_preio (
            .PADOEN(N__13098),
            .PADOUT(N__13097),
            .PADIN(N__13096),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(mem_radregZ0Z_11),
            .DOUT0(),
            .INPUTCLK(N__4932),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_4_iopad (
            .OE(N__13089),
            .DIN(N__13088),
            .DOUT(N__13087),
            .PACKAGEPIN(raddr[4]));
    defparam raddr_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_4_preio (
            .PADOEN(N__13089),
            .PADOUT(N__13088),
            .PADIN(N__13087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_8_iopad (
            .OE(N__13080),
            .DIN(N__13079),
            .DOUT(N__13078),
            .PACKAGEPIN(waddr[8]));
    defparam waddr_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_8_preio (
            .PADOEN(N__13080),
            .PADOUT(N__13079),
            .PADIN(N__13078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout_obuf_2_iopad (
            .OE(N__13071),
            .DIN(N__13070),
            .DOUT(N__13069),
            .PACKAGEPIN(dout[2]));
    defparam dout_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam dout_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO dout_obuf_2_preio (
            .PADOEN(N__13071),
            .PADOUT(N__13070),
            .PADIN(N__13069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11102),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_13_iopad (
            .OE(N__13062),
            .DIN(N__13061),
            .DOUT(N__13060),
            .PACKAGEPIN(waddr[13]));
    defparam waddr_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_13_preio (
            .PADOEN(N__13062),
            .PADOUT(N__13061),
            .PADIN(N__13060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD din_ibuf_4_iopad (
            .OE(N__13053),
            .DIN(N__13052),
            .DOUT(N__13051),
            .PACKAGEPIN(din[4]));
    defparam din_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam din_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO din_ibuf_4_preio (
            .PADOEN(N__13053),
            .PADOUT(N__13052),
            .PADIN(N__13051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(din_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_7_iopad (
            .OE(N__13044),
            .DIN(N__13043),
            .DOUT(N__13042),
            .PACKAGEPIN(waddr[7]));
    defparam waddr_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_7_preio (
            .PADOEN(N__13044),
            .PADOUT(N__13043),
            .PADIN(N__13042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout_obuf_5_iopad (
            .OE(N__13035),
            .DIN(N__13034),
            .DOUT(N__13033),
            .PACKAGEPIN(dout[5]));
    defparam dout_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam dout_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO dout_obuf_5_preio (
            .PADOEN(N__13035),
            .PADOUT(N__13034),
            .PADIN(N__13033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12482),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_0_iopad (
            .OE(N__13026),
            .DIN(N__13025),
            .DOUT(N__13024),
            .PACKAGEPIN(raddr[0]));
    defparam raddr_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_0_preio (
            .PADOEN(N__13026),
            .PADOUT(N__13025),
            .PADIN(N__13024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD din_ibuf_1_iopad (
            .OE(N__13017),
            .DIN(N__13016),
            .DOUT(N__13015),
            .PACKAGEPIN(din[1]));
    defparam din_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam din_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO din_ibuf_1_preio (
            .PADOEN(N__13017),
            .PADOUT(N__13016),
            .PADIN(N__13015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(din_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_2_iopad (
            .OE(N__13008),
            .DIN(N__13007),
            .DOUT(N__13006),
            .PACKAGEPIN(waddr[2]));
    defparam waddr_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_2_preio (
            .PADOEN(N__13008),
            .PADOUT(N__13007),
            .PADIN(N__13006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_10_iopad (
            .OE(N__12999),
            .DIN(N__12998),
            .DOUT(N__12997),
            .PACKAGEPIN(raddr[10]));
    defparam raddr_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_10_preio (
            .PADOEN(N__12999),
            .PADOUT(N__12998),
            .PADIN(N__12997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_5_iopad (
            .OE(N__12990),
            .DIN(N__12989),
            .DOUT(N__12988),
            .PACKAGEPIN(raddr[5]));
    defparam raddr_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_5_preio (
            .PADOEN(N__12990),
            .PADOUT(N__12989),
            .PADIN(N__12988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout_obuf_1_iopad (
            .OE(N__12981),
            .DIN(N__12980),
            .DOUT(N__12979),
            .PACKAGEPIN(dout[1]));
    defparam dout_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam dout_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO dout_obuf_1_preio (
            .PADOEN(N__12981),
            .PADOUT(N__12980),
            .PADIN(N__12979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10370),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD din_ibuf_5_iopad (
            .OE(N__12972),
            .DIN(N__12971),
            .DOUT(N__12970),
            .PACKAGEPIN(din[5]));
    defparam din_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam din_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO din_ibuf_5_preio (
            .PADOEN(N__12972),
            .PADOUT(N__12971),
            .PADIN(N__12970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(din_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_6_iopad (
            .OE(N__12963),
            .DIN(N__12962),
            .DOUT(N__12961),
            .PACKAGEPIN(waddr[6]));
    defparam waddr_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_6_preio (
            .PADOEN(N__12963),
            .PADOUT(N__12962),
            .PADIN(N__12961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout_obuf_4_iopad (
            .OE(N__12954),
            .DIN(N__12953),
            .DOUT(N__12952),
            .PACKAGEPIN(dout[4]));
    defparam dout_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam dout_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO dout_obuf_4_preio (
            .PADOEN(N__12954),
            .PADOUT(N__12953),
            .PADIN(N__12952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11552),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_1_iopad (
            .OE(N__12945),
            .DIN(N__12944),
            .DOUT(N__12943),
            .PACKAGEPIN(raddr[1]));
    defparam raddr_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_1_preio (
            .PADOEN(N__12945),
            .PADOUT(N__12944),
            .PADIN(N__12943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_8_iopad (
            .OE(N__12936),
            .DIN(N__12935),
            .DOUT(N__12934),
            .PACKAGEPIN(raddr[8]));
    defparam raddr_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_8_preio (
            .PADOEN(N__12936),
            .PADOUT(N__12935),
            .PADIN(N__12934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_10_iopad (
            .OE(N__12927),
            .DIN(N__12926),
            .DOUT(N__12925),
            .PACKAGEPIN(waddr[10]));
    defparam waddr_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_10_preio (
            .PADOEN(N__12927),
            .PADOUT(N__12926),
            .PADIN(N__12925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD din_ibuf_2_iopad (
            .OE(N__12918),
            .DIN(N__12917),
            .DOUT(N__12916),
            .PACKAGEPIN(din[2]));
    defparam din_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam din_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO din_ibuf_2_preio (
            .PADOEN(N__12918),
            .PADOUT(N__12917),
            .PADIN(N__12916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(din_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_13_iopad (
            .OE(N__12909),
            .DIN(N__12908),
            .DOUT(N__12907),
            .PACKAGEPIN(raddr[13]));
    defparam raddr_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_13_preio.PIN_TYPE=6'b000000;
    PRE_IO raddr_ibuf_13_preio (
            .PADOEN(N__12909),
            .PADOUT(N__12908),
            .PADIN(N__12907),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(mem_radregZ0Z_13),
            .DOUT0(),
            .INPUTCLK(N__4934),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout_obuf_0_iopad (
            .OE(N__12900),
            .DIN(N__12899),
            .DOUT(N__12898),
            .PACKAGEPIN(dout[0]));
    defparam dout_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam dout_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO dout_obuf_0_preio (
            .PADOEN(N__12900),
            .PADOUT(N__12899),
            .PADIN(N__12898),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10343),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD din_ibuf_6_iopad (
            .OE(N__12891),
            .DIN(N__12890),
            .DOUT(N__12889),
            .PACKAGEPIN(din[6]));
    defparam din_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam din_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO din_ibuf_6_preio (
            .PADOEN(N__12891),
            .PADOUT(N__12890),
            .PADIN(N__12889),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(din_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_1_iopad (
            .OE(N__12882),
            .DIN(N__12881),
            .DOUT(N__12880),
            .PACKAGEPIN(waddr[1]));
    defparam waddr_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_1_preio (
            .PADOEN(N__12882),
            .PADOUT(N__12881),
            .PADIN(N__12880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_6_iopad (
            .OE(N__12873),
            .DIN(N__12872),
            .DOUT(N__12871),
            .PACKAGEPIN(raddr[6]));
    defparam raddr_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_6_preio (
            .PADOEN(N__12873),
            .PADOUT(N__12872),
            .PADIN(N__12871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_9_iopad (
            .OE(N__12864),
            .DIN(N__12863),
            .DOUT(N__12862),
            .PACKAGEPIN(raddr[9]));
    defparam raddr_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_9_preio (
            .PADOEN(N__12864),
            .PADOUT(N__12863),
            .PADIN(N__12862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_11_iopad (
            .OE(N__12855),
            .DIN(N__12854),
            .DOUT(N__12853),
            .PACKAGEPIN(waddr[11]));
    defparam waddr_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_11_preio (
            .PADOEN(N__12855),
            .PADOUT(N__12854),
            .PADIN(N__12853),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD din_ibuf_3_iopad (
            .OE(N__12846),
            .DIN(N__12845),
            .DOUT(N__12844),
            .PACKAGEPIN(din[3]));
    defparam din_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam din_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO din_ibuf_3_preio (
            .PADOEN(N__12846),
            .PADOUT(N__12845),
            .PADIN(N__12844),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(din_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_12_iopad (
            .OE(N__12837),
            .DIN(N__12836),
            .DOUT(N__12835),
            .PACKAGEPIN(raddr[12]));
    defparam raddr_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_12_preio.PIN_TYPE=6'b000000;
    PRE_IO raddr_ibuf_12_preio (
            .PADOEN(N__12837),
            .PADOUT(N__12836),
            .PADIN(N__12835),
            .CLOCKENABLE(VCCG0),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(mem_radregZ0Z_12),
            .DOUT0(),
            .INPUTCLK(N__4933),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_5_iopad (
            .OE(N__12828),
            .DIN(N__12827),
            .DOUT(N__12826),
            .PACKAGEPIN(waddr[5]));
    defparam waddr_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_5_preio (
            .PADOEN(N__12828),
            .PADOUT(N__12827),
            .PADIN(N__12826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD write_en_ibuf_iopad (
            .OE(N__12819),
            .DIN(N__12818),
            .DOUT(N__12817),
            .PACKAGEPIN(write_en));
    defparam write_en_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam write_en_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO write_en_ibuf_preio (
            .PADOEN(N__12819),
            .PADOUT(N__12818),
            .PADIN(N__12817),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(write_en_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout_obuf_7_iopad (
            .OE(N__12810),
            .DIN(N__12809),
            .DOUT(N__12808),
            .PACKAGEPIN(dout[7]));
    defparam dout_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam dout_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO dout_obuf_7_preio (
            .PADOEN(N__12810),
            .PADOUT(N__12809),
            .PADIN(N__12808),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11048),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_2_iopad (
            .OE(N__12801),
            .DIN(N__12800),
            .DOUT(N__12799),
            .PACKAGEPIN(raddr[2]));
    defparam raddr_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_2_preio (
            .PADOEN(N__12801),
            .PADOUT(N__12800),
            .PADIN(N__12799),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD din_ibuf_7_iopad (
            .OE(N__12792),
            .DIN(N__12791),
            .DOUT(N__12790),
            .PACKAGEPIN(din[7]));
    defparam din_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam din_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO din_ibuf_7_preio (
            .PADOEN(N__12792),
            .PADOUT(N__12791),
            .PADIN(N__12790),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(din_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD raddr_ibuf_7_iopad (
            .OE(N__12783),
            .DIN(N__12782),
            .DOUT(N__12781),
            .PACKAGEPIN(raddr[7]));
    defparam raddr_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam raddr_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO raddr_ibuf_7_preio (
            .PADOEN(N__12783),
            .PADOUT(N__12782),
            .PADIN(N__12781),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(raddr_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD waddr_ibuf_9_iopad (
            .OE(N__12774),
            .DIN(N__12773),
            .DOUT(N__12772),
            .PACKAGEPIN(waddr[9]));
    defparam waddr_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam waddr_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO waddr_ibuf_9_preio (
            .PADOEN(N__12774),
            .PADOUT(N__12773),
            .PADIN(N__12772),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(waddr_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3118 (
            .O(N__12755),
            .I(N__12752));
    LocalMux I__3117 (
            .O(N__12752),
            .I(N__12744));
    InMux I__3116 (
            .O(N__12751),
            .I(N__12739));
    InMux I__3115 (
            .O(N__12750),
            .I(N__12739));
    InMux I__3114 (
            .O(N__12749),
            .I(N__12736));
    InMux I__3113 (
            .O(N__12748),
            .I(N__12731));
    InMux I__3112 (
            .O(N__12747),
            .I(N__12731));
    Span4Mux_v I__3111 (
            .O(N__12744),
            .I(N__12719));
    LocalMux I__3110 (
            .O(N__12739),
            .I(N__12719));
    LocalMux I__3109 (
            .O(N__12736),
            .I(N__12719));
    LocalMux I__3108 (
            .O(N__12731),
            .I(N__12719));
    InMux I__3107 (
            .O(N__12730),
            .I(N__12716));
    InMux I__3106 (
            .O(N__12729),
            .I(N__12708));
    InMux I__3105 (
            .O(N__12728),
            .I(N__12705));
    Span4Mux_h I__3104 (
            .O(N__12719),
            .I(N__12700));
    LocalMux I__3103 (
            .O(N__12716),
            .I(N__12700));
    InMux I__3102 (
            .O(N__12715),
            .I(N__12697));
    InMux I__3101 (
            .O(N__12714),
            .I(N__12694));
    InMux I__3100 (
            .O(N__12713),
            .I(N__12691));
    InMux I__3099 (
            .O(N__12712),
            .I(N__12688));
    InMux I__3098 (
            .O(N__12711),
            .I(N__12685));
    LocalMux I__3097 (
            .O(N__12708),
            .I(N__12680));
    LocalMux I__3096 (
            .O(N__12705),
            .I(N__12677));
    Span4Mux_v I__3095 (
            .O(N__12700),
            .I(N__12674));
    LocalMux I__3094 (
            .O(N__12697),
            .I(N__12667));
    LocalMux I__3093 (
            .O(N__12694),
            .I(N__12667));
    LocalMux I__3092 (
            .O(N__12691),
            .I(N__12667));
    LocalMux I__3091 (
            .O(N__12688),
            .I(N__12662));
    LocalMux I__3090 (
            .O(N__12685),
            .I(N__12662));
    InMux I__3089 (
            .O(N__12684),
            .I(N__12659));
    InMux I__3088 (
            .O(N__12683),
            .I(N__12656));
    Span4Mux_v I__3087 (
            .O(N__12680),
            .I(N__12651));
    Span4Mux_v I__3086 (
            .O(N__12677),
            .I(N__12651));
    Span4Mux_h I__3085 (
            .O(N__12674),
            .I(N__12648));
    Span4Mux_h I__3084 (
            .O(N__12667),
            .I(N__12645));
    Span4Mux_h I__3083 (
            .O(N__12662),
            .I(N__12638));
    LocalMux I__3082 (
            .O(N__12659),
            .I(N__12638));
    LocalMux I__3081 (
            .O(N__12656),
            .I(N__12638));
    Span4Mux_h I__3080 (
            .O(N__12651),
            .I(N__12635));
    Span4Mux_h I__3079 (
            .O(N__12648),
            .I(N__12632));
    Span4Mux_h I__3078 (
            .O(N__12645),
            .I(N__12629));
    Span4Mux_h I__3077 (
            .O(N__12638),
            .I(N__12626));
    Sp12to4 I__3076 (
            .O(N__12635),
            .I(N__12623));
    Sp12to4 I__3075 (
            .O(N__12632),
            .I(N__12620));
    Sp12to4 I__3074 (
            .O(N__12629),
            .I(N__12615));
    Sp12to4 I__3073 (
            .O(N__12626),
            .I(N__12615));
    Span12Mux_h I__3072 (
            .O(N__12623),
            .I(N__12612));
    Span12Mux_h I__3071 (
            .O(N__12620),
            .I(N__12609));
    Span12Mux_v I__3070 (
            .O(N__12615),
            .I(N__12606));
    Span12Mux_v I__3069 (
            .O(N__12612),
            .I(N__12603));
    Span12Mux_v I__3068 (
            .O(N__12609),
            .I(N__12598));
    Span12Mux_h I__3067 (
            .O(N__12606),
            .I(N__12598));
    Odrv12 I__3066 (
            .O(N__12603),
            .I(mem_radregZ0Z_12));
    Odrv12 I__3065 (
            .O(N__12598),
            .I(mem_radregZ0Z_12));
    CascadeMux I__3064 (
            .O(N__12593),
            .I(dout_obuf_RNO_2Z0Z_5_cascade_));
    InMux I__3063 (
            .O(N__12590),
            .I(N__12587));
    LocalMux I__3062 (
            .O(N__12587),
            .I(mem_N_140));
    InMux I__3061 (
            .O(N__12584),
            .I(N__12581));
    LocalMux I__3060 (
            .O(N__12581),
            .I(N__12575));
    InMux I__3059 (
            .O(N__12580),
            .I(N__12572));
    InMux I__3058 (
            .O(N__12579),
            .I(N__12567));
    InMux I__3057 (
            .O(N__12578),
            .I(N__12567));
    Span4Mux_v I__3056 (
            .O(N__12575),
            .I(N__12561));
    LocalMux I__3055 (
            .O(N__12572),
            .I(N__12561));
    LocalMux I__3054 (
            .O(N__12567),
            .I(N__12555));
    InMux I__3053 (
            .O(N__12566),
            .I(N__12552));
    Span4Mux_v I__3052 (
            .O(N__12561),
            .I(N__12549));
    InMux I__3051 (
            .O(N__12560),
            .I(N__12546));
    InMux I__3050 (
            .O(N__12559),
            .I(N__12543));
    InMux I__3049 (
            .O(N__12558),
            .I(N__12540));
    Span4Mux_v I__3048 (
            .O(N__12555),
            .I(N__12535));
    LocalMux I__3047 (
            .O(N__12552),
            .I(N__12535));
    Span4Mux_h I__3046 (
            .O(N__12549),
            .I(N__12532));
    LocalMux I__3045 (
            .O(N__12546),
            .I(N__12529));
    LocalMux I__3044 (
            .O(N__12543),
            .I(N__12524));
    LocalMux I__3043 (
            .O(N__12540),
            .I(N__12524));
    Span4Mux_h I__3042 (
            .O(N__12535),
            .I(N__12521));
    Sp12to4 I__3041 (
            .O(N__12532),
            .I(N__12516));
    Span12Mux_h I__3040 (
            .O(N__12529),
            .I(N__12516));
    Span12Mux_h I__3039 (
            .O(N__12524),
            .I(N__12513));
    Sp12to4 I__3038 (
            .O(N__12521),
            .I(N__12510));
    Span12Mux_h I__3037 (
            .O(N__12516),
            .I(N__12507));
    Span12Mux_h I__3036 (
            .O(N__12513),
            .I(N__12504));
    Span12Mux_v I__3035 (
            .O(N__12510),
            .I(N__12501));
    Span12Mux_v I__3034 (
            .O(N__12507),
            .I(N__12498));
    Span12Mux_v I__3033 (
            .O(N__12504),
            .I(N__12493));
    Span12Mux_h I__3032 (
            .O(N__12501),
            .I(N__12493));
    Odrv12 I__3031 (
            .O(N__12498),
            .I(mem_radregZ0Z_11));
    Odrv12 I__3030 (
            .O(N__12493),
            .I(mem_radregZ0Z_11));
    InMux I__3029 (
            .O(N__12488),
            .I(N__12485));
    LocalMux I__3028 (
            .O(N__12485),
            .I(mem_N_139));
    IoInMux I__3027 (
            .O(N__12482),
            .I(N__12479));
    LocalMux I__3026 (
            .O(N__12479),
            .I(N__12476));
    IoSpan4Mux I__3025 (
            .O(N__12476),
            .I(N__12473));
    Span4Mux_s2_h I__3024 (
            .O(N__12473),
            .I(N__12470));
    Span4Mux_h I__3023 (
            .O(N__12470),
            .I(N__12467));
    Span4Mux_h I__3022 (
            .O(N__12467),
            .I(N__12464));
    Odrv4 I__3021 (
            .O(N__12464),
            .I(dout_c_5));
    InMux I__3020 (
            .O(N__12461),
            .I(N__12458));
    LocalMux I__3019 (
            .O(N__12458),
            .I(N__12455));
    Odrv12 I__3018 (
            .O(N__12455),
            .I(mem_out_bus6_5));
    InMux I__3017 (
            .O(N__12452),
            .I(N__12449));
    LocalMux I__3016 (
            .O(N__12449),
            .I(N__12446));
    Span12Mux_h I__3015 (
            .O(N__12446),
            .I(N__12443));
    Odrv12 I__3014 (
            .O(N__12443),
            .I(mem_out_bus2_5));
    InMux I__3013 (
            .O(N__12440),
            .I(N__12437));
    LocalMux I__3012 (
            .O(N__12437),
            .I(N__12434));
    Odrv12 I__3011 (
            .O(N__12434),
            .I(dout_obuf_RNO_5Z0Z_5));
    InMux I__3010 (
            .O(N__12431),
            .I(N__12425));
    InMux I__3009 (
            .O(N__12430),
            .I(N__12425));
    LocalMux I__3008 (
            .O(N__12425),
            .I(N__12420));
    InMux I__3007 (
            .O(N__12424),
            .I(N__12415));
    InMux I__3006 (
            .O(N__12423),
            .I(N__12415));
    Span4Mux_s2_v I__3005 (
            .O(N__12420),
            .I(N__12408));
    LocalMux I__3004 (
            .O(N__12415),
            .I(N__12408));
    InMux I__3003 (
            .O(N__12414),
            .I(N__12403));
    InMux I__3002 (
            .O(N__12413),
            .I(N__12403));
    Span4Mux_v I__3001 (
            .O(N__12408),
            .I(N__12394));
    LocalMux I__3000 (
            .O(N__12403),
            .I(N__12394));
    InMux I__2999 (
            .O(N__12402),
            .I(N__12391));
    CascadeMux I__2998 (
            .O(N__12401),
            .I(N__12388));
    CascadeMux I__2997 (
            .O(N__12400),
            .I(N__12385));
    InMux I__2996 (
            .O(N__12399),
            .I(N__12381));
    Span4Mux_v I__2995 (
            .O(N__12394),
            .I(N__12376));
    LocalMux I__2994 (
            .O(N__12391),
            .I(N__12376));
    InMux I__2993 (
            .O(N__12388),
            .I(N__12369));
    InMux I__2992 (
            .O(N__12385),
            .I(N__12369));
    InMux I__2991 (
            .O(N__12384),
            .I(N__12369));
    LocalMux I__2990 (
            .O(N__12381),
            .I(N__12366));
    Span4Mux_v I__2989 (
            .O(N__12376),
            .I(N__12359));
    LocalMux I__2988 (
            .O(N__12369),
            .I(N__12359));
    Span4Mux_v I__2987 (
            .O(N__12366),
            .I(N__12354));
    InMux I__2986 (
            .O(N__12365),
            .I(N__12351));
    CascadeMux I__2985 (
            .O(N__12364),
            .I(N__12346));
    Span4Mux_v I__2984 (
            .O(N__12359),
            .I(N__12342));
    InMux I__2983 (
            .O(N__12358),
            .I(N__12339));
    InMux I__2982 (
            .O(N__12357),
            .I(N__12336));
    Span4Mux_v I__2981 (
            .O(N__12354),
            .I(N__12330));
    LocalMux I__2980 (
            .O(N__12351),
            .I(N__12330));
    InMux I__2979 (
            .O(N__12350),
            .I(N__12322));
    InMux I__2978 (
            .O(N__12349),
            .I(N__12322));
    InMux I__2977 (
            .O(N__12346),
            .I(N__12315));
    InMux I__2976 (
            .O(N__12345),
            .I(N__12315));
    Span4Mux_v I__2975 (
            .O(N__12342),
            .I(N__12306));
    LocalMux I__2974 (
            .O(N__12339),
            .I(N__12306));
    LocalMux I__2973 (
            .O(N__12336),
            .I(N__12306));
    InMux I__2972 (
            .O(N__12335),
            .I(N__12303));
    Span4Mux_v I__2971 (
            .O(N__12330),
            .I(N__12300));
    InMux I__2970 (
            .O(N__12329),
            .I(N__12297));
    InMux I__2969 (
            .O(N__12328),
            .I(N__12294));
    InMux I__2968 (
            .O(N__12327),
            .I(N__12291));
    LocalMux I__2967 (
            .O(N__12322),
            .I(N__12286));
    InMux I__2966 (
            .O(N__12321),
            .I(N__12283));
    InMux I__2965 (
            .O(N__12320),
            .I(N__12280));
    LocalMux I__2964 (
            .O(N__12315),
            .I(N__12275));
    InMux I__2963 (
            .O(N__12314),
            .I(N__12270));
    InMux I__2962 (
            .O(N__12313),
            .I(N__12270));
    Span4Mux_v I__2961 (
            .O(N__12306),
            .I(N__12265));
    LocalMux I__2960 (
            .O(N__12303),
            .I(N__12265));
    Span4Mux_v I__2959 (
            .O(N__12300),
            .I(N__12258));
    LocalMux I__2958 (
            .O(N__12297),
            .I(N__12258));
    LocalMux I__2957 (
            .O(N__12294),
            .I(N__12253));
    LocalMux I__2956 (
            .O(N__12291),
            .I(N__12253));
    InMux I__2955 (
            .O(N__12290),
            .I(N__12248));
    InMux I__2954 (
            .O(N__12289),
            .I(N__12248));
    Span12Mux_h I__2953 (
            .O(N__12286),
            .I(N__12245));
    LocalMux I__2952 (
            .O(N__12283),
            .I(N__12240));
    LocalMux I__2951 (
            .O(N__12280),
            .I(N__12240));
    InMux I__2950 (
            .O(N__12279),
            .I(N__12235));
    InMux I__2949 (
            .O(N__12278),
            .I(N__12235));
    Span12Mux_h I__2948 (
            .O(N__12275),
            .I(N__12232));
    LocalMux I__2947 (
            .O(N__12270),
            .I(N__12229));
    Span4Mux_v I__2946 (
            .O(N__12265),
            .I(N__12226));
    InMux I__2945 (
            .O(N__12264),
            .I(N__12221));
    InMux I__2944 (
            .O(N__12263),
            .I(N__12221));
    Span4Mux_v I__2943 (
            .O(N__12258),
            .I(N__12218));
    Span12Mux_h I__2942 (
            .O(N__12253),
            .I(N__12215));
    LocalMux I__2941 (
            .O(N__12248),
            .I(N__12212));
    Span12Mux_h I__2940 (
            .O(N__12245),
            .I(N__12209));
    Span12Mux_h I__2939 (
            .O(N__12240),
            .I(N__12206));
    LocalMux I__2938 (
            .O(N__12235),
            .I(N__12203));
    Span12Mux_h I__2937 (
            .O(N__12232),
            .I(N__12200));
    Span12Mux_h I__2936 (
            .O(N__12229),
            .I(N__12197));
    Sp12to4 I__2935 (
            .O(N__12226),
            .I(N__12192));
    LocalMux I__2934 (
            .O(N__12221),
            .I(N__12192));
    Span4Mux_h I__2933 (
            .O(N__12218),
            .I(N__12189));
    Span12Mux_h I__2932 (
            .O(N__12215),
            .I(N__12186));
    Span12Mux_h I__2931 (
            .O(N__12212),
            .I(N__12183));
    Span12Mux_v I__2930 (
            .O(N__12209),
            .I(N__12178));
    Span12Mux_h I__2929 (
            .O(N__12206),
            .I(N__12178));
    Span12Mux_h I__2928 (
            .O(N__12203),
            .I(N__12175));
    Span12Mux_v I__2927 (
            .O(N__12200),
            .I(N__12170));
    Span12Mux_h I__2926 (
            .O(N__12197),
            .I(N__12170));
    Span12Mux_h I__2925 (
            .O(N__12192),
            .I(N__12165));
    Sp12to4 I__2924 (
            .O(N__12189),
            .I(N__12165));
    Span12Mux_v I__2923 (
            .O(N__12186),
            .I(N__12160));
    Span12Mux_h I__2922 (
            .O(N__12183),
            .I(N__12160));
    Span12Mux_v I__2921 (
            .O(N__12178),
            .I(N__12155));
    Span12Mux_h I__2920 (
            .O(N__12175),
            .I(N__12155));
    Span12Mux_v I__2919 (
            .O(N__12170),
            .I(N__12150));
    Span12Mux_h I__2918 (
            .O(N__12165),
            .I(N__12150));
    Odrv12 I__2917 (
            .O(N__12160),
            .I(mem_radregZ0Z_13));
    Odrv12 I__2916 (
            .O(N__12155),
            .I(mem_radregZ0Z_13));
    Odrv12 I__2915 (
            .O(N__12150),
            .I(mem_radregZ0Z_13));
    InMux I__2914 (
            .O(N__12143),
            .I(N__12140));
    LocalMux I__2913 (
            .O(N__12140),
            .I(N__12137));
    Odrv12 I__2912 (
            .O(N__12137),
            .I(mem_out_bus7_5));
    InMux I__2911 (
            .O(N__12134),
            .I(N__12131));
    LocalMux I__2910 (
            .O(N__12131),
            .I(N__12128));
    Span12Mux_h I__2909 (
            .O(N__12128),
            .I(N__12125));
    Odrv12 I__2908 (
            .O(N__12125),
            .I(mem_out_bus3_5));
    InMux I__2907 (
            .O(N__12122),
            .I(N__12119));
    LocalMux I__2906 (
            .O(N__12119),
            .I(N__12116));
    Span12Mux_v I__2905 (
            .O(N__12116),
            .I(N__12113));
    Odrv12 I__2904 (
            .O(N__12113),
            .I(dout_obuf_RNO_3Z0Z_5));
    InMux I__2903 (
            .O(N__12110),
            .I(N__12107));
    LocalMux I__2902 (
            .O(N__12107),
            .I(N__12104));
    Span4Mux_v I__2901 (
            .O(N__12104),
            .I(N__12101));
    Odrv4 I__2900 (
            .O(N__12101),
            .I(mem_out_bus6_6));
    InMux I__2899 (
            .O(N__12098),
            .I(N__12095));
    LocalMux I__2898 (
            .O(N__12095),
            .I(N__12092));
    Span4Mux_v I__2897 (
            .O(N__12092),
            .I(N__12089));
    Sp12to4 I__2896 (
            .O(N__12089),
            .I(N__12086));
    Span12Mux_h I__2895 (
            .O(N__12086),
            .I(N__12083));
    Odrv12 I__2894 (
            .O(N__12083),
            .I(mem_out_bus2_6));
    InMux I__2893 (
            .O(N__12080),
            .I(N__12077));
    LocalMux I__2892 (
            .O(N__12077),
            .I(N__12074));
    Span12Mux_v I__2891 (
            .O(N__12074),
            .I(N__12071));
    Odrv12 I__2890 (
            .O(N__12071),
            .I(dout_obuf_RNO_5Z0Z_6));
    InMux I__2889 (
            .O(N__12068),
            .I(N__12065));
    LocalMux I__2888 (
            .O(N__12065),
            .I(N__12062));
    Odrv12 I__2887 (
            .O(N__12062),
            .I(mem_out_bus6_7));
    InMux I__2886 (
            .O(N__12059),
            .I(N__12056));
    LocalMux I__2885 (
            .O(N__12056),
            .I(N__12053));
    Span12Mux_h I__2884 (
            .O(N__12053),
            .I(N__12050));
    Odrv12 I__2883 (
            .O(N__12050),
            .I(mem_out_bus2_7));
    InMux I__2882 (
            .O(N__12047),
            .I(N__12044));
    LocalMux I__2881 (
            .O(N__12044),
            .I(N__12041));
    Span4Mux_v I__2880 (
            .O(N__12041),
            .I(N__12038));
    Span4Mux_v I__2879 (
            .O(N__12038),
            .I(N__12035));
    Odrv4 I__2878 (
            .O(N__12035),
            .I(dout_obuf_RNO_5Z0Z_7));
    InMux I__2877 (
            .O(N__12032),
            .I(N__12029));
    LocalMux I__2876 (
            .O(N__12029),
            .I(N__12026));
    Odrv4 I__2875 (
            .O(N__12026),
            .I(mem_out_bus7_1));
    InMux I__2874 (
            .O(N__12023),
            .I(N__12020));
    LocalMux I__2873 (
            .O(N__12020),
            .I(N__12017));
    Span12Mux_h I__2872 (
            .O(N__12017),
            .I(N__12014));
    Odrv12 I__2871 (
            .O(N__12014),
            .I(mem_out_bus3_1));
    InMux I__2870 (
            .O(N__12011),
            .I(N__12008));
    LocalMux I__2869 (
            .O(N__12008),
            .I(N__12005));
    Sp12to4 I__2868 (
            .O(N__12005),
            .I(N__12002));
    Span12Mux_v I__2867 (
            .O(N__12002),
            .I(N__11999));
    Odrv12 I__2866 (
            .O(N__11999),
            .I(dout_obuf_RNO_3Z0Z_1));
    InMux I__2865 (
            .O(N__11996),
            .I(N__11993));
    LocalMux I__2864 (
            .O(N__11993),
            .I(N__11990));
    Span4Mux_v I__2863 (
            .O(N__11990),
            .I(N__11987));
    Odrv4 I__2862 (
            .O(N__11987),
            .I(mem_out_bus7_4));
    InMux I__2861 (
            .O(N__11984),
            .I(N__11981));
    LocalMux I__2860 (
            .O(N__11981),
            .I(N__11978));
    Span4Mux_v I__2859 (
            .O(N__11978),
            .I(N__11975));
    Sp12to4 I__2858 (
            .O(N__11975),
            .I(N__11972));
    Span12Mux_h I__2857 (
            .O(N__11972),
            .I(N__11969));
    Odrv12 I__2856 (
            .O(N__11969),
            .I(mem_out_bus3_4));
    InMux I__2855 (
            .O(N__11966),
            .I(N__11963));
    LocalMux I__2854 (
            .O(N__11963),
            .I(N__11960));
    Span4Mux_v I__2853 (
            .O(N__11960),
            .I(N__11957));
    Span4Mux_v I__2852 (
            .O(N__11957),
            .I(N__11954));
    Span4Mux_v I__2851 (
            .O(N__11954),
            .I(N__11951));
    Span4Mux_v I__2850 (
            .O(N__11951),
            .I(N__11948));
    Odrv4 I__2849 (
            .O(N__11948),
            .I(dout_obuf_RNO_3Z0Z_4));
    InMux I__2848 (
            .O(N__11945),
            .I(N__11942));
    LocalMux I__2847 (
            .O(N__11942),
            .I(N__11939));
    Odrv4 I__2846 (
            .O(N__11939),
            .I(mem_out_bus7_7));
    InMux I__2845 (
            .O(N__11936),
            .I(N__11933));
    LocalMux I__2844 (
            .O(N__11933),
            .I(N__11930));
    Span12Mux_h I__2843 (
            .O(N__11930),
            .I(N__11927));
    Odrv12 I__2842 (
            .O(N__11927),
            .I(mem_out_bus3_7));
    InMux I__2841 (
            .O(N__11924),
            .I(N__11921));
    LocalMux I__2840 (
            .O(N__11921),
            .I(N__11918));
    Sp12to4 I__2839 (
            .O(N__11918),
            .I(N__11915));
    Span12Mux_v I__2838 (
            .O(N__11915),
            .I(N__11912));
    Odrv12 I__2837 (
            .O(N__11912),
            .I(dout_obuf_RNO_3Z0Z_7));
    InMux I__2836 (
            .O(N__11909),
            .I(N__11906));
    LocalMux I__2835 (
            .O(N__11906),
            .I(N__11903));
    Span4Mux_h I__2834 (
            .O(N__11903),
            .I(N__11900));
    Odrv4 I__2833 (
            .O(N__11900),
            .I(mem_out_bus7_6));
    InMux I__2832 (
            .O(N__11897),
            .I(N__11894));
    LocalMux I__2831 (
            .O(N__11894),
            .I(N__11891));
    Span4Mux_v I__2830 (
            .O(N__11891),
            .I(N__11888));
    Sp12to4 I__2829 (
            .O(N__11888),
            .I(N__11885));
    Span12Mux_h I__2828 (
            .O(N__11885),
            .I(N__11882));
    Odrv12 I__2827 (
            .O(N__11882),
            .I(mem_out_bus3_6));
    InMux I__2826 (
            .O(N__11879),
            .I(N__11876));
    LocalMux I__2825 (
            .O(N__11876),
            .I(N__11873));
    Sp12to4 I__2824 (
            .O(N__11873),
            .I(N__11870));
    Span12Mux_v I__2823 (
            .O(N__11870),
            .I(N__11867));
    Span12Mux_v I__2822 (
            .O(N__11867),
            .I(N__11864));
    Odrv12 I__2821 (
            .O(N__11864),
            .I(dout_obuf_RNO_3Z0Z_6));
    InMux I__2820 (
            .O(N__11861),
            .I(N__11858));
    LocalMux I__2819 (
            .O(N__11858),
            .I(N__11855));
    Span12Mux_h I__2818 (
            .O(N__11855),
            .I(N__11852));
    Odrv12 I__2817 (
            .O(N__11852),
            .I(dout_obuf_RNO_4Z0Z_5));
    InMux I__2816 (
            .O(N__11849),
            .I(N__11846));
    LocalMux I__2815 (
            .O(N__11846),
            .I(N__11843));
    Span12Mux_h I__2814 (
            .O(N__11843),
            .I(N__11840));
    Odrv12 I__2813 (
            .O(N__11840),
            .I(mem_out_bus1_5));
    InMux I__2812 (
            .O(N__11837),
            .I(N__11834));
    LocalMux I__2811 (
            .O(N__11834),
            .I(N__11831));
    Odrv12 I__2810 (
            .O(N__11831),
            .I(mem_out_bus5_5));
    InMux I__2809 (
            .O(N__11828),
            .I(N__11825));
    LocalMux I__2808 (
            .O(N__11825),
            .I(mem_N_174));
    CascadeMux I__2807 (
            .O(N__11822),
            .I(mem_N_172_cascade_));
    IoInMux I__2806 (
            .O(N__11819),
            .I(N__11816));
    LocalMux I__2805 (
            .O(N__11816),
            .I(N__11813));
    Span12Mux_s8_h I__2804 (
            .O(N__11813),
            .I(N__11810));
    Odrv12 I__2803 (
            .O(N__11810),
            .I(dout_c_3));
    InMux I__2802 (
            .O(N__11807),
            .I(N__11804));
    LocalMux I__2801 (
            .O(N__11804),
            .I(N__11801));
    Span12Mux_v I__2800 (
            .O(N__11801),
            .I(N__11798));
    Odrv12 I__2799 (
            .O(N__11798),
            .I(dout_obuf_RNO_4Z0Z_2));
    InMux I__2798 (
            .O(N__11795),
            .I(N__11792));
    LocalMux I__2797 (
            .O(N__11792),
            .I(mem_N_168));
    InMux I__2796 (
            .O(N__11789),
            .I(N__11786));
    LocalMux I__2795 (
            .O(N__11786),
            .I(N__11783));
    Span4Mux_v I__2794 (
            .O(N__11783),
            .I(N__11780));
    Sp12to4 I__2793 (
            .O(N__11780),
            .I(N__11777));
    Span12Mux_h I__2792 (
            .O(N__11777),
            .I(N__11774));
    Odrv12 I__2791 (
            .O(N__11774),
            .I(mem_out_bus1_4));
    InMux I__2790 (
            .O(N__11771),
            .I(N__11768));
    LocalMux I__2789 (
            .O(N__11768),
            .I(N__11765));
    Span4Mux_v I__2788 (
            .O(N__11765),
            .I(N__11762));
    Odrv4 I__2787 (
            .O(N__11762),
            .I(mem_out_bus5_4));
    CascadeMux I__2786 (
            .O(N__11759),
            .I(dout_obuf_RNO_2Z0Z_4_cascade_));
    InMux I__2785 (
            .O(N__11756),
            .I(N__11753));
    LocalMux I__2784 (
            .O(N__11753),
            .I(N__11750));
    Span4Mux_v I__2783 (
            .O(N__11750),
            .I(N__11747));
    Odrv4 I__2782 (
            .O(N__11747),
            .I(mem_N_178));
    InMux I__2781 (
            .O(N__11744),
            .I(N__11741));
    LocalMux I__2780 (
            .O(N__11741),
            .I(N__11738));
    Span4Mux_v I__2779 (
            .O(N__11738),
            .I(N__11735));
    Sp12to4 I__2778 (
            .O(N__11735),
            .I(N__11732));
    Span12Mux_h I__2777 (
            .O(N__11732),
            .I(N__11729));
    Odrv12 I__2776 (
            .O(N__11729),
            .I(mem_out_bus1_6));
    InMux I__2775 (
            .O(N__11726),
            .I(N__11723));
    LocalMux I__2774 (
            .O(N__11723),
            .I(N__11720));
    Span4Mux_v I__2773 (
            .O(N__11720),
            .I(N__11717));
    Odrv4 I__2772 (
            .O(N__11717),
            .I(mem_out_bus5_6));
    CascadeMux I__2771 (
            .O(N__11714),
            .I(dout_obuf_RNO_2Z0Z_6_cascade_));
    InMux I__2770 (
            .O(N__11711),
            .I(N__11708));
    LocalMux I__2769 (
            .O(N__11708),
            .I(N__11705));
    Span4Mux_v I__2768 (
            .O(N__11705),
            .I(N__11702));
    Odrv4 I__2767 (
            .O(N__11702),
            .I(mem_N_144));
    InMux I__2766 (
            .O(N__11699),
            .I(N__11696));
    LocalMux I__2765 (
            .O(N__11696),
            .I(N__11693));
    Span4Mux_v I__2764 (
            .O(N__11693),
            .I(N__11690));
    Odrv4 I__2763 (
            .O(N__11690),
            .I(mem_out_bus6_4));
    InMux I__2762 (
            .O(N__11687),
            .I(N__11684));
    LocalMux I__2761 (
            .O(N__11684),
            .I(N__11681));
    Span4Mux_v I__2760 (
            .O(N__11681),
            .I(N__11678));
    Sp12to4 I__2759 (
            .O(N__11678),
            .I(N__11675));
    Span12Mux_h I__2758 (
            .O(N__11675),
            .I(N__11672));
    Odrv12 I__2757 (
            .O(N__11672),
            .I(mem_out_bus2_4));
    InMux I__2756 (
            .O(N__11669),
            .I(N__11666));
    LocalMux I__2755 (
            .O(N__11666),
            .I(N__11663));
    Span12Mux_v I__2754 (
            .O(N__11663),
            .I(N__11660));
    Odrv12 I__2753 (
            .O(N__11660),
            .I(dout_obuf_RNO_5Z0Z_4));
    InMux I__2752 (
            .O(N__11657),
            .I(N__11654));
    LocalMux I__2751 (
            .O(N__11654),
            .I(N__11651));
    Span4Mux_v I__2750 (
            .O(N__11651),
            .I(N__11648));
    Sp12to4 I__2749 (
            .O(N__11648),
            .I(N__11645));
    Span12Mux_h I__2748 (
            .O(N__11645),
            .I(N__11642));
    Odrv12 I__2747 (
            .O(N__11642),
            .I(mem_out_bus2_2));
    InMux I__2746 (
            .O(N__11639),
            .I(N__11636));
    LocalMux I__2745 (
            .O(N__11636),
            .I(N__11633));
    Span4Mux_v I__2744 (
            .O(N__11633),
            .I(N__11630));
    Odrv4 I__2743 (
            .O(N__11630),
            .I(mem_out_bus6_2));
    InMux I__2742 (
            .O(N__11627),
            .I(N__11624));
    LocalMux I__2741 (
            .O(N__11624),
            .I(N__11621));
    Odrv12 I__2740 (
            .O(N__11621),
            .I(dout_obuf_RNO_5Z0Z_2));
    InMux I__2739 (
            .O(N__11618),
            .I(N__11615));
    LocalMux I__2738 (
            .O(N__11615),
            .I(N__11612));
    Odrv4 I__2737 (
            .O(N__11612),
            .I(mem_out_bus4_5));
    InMux I__2736 (
            .O(N__11609),
            .I(N__11606));
    LocalMux I__2735 (
            .O(N__11606),
            .I(N__11603));
    Span12Mux_h I__2734 (
            .O(N__11603),
            .I(N__11600));
    Odrv12 I__2733 (
            .O(N__11600),
            .I(mem_out_bus0_5));
    InMux I__2732 (
            .O(N__11597),
            .I(N__11594));
    LocalMux I__2731 (
            .O(N__11594),
            .I(N__11591));
    Span4Mux_v I__2730 (
            .O(N__11591),
            .I(N__11588));
    Sp12to4 I__2729 (
            .O(N__11588),
            .I(N__11585));
    Span12Mux_h I__2728 (
            .O(N__11585),
            .I(N__11582));
    Odrv12 I__2727 (
            .O(N__11582),
            .I(mem_out_bus0_4));
    InMux I__2726 (
            .O(N__11579),
            .I(N__11576));
    LocalMux I__2725 (
            .O(N__11576),
            .I(N__11573));
    Span4Mux_v I__2724 (
            .O(N__11573),
            .I(N__11570));
    Odrv4 I__2723 (
            .O(N__11570),
            .I(mem_out_bus4_4));
    InMux I__2722 (
            .O(N__11567),
            .I(N__11564));
    LocalMux I__2721 (
            .O(N__11564),
            .I(N__11561));
    Span4Mux_v I__2720 (
            .O(N__11561),
            .I(N__11558));
    Odrv4 I__2719 (
            .O(N__11558),
            .I(dout_obuf_RNO_4Z0Z_4));
    CascadeMux I__2718 (
            .O(N__11555),
            .I(mem_N_180_cascade_));
    IoInMux I__2717 (
            .O(N__11552),
            .I(N__11549));
    LocalMux I__2716 (
            .O(N__11549),
            .I(N__11546));
    Span4Mux_s2_h I__2715 (
            .O(N__11546),
            .I(N__11543));
    Span4Mux_h I__2714 (
            .O(N__11543),
            .I(N__11540));
    Span4Mux_h I__2713 (
            .O(N__11540),
            .I(N__11537));
    Odrv4 I__2712 (
            .O(N__11537),
            .I(dout_c_4));
    InMux I__2711 (
            .O(N__11534),
            .I(N__11531));
    LocalMux I__2710 (
            .O(N__11531),
            .I(N__11528));
    Odrv4 I__2709 (
            .O(N__11528),
            .I(dout_obuf_RNO_4Z0Z_6));
    CascadeMux I__2708 (
            .O(N__11525),
            .I(mem_N_145_cascade_));
    IoInMux I__2707 (
            .O(N__11522),
            .I(N__11519));
    LocalMux I__2706 (
            .O(N__11519),
            .I(N__11516));
    Span4Mux_s2_h I__2705 (
            .O(N__11516),
            .I(N__11513));
    Span4Mux_h I__2704 (
            .O(N__11513),
            .I(N__11510));
    Span4Mux_h I__2703 (
            .O(N__11510),
            .I(N__11507));
    Odrv4 I__2702 (
            .O(N__11507),
            .I(dout_c_6));
    InMux I__2701 (
            .O(N__11504),
            .I(N__11501));
    LocalMux I__2700 (
            .O(N__11501),
            .I(N__11498));
    Sp12to4 I__2699 (
            .O(N__11498),
            .I(N__11495));
    Odrv12 I__2698 (
            .O(N__11495),
            .I(dout_obuf_RNO_4Z0Z_3));
    InMux I__2697 (
            .O(N__11492),
            .I(N__11489));
    LocalMux I__2696 (
            .O(N__11489),
            .I(N__11486));
    Span4Mux_v I__2695 (
            .O(N__11486),
            .I(N__11483));
    Odrv4 I__2694 (
            .O(N__11483),
            .I(dout_obuf_RNO_5Z0Z_3));
    InMux I__2693 (
            .O(N__11480),
            .I(N__11477));
    LocalMux I__2692 (
            .O(N__11477),
            .I(N__11474));
    Odrv4 I__2691 (
            .O(N__11474),
            .I(mem_out_bus5_3));
    InMux I__2690 (
            .O(N__11471),
            .I(N__11468));
    LocalMux I__2689 (
            .O(N__11468),
            .I(N__11465));
    Span12Mux_h I__2688 (
            .O(N__11465),
            .I(N__11462));
    Span12Mux_h I__2687 (
            .O(N__11462),
            .I(N__11459));
    Odrv12 I__2686 (
            .O(N__11459),
            .I(mem_out_bus1_3));
    InMux I__2685 (
            .O(N__11456),
            .I(N__11453));
    LocalMux I__2684 (
            .O(N__11453),
            .I(N__11450));
    Span12Mux_v I__2683 (
            .O(N__11450),
            .I(N__11447));
    Span12Mux_v I__2682 (
            .O(N__11447),
            .I(N__11444));
    Odrv12 I__2681 (
            .O(N__11444),
            .I(dout_obuf_RNO_3Z0Z_3));
    CascadeMux I__2680 (
            .O(N__11441),
            .I(dout_obuf_RNO_2Z0Z_3_cascade_));
    InMux I__2679 (
            .O(N__11438),
            .I(N__11435));
    LocalMux I__2678 (
            .O(N__11435),
            .I(N__11432));
    Span12Mux_h I__2677 (
            .O(N__11432),
            .I(N__11429));
    Span12Mux_h I__2676 (
            .O(N__11429),
            .I(N__11426));
    Odrv12 I__2675 (
            .O(N__11426),
            .I(mem_out_bus2_1));
    InMux I__2674 (
            .O(N__11423),
            .I(N__11420));
    LocalMux I__2673 (
            .O(N__11420),
            .I(N__11417));
    Odrv12 I__2672 (
            .O(N__11417),
            .I(mem_out_bus6_1));
    InMux I__2671 (
            .O(N__11414),
            .I(N__11411));
    LocalMux I__2670 (
            .O(N__11411),
            .I(N__11408));
    Span4Mux_v I__2669 (
            .O(N__11408),
            .I(N__11405));
    Odrv4 I__2668 (
            .O(N__11405),
            .I(dout_obuf_RNO_5Z0Z_1));
    InMux I__2667 (
            .O(N__11402),
            .I(N__11399));
    LocalMux I__2666 (
            .O(N__11399),
            .I(N__11396));
    Span4Mux_h I__2665 (
            .O(N__11396),
            .I(N__11393));
    Odrv4 I__2664 (
            .O(N__11393),
            .I(mem_out_bus6_0));
    InMux I__2663 (
            .O(N__11390),
            .I(N__11387));
    LocalMux I__2662 (
            .O(N__11387),
            .I(N__11384));
    Span4Mux_v I__2661 (
            .O(N__11384),
            .I(N__11381));
    Sp12to4 I__2660 (
            .O(N__11381),
            .I(N__11378));
    Span12Mux_h I__2659 (
            .O(N__11378),
            .I(N__11375));
    Odrv12 I__2658 (
            .O(N__11375),
            .I(mem_out_bus2_0));
    InMux I__2657 (
            .O(N__11372),
            .I(N__11369));
    LocalMux I__2656 (
            .O(N__11369),
            .I(N__11366));
    Odrv12 I__2655 (
            .O(N__11366),
            .I(dout_obuf_RNO_5Z0Z_0));
    InMux I__2654 (
            .O(N__11363),
            .I(N__11360));
    LocalMux I__2653 (
            .O(N__11360),
            .I(N__11357));
    Span4Mux_v I__2652 (
            .O(N__11357),
            .I(N__11354));
    Odrv4 I__2651 (
            .O(N__11354),
            .I(mem_out_bus6_3));
    InMux I__2650 (
            .O(N__11351),
            .I(N__11348));
    LocalMux I__2649 (
            .O(N__11348),
            .I(N__11345));
    Span4Mux_v I__2648 (
            .O(N__11345),
            .I(N__11342));
    Sp12to4 I__2647 (
            .O(N__11342),
            .I(N__11339));
    Span12Mux_h I__2646 (
            .O(N__11339),
            .I(N__11336));
    Odrv12 I__2645 (
            .O(N__11336),
            .I(mem_out_bus2_3));
    InMux I__2644 (
            .O(N__11333),
            .I(N__11330));
    LocalMux I__2643 (
            .O(N__11330),
            .I(N__11327));
    Span4Mux_h I__2642 (
            .O(N__11327),
            .I(N__11324));
    Odrv4 I__2641 (
            .O(N__11324),
            .I(mem_out_bus7_0));
    InMux I__2640 (
            .O(N__11321),
            .I(N__11318));
    LocalMux I__2639 (
            .O(N__11318),
            .I(N__11315));
    Span4Mux_v I__2638 (
            .O(N__11315),
            .I(N__11312));
    Sp12to4 I__2637 (
            .O(N__11312),
            .I(N__11309));
    Span12Mux_h I__2636 (
            .O(N__11309),
            .I(N__11306));
    Odrv12 I__2635 (
            .O(N__11306),
            .I(mem_out_bus3_0));
    InMux I__2634 (
            .O(N__11303),
            .I(N__11300));
    LocalMux I__2633 (
            .O(N__11300),
            .I(N__11297));
    Span12Mux_v I__2632 (
            .O(N__11297),
            .I(N__11294));
    Odrv12 I__2631 (
            .O(N__11294),
            .I(dout_obuf_RNO_3Z0Z_0));
    InMux I__2630 (
            .O(N__11291),
            .I(N__11288));
    LocalMux I__2629 (
            .O(N__11288),
            .I(N__11285));
    Span4Mux_h I__2628 (
            .O(N__11285),
            .I(N__11282));
    Odrv4 I__2627 (
            .O(N__11282),
            .I(mem_out_bus7_2));
    InMux I__2626 (
            .O(N__11279),
            .I(N__11276));
    LocalMux I__2625 (
            .O(N__11276),
            .I(N__11273));
    Span4Mux_v I__2624 (
            .O(N__11273),
            .I(N__11270));
    Sp12to4 I__2623 (
            .O(N__11270),
            .I(N__11267));
    Span12Mux_h I__2622 (
            .O(N__11267),
            .I(N__11264));
    Odrv12 I__2621 (
            .O(N__11264),
            .I(mem_out_bus3_2));
    InMux I__2620 (
            .O(N__11261),
            .I(N__11258));
    LocalMux I__2619 (
            .O(N__11258),
            .I(N__11255));
    Span12Mux_v I__2618 (
            .O(N__11255),
            .I(N__11252));
    Span12Mux_v I__2617 (
            .O(N__11252),
            .I(N__11249));
    Odrv12 I__2616 (
            .O(N__11249),
            .I(dout_obuf_RNO_3Z0Z_2));
    InMux I__2615 (
            .O(N__11246),
            .I(N__11243));
    LocalMux I__2614 (
            .O(N__11243),
            .I(N__11240));
    Odrv4 I__2613 (
            .O(N__11240),
            .I(mem_out_bus7_3));
    InMux I__2612 (
            .O(N__11237),
            .I(N__11234));
    LocalMux I__2611 (
            .O(N__11234),
            .I(N__11231));
    Span12Mux_h I__2610 (
            .O(N__11231),
            .I(N__11228));
    Span12Mux_h I__2609 (
            .O(N__11228),
            .I(N__11225));
    Odrv12 I__2608 (
            .O(N__11225),
            .I(mem_out_bus3_3));
    InMux I__2607 (
            .O(N__11222),
            .I(N__11219));
    LocalMux I__2606 (
            .O(N__11219),
            .I(N__11216));
    Span4Mux_s3_v I__2605 (
            .O(N__11216),
            .I(N__11213));
    Odrv4 I__2604 (
            .O(N__11213),
            .I(mem_out_bus4_2));
    InMux I__2603 (
            .O(N__11210),
            .I(N__11207));
    LocalMux I__2602 (
            .O(N__11207),
            .I(N__11204));
    Span4Mux_s3_v I__2601 (
            .O(N__11204),
            .I(N__11201));
    Sp12to4 I__2600 (
            .O(N__11201),
            .I(N__11198));
    Span12Mux_h I__2599 (
            .O(N__11198),
            .I(N__11195));
    Odrv12 I__2598 (
            .O(N__11195),
            .I(mem_out_bus0_2));
    InMux I__2597 (
            .O(N__11192),
            .I(N__11189));
    LocalMux I__2596 (
            .O(N__11189),
            .I(N__11186));
    Odrv4 I__2595 (
            .O(N__11186),
            .I(mem_out_bus4_3));
    InMux I__2594 (
            .O(N__11183),
            .I(N__11180));
    LocalMux I__2593 (
            .O(N__11180),
            .I(N__11177));
    Span12Mux_h I__2592 (
            .O(N__11177),
            .I(N__11174));
    Odrv12 I__2591 (
            .O(N__11174),
            .I(mem_out_bus0_3));
    InMux I__2590 (
            .O(N__11171),
            .I(N__11168));
    LocalMux I__2589 (
            .O(N__11168),
            .I(N__11165));
    Odrv12 I__2588 (
            .O(N__11165),
            .I(dout_obuf_RNO_2Z0Z_1));
    InMux I__2587 (
            .O(N__11162),
            .I(N__11159));
    LocalMux I__2586 (
            .O(N__11159),
            .I(mem_N_160));
    InMux I__2585 (
            .O(N__11156),
            .I(N__11153));
    LocalMux I__2584 (
            .O(N__11153),
            .I(N__11150));
    Odrv4 I__2583 (
            .O(N__11150),
            .I(dout_obuf_RNO_2Z0Z_0));
    InMux I__2582 (
            .O(N__11147),
            .I(N__11144));
    LocalMux I__2581 (
            .O(N__11144),
            .I(mem_N_154));
    InMux I__2580 (
            .O(N__11141),
            .I(N__11138));
    LocalMux I__2579 (
            .O(N__11138),
            .I(N__11135));
    Span4Mux_h I__2578 (
            .O(N__11135),
            .I(N__11132));
    Odrv4 I__2577 (
            .O(N__11132),
            .I(mem_out_bus5_2));
    InMux I__2576 (
            .O(N__11129),
            .I(N__11126));
    LocalMux I__2575 (
            .O(N__11126),
            .I(N__11123));
    Span4Mux_v I__2574 (
            .O(N__11123),
            .I(N__11120));
    Sp12to4 I__2573 (
            .O(N__11120),
            .I(N__11117));
    Span12Mux_h I__2572 (
            .O(N__11117),
            .I(N__11114));
    Odrv12 I__2571 (
            .O(N__11114),
            .I(mem_out_bus1_2));
    InMux I__2570 (
            .O(N__11111),
            .I(N__11108));
    LocalMux I__2569 (
            .O(N__11108),
            .I(dout_obuf_RNO_2Z0Z_2));
    CascadeMux I__2568 (
            .O(N__11105),
            .I(mem_N_166_cascade_));
    IoInMux I__2567 (
            .O(N__11102),
            .I(N__11099));
    LocalMux I__2566 (
            .O(N__11099),
            .I(N__11096));
    Odrv12 I__2565 (
            .O(N__11096),
            .I(dout_c_2));
    InMux I__2564 (
            .O(N__11093),
            .I(N__11090));
    LocalMux I__2563 (
            .O(N__11090),
            .I(N__11087));
    Odrv12 I__2562 (
            .O(N__11087),
            .I(dout_obuf_RNO_4Z0Z_7));
    InMux I__2561 (
            .O(N__11084),
            .I(N__11081));
    LocalMux I__2560 (
            .O(N__11081),
            .I(N__11078));
    Odrv4 I__2559 (
            .O(N__11078),
            .I(mem_out_bus5_7));
    InMux I__2558 (
            .O(N__11075),
            .I(N__11072));
    LocalMux I__2557 (
            .O(N__11072),
            .I(N__11069));
    Span12Mux_h I__2556 (
            .O(N__11069),
            .I(N__11066));
    Span12Mux_h I__2555 (
            .O(N__11066),
            .I(N__11063));
    Odrv12 I__2554 (
            .O(N__11063),
            .I(mem_out_bus1_7));
    CascadeMux I__2553 (
            .O(N__11060),
            .I(dout_obuf_RNO_2Z0Z_7_cascade_));
    InMux I__2552 (
            .O(N__11057),
            .I(N__11054));
    LocalMux I__2551 (
            .O(N__11054),
            .I(mem_N_150));
    CascadeMux I__2550 (
            .O(N__11051),
            .I(mem_N_149_cascade_));
    IoInMux I__2549 (
            .O(N__11048),
            .I(N__11045));
    LocalMux I__2548 (
            .O(N__11045),
            .I(N__11042));
    IoSpan4Mux I__2547 (
            .O(N__11042),
            .I(N__11039));
    Span4Mux_s3_h I__2546 (
            .O(N__11039),
            .I(N__11036));
    Span4Mux_h I__2545 (
            .O(N__11036),
            .I(N__11033));
    Odrv4 I__2544 (
            .O(N__11033),
            .I(dout_c_7));
    InMux I__2543 (
            .O(N__11030),
            .I(N__11027));
    LocalMux I__2542 (
            .O(N__11027),
            .I(N__11024));
    Span4Mux_v I__2541 (
            .O(N__11024),
            .I(N__11021));
    Sp12to4 I__2540 (
            .O(N__11021),
            .I(N__11018));
    Span12Mux_h I__2539 (
            .O(N__11018),
            .I(N__11015));
    Odrv12 I__2538 (
            .O(N__11015),
            .I(mem_out_bus0_6));
    InMux I__2537 (
            .O(N__11012),
            .I(N__11009));
    LocalMux I__2536 (
            .O(N__11009),
            .I(N__11006));
    Span4Mux_h I__2535 (
            .O(N__11006),
            .I(N__11003));
    Odrv4 I__2534 (
            .O(N__11003),
            .I(mem_out_bus4_6));
    SRMux I__2533 (
            .O(N__11000),
            .I(N__10995));
    SRMux I__2532 (
            .O(N__10999),
            .I(N__10992));
    SRMux I__2531 (
            .O(N__10998),
            .I(N__10987));
    LocalMux I__2530 (
            .O(N__10995),
            .I(N__10980));
    LocalMux I__2529 (
            .O(N__10992),
            .I(N__10980));
    SRMux I__2528 (
            .O(N__10991),
            .I(N__10977));
    SRMux I__2527 (
            .O(N__10990),
            .I(N__10974));
    LocalMux I__2526 (
            .O(N__10987),
            .I(N__10971));
    SRMux I__2525 (
            .O(N__10986),
            .I(N__10968));
    SRMux I__2524 (
            .O(N__10985),
            .I(N__10965));
    Span4Mux_s3_v I__2523 (
            .O(N__10980),
            .I(N__10953));
    LocalMux I__2522 (
            .O(N__10977),
            .I(N__10953));
    LocalMux I__2521 (
            .O(N__10974),
            .I(N__10953));
    Span4Mux_s3_v I__2520 (
            .O(N__10971),
            .I(N__10946));
    LocalMux I__2519 (
            .O(N__10968),
            .I(N__10946));
    LocalMux I__2518 (
            .O(N__10965),
            .I(N__10946));
    SRMux I__2517 (
            .O(N__10964),
            .I(N__10943));
    SRMux I__2516 (
            .O(N__10963),
            .I(N__10940));
    SRMux I__2515 (
            .O(N__10962),
            .I(N__10937));
    SRMux I__2514 (
            .O(N__10961),
            .I(N__10934));
    SRMux I__2513 (
            .O(N__10960),
            .I(N__10928));
    Span4Mux_v I__2512 (
            .O(N__10953),
            .I(N__10911));
    Span4Mux_v I__2511 (
            .O(N__10946),
            .I(N__10911));
    LocalMux I__2510 (
            .O(N__10943),
            .I(N__10911));
    LocalMux I__2509 (
            .O(N__10940),
            .I(N__10911));
    LocalMux I__2508 (
            .O(N__10937),
            .I(N__10906));
    LocalMux I__2507 (
            .O(N__10934),
            .I(N__10906));
    SRMux I__2506 (
            .O(N__10933),
            .I(N__10903));
    SRMux I__2505 (
            .O(N__10932),
            .I(N__10900));
    SRMux I__2504 (
            .O(N__10931),
            .I(N__10895));
    LocalMux I__2503 (
            .O(N__10928),
            .I(N__10892));
    SRMux I__2502 (
            .O(N__10927),
            .I(N__10889));
    SRMux I__2501 (
            .O(N__10926),
            .I(N__10886));
    SRMux I__2500 (
            .O(N__10925),
            .I(N__10882));
    SRMux I__2499 (
            .O(N__10924),
            .I(N__10879));
    SRMux I__2498 (
            .O(N__10923),
            .I(N__10873));
    SRMux I__2497 (
            .O(N__10922),
            .I(N__10870));
    SRMux I__2496 (
            .O(N__10921),
            .I(N__10865));
    SRMux I__2495 (
            .O(N__10920),
            .I(N__10859));
    Span4Mux_v I__2494 (
            .O(N__10911),
            .I(N__10849));
    Span4Mux_v I__2493 (
            .O(N__10906),
            .I(N__10849));
    LocalMux I__2492 (
            .O(N__10903),
            .I(N__10849));
    LocalMux I__2491 (
            .O(N__10900),
            .I(N__10849));
    SRMux I__2490 (
            .O(N__10899),
            .I(N__10846));
    SRMux I__2489 (
            .O(N__10898),
            .I(N__10843));
    LocalMux I__2488 (
            .O(N__10895),
            .I(N__10835));
    Span4Mux_s0_v I__2487 (
            .O(N__10892),
            .I(N__10835));
    LocalMux I__2486 (
            .O(N__10889),
            .I(N__10835));
    LocalMux I__2485 (
            .O(N__10886),
            .I(N__10832));
    SRMux I__2484 (
            .O(N__10885),
            .I(N__10829));
    LocalMux I__2483 (
            .O(N__10882),
            .I(N__10823));
    LocalMux I__2482 (
            .O(N__10879),
            .I(N__10823));
    SRMux I__2481 (
            .O(N__10878),
            .I(N__10820));
    SRMux I__2480 (
            .O(N__10877),
            .I(N__10817));
    SRMux I__2479 (
            .O(N__10876),
            .I(N__10813));
    LocalMux I__2478 (
            .O(N__10873),
            .I(N__10808));
    LocalMux I__2477 (
            .O(N__10870),
            .I(N__10805));
    SRMux I__2476 (
            .O(N__10869),
            .I(N__10802));
    SRMux I__2475 (
            .O(N__10868),
            .I(N__10799));
    LocalMux I__2474 (
            .O(N__10865),
            .I(N__10795));
    SRMux I__2473 (
            .O(N__10864),
            .I(N__10792));
    SRMux I__2472 (
            .O(N__10863),
            .I(N__10789));
    SRMux I__2471 (
            .O(N__10862),
            .I(N__10783));
    LocalMux I__2470 (
            .O(N__10859),
            .I(N__10780));
    SRMux I__2469 (
            .O(N__10858),
            .I(N__10777));
    Span4Mux_v I__2468 (
            .O(N__10849),
            .I(N__10770));
    LocalMux I__2467 (
            .O(N__10846),
            .I(N__10770));
    LocalMux I__2466 (
            .O(N__10843),
            .I(N__10770));
    SRMux I__2465 (
            .O(N__10842),
            .I(N__10767));
    Span4Mux_v I__2464 (
            .O(N__10835),
            .I(N__10760));
    Span4Mux_v I__2463 (
            .O(N__10832),
            .I(N__10760));
    LocalMux I__2462 (
            .O(N__10829),
            .I(N__10760));
    SRMux I__2461 (
            .O(N__10828),
            .I(N__10757));
    Span4Mux_v I__2460 (
            .O(N__10823),
            .I(N__10750));
    LocalMux I__2459 (
            .O(N__10820),
            .I(N__10750));
    LocalMux I__2458 (
            .O(N__10817),
            .I(N__10750));
    SRMux I__2457 (
            .O(N__10816),
            .I(N__10747));
    LocalMux I__2456 (
            .O(N__10813),
            .I(N__10744));
    SRMux I__2455 (
            .O(N__10812),
            .I(N__10741));
    SRMux I__2454 (
            .O(N__10811),
            .I(N__10737));
    Span4Mux_s3_v I__2453 (
            .O(N__10808),
            .I(N__10727));
    Span4Mux_s3_v I__2452 (
            .O(N__10805),
            .I(N__10727));
    LocalMux I__2451 (
            .O(N__10802),
            .I(N__10727));
    LocalMux I__2450 (
            .O(N__10799),
            .I(N__10727));
    SRMux I__2449 (
            .O(N__10798),
            .I(N__10724));
    Span4Mux_s3_v I__2448 (
            .O(N__10795),
            .I(N__10717));
    LocalMux I__2447 (
            .O(N__10792),
            .I(N__10717));
    LocalMux I__2446 (
            .O(N__10789),
            .I(N__10717));
    SRMux I__2445 (
            .O(N__10788),
            .I(N__10714));
    SRMux I__2444 (
            .O(N__10787),
            .I(N__10711));
    SRMux I__2443 (
            .O(N__10786),
            .I(N__10706));
    LocalMux I__2442 (
            .O(N__10783),
            .I(N__10696));
    Span4Mux_h I__2441 (
            .O(N__10780),
            .I(N__10696));
    LocalMux I__2440 (
            .O(N__10777),
            .I(N__10696));
    Span4Mux_v I__2439 (
            .O(N__10770),
            .I(N__10687));
    LocalMux I__2438 (
            .O(N__10767),
            .I(N__10687));
    Span4Mux_v I__2437 (
            .O(N__10760),
            .I(N__10687));
    LocalMux I__2436 (
            .O(N__10757),
            .I(N__10687));
    Span4Mux_v I__2435 (
            .O(N__10750),
            .I(N__10678));
    LocalMux I__2434 (
            .O(N__10747),
            .I(N__10678));
    Span4Mux_h I__2433 (
            .O(N__10744),
            .I(N__10678));
    LocalMux I__2432 (
            .O(N__10741),
            .I(N__10678));
    SRMux I__2431 (
            .O(N__10740),
            .I(N__10675));
    LocalMux I__2430 (
            .O(N__10737),
            .I(N__10672));
    SRMux I__2429 (
            .O(N__10736),
            .I(N__10669));
    Span4Mux_v I__2428 (
            .O(N__10727),
            .I(N__10664));
    LocalMux I__2427 (
            .O(N__10724),
            .I(N__10664));
    Span4Mux_v I__2426 (
            .O(N__10717),
            .I(N__10657));
    LocalMux I__2425 (
            .O(N__10714),
            .I(N__10657));
    LocalMux I__2424 (
            .O(N__10711),
            .I(N__10657));
    SRMux I__2423 (
            .O(N__10710),
            .I(N__10654));
    SRMux I__2422 (
            .O(N__10709),
            .I(N__10651));
    LocalMux I__2421 (
            .O(N__10706),
            .I(N__10648));
    SRMux I__2420 (
            .O(N__10705),
            .I(N__10645));
    SRMux I__2419 (
            .O(N__10704),
            .I(N__10642));
    SRMux I__2418 (
            .O(N__10703),
            .I(N__10633));
    Span4Mux_v I__2417 (
            .O(N__10696),
            .I(N__10624));
    Span4Mux_v I__2416 (
            .O(N__10687),
            .I(N__10624));
    Span4Mux_v I__2415 (
            .O(N__10678),
            .I(N__10624));
    LocalMux I__2414 (
            .O(N__10675),
            .I(N__10617));
    Span4Mux_h I__2413 (
            .O(N__10672),
            .I(N__10617));
    LocalMux I__2412 (
            .O(N__10669),
            .I(N__10617));
    Span4Mux_v I__2411 (
            .O(N__10664),
            .I(N__10608));
    Span4Mux_v I__2410 (
            .O(N__10657),
            .I(N__10608));
    LocalMux I__2409 (
            .O(N__10654),
            .I(N__10608));
    LocalMux I__2408 (
            .O(N__10651),
            .I(N__10608));
    Span4Mux_v I__2407 (
            .O(N__10648),
            .I(N__10601));
    LocalMux I__2406 (
            .O(N__10645),
            .I(N__10601));
    LocalMux I__2405 (
            .O(N__10642),
            .I(N__10601));
    SRMux I__2404 (
            .O(N__10641),
            .I(N__10598));
    SRMux I__2403 (
            .O(N__10640),
            .I(N__10595));
    SRMux I__2402 (
            .O(N__10639),
            .I(N__10591));
    SRMux I__2401 (
            .O(N__10638),
            .I(N__10586));
    SRMux I__2400 (
            .O(N__10637),
            .I(N__10583));
    SRMux I__2399 (
            .O(N__10636),
            .I(N__10579));
    LocalMux I__2398 (
            .O(N__10633),
            .I(N__10576));
    SRMux I__2397 (
            .O(N__10632),
            .I(N__10573));
    SRMux I__2396 (
            .O(N__10631),
            .I(N__10570));
    Span4Mux_h I__2395 (
            .O(N__10624),
            .I(N__10567));
    Span4Mux_v I__2394 (
            .O(N__10617),
            .I(N__10564));
    Span4Mux_v I__2393 (
            .O(N__10608),
            .I(N__10555));
    Span4Mux_v I__2392 (
            .O(N__10601),
            .I(N__10555));
    LocalMux I__2391 (
            .O(N__10598),
            .I(N__10555));
    LocalMux I__2390 (
            .O(N__10595),
            .I(N__10555));
    SRMux I__2389 (
            .O(N__10594),
            .I(N__10552));
    LocalMux I__2388 (
            .O(N__10591),
            .I(N__10549));
    SRMux I__2387 (
            .O(N__10590),
            .I(N__10546));
    SRMux I__2386 (
            .O(N__10589),
            .I(N__10543));
    LocalMux I__2385 (
            .O(N__10586),
            .I(N__10540));
    LocalMux I__2384 (
            .O(N__10583),
            .I(N__10537));
    SRMux I__2383 (
            .O(N__10582),
            .I(N__10534));
    LocalMux I__2382 (
            .O(N__10579),
            .I(N__10531));
    Span4Mux_h I__2381 (
            .O(N__10576),
            .I(N__10527));
    LocalMux I__2380 (
            .O(N__10573),
            .I(N__10524));
    LocalMux I__2379 (
            .O(N__10570),
            .I(N__10521));
    Span4Mux_h I__2378 (
            .O(N__10567),
            .I(N__10518));
    Span4Mux_v I__2377 (
            .O(N__10564),
            .I(N__10513));
    Span4Mux_v I__2376 (
            .O(N__10555),
            .I(N__10513));
    LocalMux I__2375 (
            .O(N__10552),
            .I(N__10510));
    Span4Mux_h I__2374 (
            .O(N__10549),
            .I(N__10507));
    LocalMux I__2373 (
            .O(N__10546),
            .I(N__10504));
    LocalMux I__2372 (
            .O(N__10543),
            .I(N__10501));
    Span4Mux_h I__2371 (
            .O(N__10540),
            .I(N__10496));
    Span4Mux_h I__2370 (
            .O(N__10537),
            .I(N__10496));
    LocalMux I__2369 (
            .O(N__10534),
            .I(N__10493));
    Span4Mux_h I__2368 (
            .O(N__10531),
            .I(N__10490));
    SRMux I__2367 (
            .O(N__10530),
            .I(N__10487));
    Span4Mux_v I__2366 (
            .O(N__10527),
            .I(N__10480));
    Span4Mux_h I__2365 (
            .O(N__10524),
            .I(N__10480));
    Span4Mux_h I__2364 (
            .O(N__10521),
            .I(N__10480));
    Span4Mux_h I__2363 (
            .O(N__10518),
            .I(N__10475));
    Span4Mux_v I__2362 (
            .O(N__10513),
            .I(N__10475));
    Span4Mux_h I__2361 (
            .O(N__10510),
            .I(N__10472));
    Span4Mux_v I__2360 (
            .O(N__10507),
            .I(N__10465));
    Span4Mux_h I__2359 (
            .O(N__10504),
            .I(N__10465));
    Span4Mux_h I__2358 (
            .O(N__10501),
            .I(N__10465));
    Sp12to4 I__2357 (
            .O(N__10496),
            .I(N__10460));
    Span12Mux_s9_h I__2356 (
            .O(N__10493),
            .I(N__10460));
    Span4Mux_v I__2355 (
            .O(N__10490),
            .I(N__10455));
    LocalMux I__2354 (
            .O(N__10487),
            .I(N__10455));
    Span4Mux_v I__2353 (
            .O(N__10480),
            .I(N__10452));
    Odrv4 I__2352 (
            .O(N__10475),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2351 (
            .O(N__10472),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2350 (
            .O(N__10465),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2349 (
            .O(N__10460),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2348 (
            .O(N__10455),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2347 (
            .O(N__10452),
            .I(CONSTANT_ONE_NET));
    InMux I__2346 (
            .O(N__10439),
            .I(N__10436));
    LocalMux I__2345 (
            .O(N__10436),
            .I(N__10433));
    Odrv4 I__2344 (
            .O(N__10433),
            .I(mem_out_bus5_1));
    InMux I__2343 (
            .O(N__10430),
            .I(N__10427));
    LocalMux I__2342 (
            .O(N__10427),
            .I(N__10424));
    Span12Mux_h I__2341 (
            .O(N__10424),
            .I(N__10421));
    Span12Mux_h I__2340 (
            .O(N__10421),
            .I(N__10418));
    Odrv12 I__2339 (
            .O(N__10418),
            .I(mem_out_bus1_1));
    InMux I__2338 (
            .O(N__10415),
            .I(N__10412));
    LocalMux I__2337 (
            .O(N__10412),
            .I(N__10409));
    Span4Mux_h I__2336 (
            .O(N__10409),
            .I(N__10406));
    Odrv4 I__2335 (
            .O(N__10406),
            .I(mem_out_bus5_0));
    InMux I__2334 (
            .O(N__10403),
            .I(N__10400));
    LocalMux I__2333 (
            .O(N__10400),
            .I(N__10397));
    Span4Mux_v I__2332 (
            .O(N__10397),
            .I(N__10394));
    Sp12to4 I__2331 (
            .O(N__10394),
            .I(N__10391));
    Span12Mux_h I__2330 (
            .O(N__10391),
            .I(N__10388));
    Odrv12 I__2329 (
            .O(N__10388),
            .I(mem_out_bus1_0));
    InMux I__2328 (
            .O(N__10385),
            .I(N__10382));
    LocalMux I__2327 (
            .O(N__10382),
            .I(N__10379));
    Span12Mux_v I__2326 (
            .O(N__10379),
            .I(N__10376));
    Odrv12 I__2325 (
            .O(N__10376),
            .I(dout_obuf_RNO_4Z0Z_1));
    CascadeMux I__2324 (
            .O(N__10373),
            .I(mem_N_162_cascade_));
    IoInMux I__2323 (
            .O(N__10370),
            .I(N__10367));
    LocalMux I__2322 (
            .O(N__10367),
            .I(N__10364));
    Span12Mux_s9_h I__2321 (
            .O(N__10364),
            .I(N__10361));
    Odrv12 I__2320 (
            .O(N__10361),
            .I(dout_c_1));
    InMux I__2319 (
            .O(N__10358),
            .I(N__10355));
    LocalMux I__2318 (
            .O(N__10355),
            .I(N__10352));
    Span12Mux_v I__2317 (
            .O(N__10352),
            .I(N__10349));
    Odrv12 I__2316 (
            .O(N__10349),
            .I(dout_obuf_RNO_4Z0Z_0));
    CascadeMux I__2315 (
            .O(N__10346),
            .I(mem_N_156_cascade_));
    IoInMux I__2314 (
            .O(N__10343),
            .I(N__10340));
    LocalMux I__2313 (
            .O(N__10340),
            .I(N__10337));
    Span4Mux_s2_h I__2312 (
            .O(N__10337),
            .I(N__10334));
    Sp12to4 I__2311 (
            .O(N__10334),
            .I(N__10331));
    Span12Mux_s10_v I__2310 (
            .O(N__10331),
            .I(N__10328));
    Odrv12 I__2309 (
            .O(N__10328),
            .I(dout_c_0));
    CEMux I__2308 (
            .O(N__10325),
            .I(N__10321));
    CEMux I__2307 (
            .O(N__10324),
            .I(N__10318));
    LocalMux I__2306 (
            .O(N__10321),
            .I(N__10314));
    LocalMux I__2305 (
            .O(N__10318),
            .I(N__10311));
    CEMux I__2304 (
            .O(N__10317),
            .I(N__10308));
    Span4Mux_v I__2303 (
            .O(N__10314),
            .I(N__10301));
    Span4Mux_h I__2302 (
            .O(N__10311),
            .I(N__10301));
    LocalMux I__2301 (
            .O(N__10308),
            .I(N__10301));
    Span4Mux_v I__2300 (
            .O(N__10301),
            .I(N__10297));
    CEMux I__2299 (
            .O(N__10300),
            .I(N__10294));
    Odrv4 I__2298 (
            .O(N__10297),
            .I(mem_WE_8));
    LocalMux I__2297 (
            .O(N__10294),
            .I(mem_WE_8));
    CEMux I__2296 (
            .O(N__10289),
            .I(N__10285));
    CEMux I__2295 (
            .O(N__10288),
            .I(N__10282));
    LocalMux I__2294 (
            .O(N__10285),
            .I(N__10276));
    LocalMux I__2293 (
            .O(N__10282),
            .I(N__10276));
    CEMux I__2292 (
            .O(N__10281),
            .I(N__10273));
    Span4Mux_v I__2291 (
            .O(N__10276),
            .I(N__10267));
    LocalMux I__2290 (
            .O(N__10273),
            .I(N__10267));
    CEMux I__2289 (
            .O(N__10272),
            .I(N__10264));
    Span4Mux_v I__2288 (
            .O(N__10267),
            .I(N__10261));
    LocalMux I__2287 (
            .O(N__10264),
            .I(N__10258));
    Span4Mux_v I__2286 (
            .O(N__10261),
            .I(N__10255));
    Span12Mux_h I__2285 (
            .O(N__10258),
            .I(N__10252));
    Odrv4 I__2284 (
            .O(N__10255),
            .I(mem_WE_12));
    Odrv12 I__2283 (
            .O(N__10252),
            .I(mem_WE_12));
    CEMux I__2282 (
            .O(N__10247),
            .I(N__10243));
    CEMux I__2281 (
            .O(N__10246),
            .I(N__10240));
    LocalMux I__2280 (
            .O(N__10243),
            .I(N__10233));
    LocalMux I__2279 (
            .O(N__10240),
            .I(N__10233));
    CEMux I__2278 (
            .O(N__10239),
            .I(N__10230));
    CEMux I__2277 (
            .O(N__10238),
            .I(N__10227));
    Span4Mux_s3_v I__2276 (
            .O(N__10233),
            .I(N__10220));
    LocalMux I__2275 (
            .O(N__10230),
            .I(N__10220));
    LocalMux I__2274 (
            .O(N__10227),
            .I(N__10220));
    Span4Mux_v I__2273 (
            .O(N__10220),
            .I(N__10217));
    Span4Mux_v I__2272 (
            .O(N__10217),
            .I(N__10214));
    Span4Mux_v I__2271 (
            .O(N__10214),
            .I(N__10211));
    Sp12to4 I__2270 (
            .O(N__10211),
            .I(N__10208));
    Span12Mux_h I__2269 (
            .O(N__10208),
            .I(N__10205));
    Odrv12 I__2268 (
            .O(N__10205),
            .I(mem_WE_16));
    CEMux I__2267 (
            .O(N__10202),
            .I(N__10199));
    LocalMux I__2266 (
            .O(N__10199),
            .I(N__10193));
    CEMux I__2265 (
            .O(N__10198),
            .I(N__10190));
    CEMux I__2264 (
            .O(N__10197),
            .I(N__10187));
    CEMux I__2263 (
            .O(N__10196),
            .I(N__10184));
    Span4Mux_v I__2262 (
            .O(N__10193),
            .I(N__10181));
    LocalMux I__2261 (
            .O(N__10190),
            .I(N__10178));
    LocalMux I__2260 (
            .O(N__10187),
            .I(N__10173));
    LocalMux I__2259 (
            .O(N__10184),
            .I(N__10173));
    Span4Mux_h I__2258 (
            .O(N__10181),
            .I(N__10168));
    Span4Mux_h I__2257 (
            .O(N__10178),
            .I(N__10168));
    Span4Mux_v I__2256 (
            .O(N__10173),
            .I(N__10165));
    Span4Mux_h I__2255 (
            .O(N__10168),
            .I(N__10162));
    Span4Mux_h I__2254 (
            .O(N__10165),
            .I(N__10159));
    Sp12to4 I__2253 (
            .O(N__10162),
            .I(N__10156));
    Sp12to4 I__2252 (
            .O(N__10159),
            .I(N__10153));
    Span12Mux_v I__2251 (
            .O(N__10156),
            .I(N__10148));
    Span12Mux_h I__2250 (
            .O(N__10153),
            .I(N__10148));
    Odrv12 I__2249 (
            .O(N__10148),
            .I(mem_WE_20));
    CEMux I__2248 (
            .O(N__10145),
            .I(N__10141));
    CEMux I__2247 (
            .O(N__10144),
            .I(N__10138));
    LocalMux I__2246 (
            .O(N__10141),
            .I(N__10131));
    LocalMux I__2245 (
            .O(N__10138),
            .I(N__10131));
    CEMux I__2244 (
            .O(N__10137),
            .I(N__10128));
    CEMux I__2243 (
            .O(N__10136),
            .I(N__10125));
    Span4Mux_v I__2242 (
            .O(N__10131),
            .I(N__10118));
    LocalMux I__2241 (
            .O(N__10128),
            .I(N__10118));
    LocalMux I__2240 (
            .O(N__10125),
            .I(N__10118));
    Span4Mux_v I__2239 (
            .O(N__10118),
            .I(N__10115));
    Span4Mux_h I__2238 (
            .O(N__10115),
            .I(N__10112));
    Span4Mux_h I__2237 (
            .O(N__10112),
            .I(N__10109));
    Span4Mux_h I__2236 (
            .O(N__10109),
            .I(N__10106));
    Span4Mux_h I__2235 (
            .O(N__10106),
            .I(N__10103));
    Odrv4 I__2234 (
            .O(N__10103),
            .I(mem_WE_24));
    InMux I__2233 (
            .O(N__10100),
            .I(N__10076));
    InMux I__2232 (
            .O(N__10099),
            .I(N__10076));
    InMux I__2231 (
            .O(N__10098),
            .I(N__10076));
    InMux I__2230 (
            .O(N__10097),
            .I(N__10076));
    InMux I__2229 (
            .O(N__10096),
            .I(N__10076));
    InMux I__2228 (
            .O(N__10095),
            .I(N__10076));
    InMux I__2227 (
            .O(N__10094),
            .I(N__10076));
    InMux I__2226 (
            .O(N__10093),
            .I(N__10076));
    LocalMux I__2225 (
            .O(N__10076),
            .I(N__10073));
    Span4Mux_v I__2224 (
            .O(N__10073),
            .I(N__10070));
    Span4Mux_h I__2223 (
            .O(N__10070),
            .I(N__10067));
    Odrv4 I__2222 (
            .O(N__10067),
            .I(write_en_c));
    InMux I__2221 (
            .O(N__10064),
            .I(N__10040));
    InMux I__2220 (
            .O(N__10063),
            .I(N__10040));
    InMux I__2219 (
            .O(N__10062),
            .I(N__10040));
    InMux I__2218 (
            .O(N__10061),
            .I(N__10040));
    InMux I__2217 (
            .O(N__10060),
            .I(N__10040));
    InMux I__2216 (
            .O(N__10059),
            .I(N__10040));
    InMux I__2215 (
            .O(N__10058),
            .I(N__10040));
    InMux I__2214 (
            .O(N__10057),
            .I(N__10040));
    LocalMux I__2213 (
            .O(N__10040),
            .I(N__10037));
    Span4Mux_v I__2212 (
            .O(N__10037),
            .I(N__10034));
    Sp12to4 I__2211 (
            .O(N__10034),
            .I(N__10031));
    Odrv12 I__2210 (
            .O(N__10031),
            .I(waddr_c_13));
    CascadeMux I__2209 (
            .O(N__10028),
            .I(N__10022));
    CascadeMux I__2208 (
            .O(N__10027),
            .I(N__10018));
    CascadeMux I__2207 (
            .O(N__10026),
            .I(N__10014));
    CascadeMux I__2206 (
            .O(N__10025),
            .I(N__10010));
    InMux I__2205 (
            .O(N__10022),
            .I(N__9992));
    InMux I__2204 (
            .O(N__10021),
            .I(N__9992));
    InMux I__2203 (
            .O(N__10018),
            .I(N__9992));
    InMux I__2202 (
            .O(N__10017),
            .I(N__9992));
    InMux I__2201 (
            .O(N__10014),
            .I(N__9992));
    InMux I__2200 (
            .O(N__10013),
            .I(N__9992));
    InMux I__2199 (
            .O(N__10010),
            .I(N__9992));
    InMux I__2198 (
            .O(N__10009),
            .I(N__9992));
    LocalMux I__2197 (
            .O(N__9992),
            .I(N__9989));
    Span4Mux_v I__2196 (
            .O(N__9989),
            .I(N__9986));
    Span4Mux_h I__2195 (
            .O(N__9986),
            .I(N__9983));
    Odrv4 I__2194 (
            .O(N__9983),
            .I(waddr_c_11));
    CascadeMux I__2193 (
            .O(N__9980),
            .I(N__9973));
    CascadeMux I__2192 (
            .O(N__9979),
            .I(N__9969));
    CascadeMux I__2191 (
            .O(N__9978),
            .I(N__9965));
    CascadeMux I__2190 (
            .O(N__9977),
            .I(N__9961));
    InMux I__2189 (
            .O(N__9976),
            .I(N__9944));
    InMux I__2188 (
            .O(N__9973),
            .I(N__9944));
    InMux I__2187 (
            .O(N__9972),
            .I(N__9944));
    InMux I__2186 (
            .O(N__9969),
            .I(N__9944));
    InMux I__2185 (
            .O(N__9968),
            .I(N__9944));
    InMux I__2184 (
            .O(N__9965),
            .I(N__9944));
    InMux I__2183 (
            .O(N__9964),
            .I(N__9944));
    InMux I__2182 (
            .O(N__9961),
            .I(N__9944));
    LocalMux I__2181 (
            .O(N__9944),
            .I(N__9941));
    Odrv12 I__2180 (
            .O(N__9941),
            .I(waddr_c_12));
    CEMux I__2179 (
            .O(N__9938),
            .I(N__9932));
    CEMux I__2178 (
            .O(N__9937),
            .I(N__9929));
    CEMux I__2177 (
            .O(N__9936),
            .I(N__9926));
    CEMux I__2176 (
            .O(N__9935),
            .I(N__9923));
    LocalMux I__2175 (
            .O(N__9932),
            .I(N__9918));
    LocalMux I__2174 (
            .O(N__9929),
            .I(N__9918));
    LocalMux I__2173 (
            .O(N__9926),
            .I(N__9913));
    LocalMux I__2172 (
            .O(N__9923),
            .I(N__9913));
    Span4Mux_v I__2171 (
            .O(N__9918),
            .I(N__9908));
    Span4Mux_v I__2170 (
            .O(N__9913),
            .I(N__9908));
    Sp12to4 I__2169 (
            .O(N__9908),
            .I(N__9905));
    Span12Mux_h I__2168 (
            .O(N__9905),
            .I(N__9902));
    Span12Mux_v I__2167 (
            .O(N__9902),
            .I(N__9899));
    Odrv12 I__2166 (
            .O(N__9899),
            .I(mem_WE_28));
    InMux I__2165 (
            .O(N__9896),
            .I(N__9893));
    LocalMux I__2164 (
            .O(N__9893),
            .I(N__9890));
    Span4Mux_s1_v I__2163 (
            .O(N__9890),
            .I(N__9887));
    Sp12to4 I__2162 (
            .O(N__9887),
            .I(N__9884));
    Span12Mux_h I__2161 (
            .O(N__9884),
            .I(N__9881));
    Odrv12 I__2160 (
            .O(N__9881),
            .I(mem_out_bus0_0));
    InMux I__2159 (
            .O(N__9878),
            .I(N__9875));
    LocalMux I__2158 (
            .O(N__9875),
            .I(N__9872));
    Span4Mux_s1_v I__2157 (
            .O(N__9872),
            .I(N__9869));
    Odrv4 I__2156 (
            .O(N__9869),
            .I(mem_out_bus4_0));
    InMux I__2155 (
            .O(N__9866),
            .I(N__9863));
    LocalMux I__2154 (
            .O(N__9863),
            .I(N__9860));
    Span12Mux_h I__2153 (
            .O(N__9860),
            .I(N__9857));
    Span12Mux_h I__2152 (
            .O(N__9857),
            .I(N__9854));
    Odrv12 I__2151 (
            .O(N__9854),
            .I(mem_out_bus0_1));
    InMux I__2150 (
            .O(N__9851),
            .I(N__9848));
    LocalMux I__2149 (
            .O(N__9848),
            .I(N__9845));
    Odrv4 I__2148 (
            .O(N__9845),
            .I(mem_out_bus4_1));
    InMux I__2147 (
            .O(N__9842),
            .I(N__9839));
    LocalMux I__2146 (
            .O(N__9839),
            .I(N__9836));
    Odrv12 I__2145 (
            .O(N__9836),
            .I(mem_out_bus4_7));
    InMux I__2144 (
            .O(N__9833),
            .I(N__9830));
    LocalMux I__2143 (
            .O(N__9830),
            .I(N__9827));
    Span12Mux_h I__2142 (
            .O(N__9827),
            .I(N__9824));
    Odrv12 I__2141 (
            .O(N__9824),
            .I(mem_out_bus0_7));
    CascadeMux I__2140 (
            .O(N__9821),
            .I(N__9818));
    CascadeBuf I__2139 (
            .O(N__9818),
            .I(N__9815));
    CascadeMux I__2138 (
            .O(N__9815),
            .I(N__9811));
    CascadeMux I__2137 (
            .O(N__9814),
            .I(N__9808));
    CascadeBuf I__2136 (
            .O(N__9811),
            .I(N__9805));
    CascadeBuf I__2135 (
            .O(N__9808),
            .I(N__9802));
    CascadeMux I__2134 (
            .O(N__9805),
            .I(N__9799));
    CascadeMux I__2133 (
            .O(N__9802),
            .I(N__9796));
    CascadeBuf I__2132 (
            .O(N__9799),
            .I(N__9793));
    CascadeBuf I__2131 (
            .O(N__9796),
            .I(N__9790));
    CascadeMux I__2130 (
            .O(N__9793),
            .I(N__9787));
    CascadeMux I__2129 (
            .O(N__9790),
            .I(N__9784));
    CascadeBuf I__2128 (
            .O(N__9787),
            .I(N__9781));
    CascadeBuf I__2127 (
            .O(N__9784),
            .I(N__9778));
    CascadeMux I__2126 (
            .O(N__9781),
            .I(N__9775));
    CascadeMux I__2125 (
            .O(N__9778),
            .I(N__9772));
    CascadeBuf I__2124 (
            .O(N__9775),
            .I(N__9769));
    CascadeBuf I__2123 (
            .O(N__9772),
            .I(N__9766));
    CascadeMux I__2122 (
            .O(N__9769),
            .I(N__9763));
    CascadeMux I__2121 (
            .O(N__9766),
            .I(N__9760));
    CascadeBuf I__2120 (
            .O(N__9763),
            .I(N__9757));
    CascadeBuf I__2119 (
            .O(N__9760),
            .I(N__9754));
    CascadeMux I__2118 (
            .O(N__9757),
            .I(N__9751));
    CascadeMux I__2117 (
            .O(N__9754),
            .I(N__9748));
    CascadeBuf I__2116 (
            .O(N__9751),
            .I(N__9745));
    CascadeBuf I__2115 (
            .O(N__9748),
            .I(N__9742));
    CascadeMux I__2114 (
            .O(N__9745),
            .I(N__9739));
    CascadeMux I__2113 (
            .O(N__9742),
            .I(N__9736));
    CascadeBuf I__2112 (
            .O(N__9739),
            .I(N__9733));
    CascadeBuf I__2111 (
            .O(N__9736),
            .I(N__9730));
    CascadeMux I__2110 (
            .O(N__9733),
            .I(N__9727));
    CascadeMux I__2109 (
            .O(N__9730),
            .I(N__9724));
    CascadeBuf I__2108 (
            .O(N__9727),
            .I(N__9721));
    CascadeBuf I__2107 (
            .O(N__9724),
            .I(N__9718));
    CascadeMux I__2106 (
            .O(N__9721),
            .I(N__9715));
    CascadeMux I__2105 (
            .O(N__9718),
            .I(N__9712));
    CascadeBuf I__2104 (
            .O(N__9715),
            .I(N__9709));
    CascadeBuf I__2103 (
            .O(N__9712),
            .I(N__9706));
    CascadeMux I__2102 (
            .O(N__9709),
            .I(N__9703));
    CascadeMux I__2101 (
            .O(N__9706),
            .I(N__9700));
    CascadeBuf I__2100 (
            .O(N__9703),
            .I(N__9697));
    CascadeBuf I__2099 (
            .O(N__9700),
            .I(N__9694));
    CascadeMux I__2098 (
            .O(N__9697),
            .I(N__9691));
    CascadeMux I__2097 (
            .O(N__9694),
            .I(N__9688));
    CascadeBuf I__2096 (
            .O(N__9691),
            .I(N__9685));
    CascadeBuf I__2095 (
            .O(N__9688),
            .I(N__9682));
    CascadeMux I__2094 (
            .O(N__9685),
            .I(N__9679));
    CascadeMux I__2093 (
            .O(N__9682),
            .I(N__9676));
    CascadeBuf I__2092 (
            .O(N__9679),
            .I(N__9673));
    CascadeBuf I__2091 (
            .O(N__9676),
            .I(N__9670));
    CascadeMux I__2090 (
            .O(N__9673),
            .I(N__9667));
    CascadeMux I__2089 (
            .O(N__9670),
            .I(N__9664));
    CascadeBuf I__2088 (
            .O(N__9667),
            .I(N__9661));
    CascadeBuf I__2087 (
            .O(N__9664),
            .I(N__9658));
    CascadeMux I__2086 (
            .O(N__9661),
            .I(N__9655));
    CascadeMux I__2085 (
            .O(N__9658),
            .I(N__9652));
    CascadeBuf I__2084 (
            .O(N__9655),
            .I(N__9649));
    CascadeBuf I__2083 (
            .O(N__9652),
            .I(N__9646));
    CascadeMux I__2082 (
            .O(N__9649),
            .I(N__9643));
    CascadeMux I__2081 (
            .O(N__9646),
            .I(N__9640));
    InMux I__2080 (
            .O(N__9643),
            .I(N__9637));
    CascadeBuf I__2079 (
            .O(N__9640),
            .I(N__9634));
    LocalMux I__2078 (
            .O(N__9637),
            .I(N__9631));
    CascadeMux I__2077 (
            .O(N__9634),
            .I(N__9628));
    Span4Mux_s2_v I__2076 (
            .O(N__9631),
            .I(N__9625));
    InMux I__2075 (
            .O(N__9628),
            .I(N__9622));
    Span4Mux_h I__2074 (
            .O(N__9625),
            .I(N__9619));
    LocalMux I__2073 (
            .O(N__9622),
            .I(N__9616));
    Sp12to4 I__2072 (
            .O(N__9619),
            .I(N__9613));
    Span4Mux_s2_v I__2071 (
            .O(N__9616),
            .I(N__9610));
    Span12Mux_h I__2070 (
            .O(N__9613),
            .I(N__9605));
    Sp12to4 I__2069 (
            .O(N__9610),
            .I(N__9605));
    Odrv12 I__2068 (
            .O(N__9605),
            .I(waddr_c_0));
    CEMux I__2067 (
            .O(N__9602),
            .I(N__9599));
    LocalMux I__2066 (
            .O(N__9599),
            .I(N__9594));
    CEMux I__2065 (
            .O(N__9598),
            .I(N__9591));
    CEMux I__2064 (
            .O(N__9597),
            .I(N__9588));
    Span4Mux_v I__2063 (
            .O(N__9594),
            .I(N__9580));
    LocalMux I__2062 (
            .O(N__9591),
            .I(N__9580));
    LocalMux I__2061 (
            .O(N__9588),
            .I(N__9580));
    CEMux I__2060 (
            .O(N__9587),
            .I(N__9577));
    Span4Mux_v I__2059 (
            .O(N__9580),
            .I(N__9572));
    LocalMux I__2058 (
            .O(N__9577),
            .I(N__9572));
    Span4Mux_h I__2057 (
            .O(N__9572),
            .I(N__9569));
    Odrv4 I__2056 (
            .O(N__9569),
            .I(mem_WE_4));
    CEMux I__2055 (
            .O(N__9566),
            .I(N__9562));
    CEMux I__2054 (
            .O(N__9565),
            .I(N__9559));
    LocalMux I__2053 (
            .O(N__9562),
            .I(N__9555));
    LocalMux I__2052 (
            .O(N__9559),
            .I(N__9552));
    CEMux I__2051 (
            .O(N__9558),
            .I(N__9549));
    Span4Mux_s2_v I__2050 (
            .O(N__9555),
            .I(N__9542));
    Span4Mux_h I__2049 (
            .O(N__9552),
            .I(N__9542));
    LocalMux I__2048 (
            .O(N__9549),
            .I(N__9542));
    Span4Mux_v I__2047 (
            .O(N__9542),
            .I(N__9538));
    CEMux I__2046 (
            .O(N__9541),
            .I(N__9535));
    Sp12to4 I__2045 (
            .O(N__9538),
            .I(N__9530));
    LocalMux I__2044 (
            .O(N__9535),
            .I(N__9530));
    Span12Mux_h I__2043 (
            .O(N__9530),
            .I(N__9527));
    Odrv12 I__2042 (
            .O(N__9527),
            .I(mem_WE_0));
    InMux I__2041 (
            .O(N__9524),
            .I(N__9517));
    InMux I__2040 (
            .O(N__9523),
            .I(N__9513));
    InMux I__2039 (
            .O(N__9522),
            .I(N__9510));
    InMux I__2038 (
            .O(N__9521),
            .I(N__9507));
    InMux I__2037 (
            .O(N__9520),
            .I(N__9504));
    LocalMux I__2036 (
            .O(N__9517),
            .I(N__9501));
    InMux I__2035 (
            .O(N__9516),
            .I(N__9498));
    LocalMux I__2034 (
            .O(N__9513),
            .I(N__9494));
    LocalMux I__2033 (
            .O(N__9510),
            .I(N__9491));
    LocalMux I__2032 (
            .O(N__9507),
            .I(N__9488));
    LocalMux I__2031 (
            .O(N__9504),
            .I(N__9484));
    Sp12to4 I__2030 (
            .O(N__9501),
            .I(N__9479));
    LocalMux I__2029 (
            .O(N__9498),
            .I(N__9479));
    InMux I__2028 (
            .O(N__9497),
            .I(N__9476));
    Span4Mux_h I__2027 (
            .O(N__9494),
            .I(N__9473));
    Span12Mux_h I__2026 (
            .O(N__9491),
            .I(N__9468));
    Span12Mux_h I__2025 (
            .O(N__9488),
            .I(N__9468));
    InMux I__2024 (
            .O(N__9487),
            .I(N__9465));
    Span12Mux_h I__2023 (
            .O(N__9484),
            .I(N__9462));
    Span12Mux_v I__2022 (
            .O(N__9479),
            .I(N__9459));
    LocalMux I__2021 (
            .O(N__9476),
            .I(N__9456));
    Span4Mux_h I__2020 (
            .O(N__9473),
            .I(N__9453));
    Span12Mux_v I__2019 (
            .O(N__9468),
            .I(N__9450));
    LocalMux I__2018 (
            .O(N__9465),
            .I(N__9447));
    Span12Mux_v I__2017 (
            .O(N__9462),
            .I(N__9442));
    Span12Mux_h I__2016 (
            .O(N__9459),
            .I(N__9442));
    Span12Mux_h I__2015 (
            .O(N__9456),
            .I(N__9439));
    Span4Mux_h I__2014 (
            .O(N__9453),
            .I(N__9436));
    Span12Mux_v I__2013 (
            .O(N__9450),
            .I(N__9431));
    Span12Mux_h I__2012 (
            .O(N__9447),
            .I(N__9431));
    Odrv12 I__2011 (
            .O(N__9442),
            .I(din_c_5));
    Odrv12 I__2010 (
            .O(N__9439),
            .I(din_c_5));
    Odrv4 I__2009 (
            .O(N__9436),
            .I(din_c_5));
    Odrv12 I__2008 (
            .O(N__9431),
            .I(din_c_5));
    CascadeMux I__2007 (
            .O(N__9422),
            .I(N__9419));
    CascadeBuf I__2006 (
            .O(N__9419),
            .I(N__9416));
    CascadeMux I__2005 (
            .O(N__9416),
            .I(N__9413));
    CascadeBuf I__2004 (
            .O(N__9413),
            .I(N__9409));
    CascadeMux I__2003 (
            .O(N__9412),
            .I(N__9406));
    CascadeMux I__2002 (
            .O(N__9409),
            .I(N__9403));
    CascadeBuf I__2001 (
            .O(N__9406),
            .I(N__9400));
    CascadeBuf I__2000 (
            .O(N__9403),
            .I(N__9397));
    CascadeMux I__1999 (
            .O(N__9400),
            .I(N__9394));
    CascadeMux I__1998 (
            .O(N__9397),
            .I(N__9391));
    CascadeBuf I__1997 (
            .O(N__9394),
            .I(N__9388));
    CascadeBuf I__1996 (
            .O(N__9391),
            .I(N__9385));
    CascadeMux I__1995 (
            .O(N__9388),
            .I(N__9382));
    CascadeMux I__1994 (
            .O(N__9385),
            .I(N__9379));
    CascadeBuf I__1993 (
            .O(N__9382),
            .I(N__9376));
    CascadeBuf I__1992 (
            .O(N__9379),
            .I(N__9373));
    CascadeMux I__1991 (
            .O(N__9376),
            .I(N__9370));
    CascadeMux I__1990 (
            .O(N__9373),
            .I(N__9367));
    CascadeBuf I__1989 (
            .O(N__9370),
            .I(N__9364));
    CascadeBuf I__1988 (
            .O(N__9367),
            .I(N__9361));
    CascadeMux I__1987 (
            .O(N__9364),
            .I(N__9358));
    CascadeMux I__1986 (
            .O(N__9361),
            .I(N__9355));
    CascadeBuf I__1985 (
            .O(N__9358),
            .I(N__9352));
    CascadeBuf I__1984 (
            .O(N__9355),
            .I(N__9349));
    CascadeMux I__1983 (
            .O(N__9352),
            .I(N__9346));
    CascadeMux I__1982 (
            .O(N__9349),
            .I(N__9343));
    CascadeBuf I__1981 (
            .O(N__9346),
            .I(N__9340));
    CascadeBuf I__1980 (
            .O(N__9343),
            .I(N__9337));
    CascadeMux I__1979 (
            .O(N__9340),
            .I(N__9334));
    CascadeMux I__1978 (
            .O(N__9337),
            .I(N__9331));
    CascadeBuf I__1977 (
            .O(N__9334),
            .I(N__9328));
    CascadeBuf I__1976 (
            .O(N__9331),
            .I(N__9325));
    CascadeMux I__1975 (
            .O(N__9328),
            .I(N__9322));
    CascadeMux I__1974 (
            .O(N__9325),
            .I(N__9319));
    CascadeBuf I__1973 (
            .O(N__9322),
            .I(N__9316));
    CascadeBuf I__1972 (
            .O(N__9319),
            .I(N__9313));
    CascadeMux I__1971 (
            .O(N__9316),
            .I(N__9310));
    CascadeMux I__1970 (
            .O(N__9313),
            .I(N__9307));
    CascadeBuf I__1969 (
            .O(N__9310),
            .I(N__9304));
    CascadeBuf I__1968 (
            .O(N__9307),
            .I(N__9301));
    CascadeMux I__1967 (
            .O(N__9304),
            .I(N__9298));
    CascadeMux I__1966 (
            .O(N__9301),
            .I(N__9295));
    CascadeBuf I__1965 (
            .O(N__9298),
            .I(N__9292));
    CascadeBuf I__1964 (
            .O(N__9295),
            .I(N__9289));
    CascadeMux I__1963 (
            .O(N__9292),
            .I(N__9286));
    CascadeMux I__1962 (
            .O(N__9289),
            .I(N__9283));
    CascadeBuf I__1961 (
            .O(N__9286),
            .I(N__9280));
    CascadeBuf I__1960 (
            .O(N__9283),
            .I(N__9277));
    CascadeMux I__1959 (
            .O(N__9280),
            .I(N__9274));
    CascadeMux I__1958 (
            .O(N__9277),
            .I(N__9271));
    CascadeBuf I__1957 (
            .O(N__9274),
            .I(N__9268));
    CascadeBuf I__1956 (
            .O(N__9271),
            .I(N__9265));
    CascadeMux I__1955 (
            .O(N__9268),
            .I(N__9262));
    CascadeMux I__1954 (
            .O(N__9265),
            .I(N__9259));
    CascadeBuf I__1953 (
            .O(N__9262),
            .I(N__9256));
    CascadeBuf I__1952 (
            .O(N__9259),
            .I(N__9253));
    CascadeMux I__1951 (
            .O(N__9256),
            .I(N__9250));
    CascadeMux I__1950 (
            .O(N__9253),
            .I(N__9247));
    CascadeBuf I__1949 (
            .O(N__9250),
            .I(N__9244));
    InMux I__1948 (
            .O(N__9247),
            .I(N__9241));
    CascadeMux I__1947 (
            .O(N__9244),
            .I(N__9238));
    LocalMux I__1946 (
            .O(N__9241),
            .I(N__9235));
    CascadeBuf I__1945 (
            .O(N__9238),
            .I(N__9232));
    Span4Mux_s3_v I__1944 (
            .O(N__9235),
            .I(N__9229));
    CascadeMux I__1943 (
            .O(N__9232),
            .I(N__9226));
    Span4Mux_v I__1942 (
            .O(N__9229),
            .I(N__9223));
    InMux I__1941 (
            .O(N__9226),
            .I(N__9220));
    Sp12to4 I__1940 (
            .O(N__9223),
            .I(N__9217));
    LocalMux I__1939 (
            .O(N__9220),
            .I(N__9214));
    Span12Mux_h I__1938 (
            .O(N__9217),
            .I(N__9211));
    Span12Mux_s7_v I__1937 (
            .O(N__9214),
            .I(N__9208));
    Odrv12 I__1936 (
            .O(N__9211),
            .I(raddr_c_5));
    Odrv12 I__1935 (
            .O(N__9208),
            .I(raddr_c_5));
    CascadeMux I__1934 (
            .O(N__9203),
            .I(N__9200));
    CascadeBuf I__1933 (
            .O(N__9200),
            .I(N__9197));
    CascadeMux I__1932 (
            .O(N__9197),
            .I(N__9194));
    CascadeBuf I__1931 (
            .O(N__9194),
            .I(N__9190));
    CascadeMux I__1930 (
            .O(N__9193),
            .I(N__9187));
    CascadeMux I__1929 (
            .O(N__9190),
            .I(N__9184));
    CascadeBuf I__1928 (
            .O(N__9187),
            .I(N__9181));
    CascadeBuf I__1927 (
            .O(N__9184),
            .I(N__9178));
    CascadeMux I__1926 (
            .O(N__9181),
            .I(N__9175));
    CascadeMux I__1925 (
            .O(N__9178),
            .I(N__9172));
    CascadeBuf I__1924 (
            .O(N__9175),
            .I(N__9169));
    CascadeBuf I__1923 (
            .O(N__9172),
            .I(N__9166));
    CascadeMux I__1922 (
            .O(N__9169),
            .I(N__9163));
    CascadeMux I__1921 (
            .O(N__9166),
            .I(N__9160));
    CascadeBuf I__1920 (
            .O(N__9163),
            .I(N__9157));
    CascadeBuf I__1919 (
            .O(N__9160),
            .I(N__9154));
    CascadeMux I__1918 (
            .O(N__9157),
            .I(N__9151));
    CascadeMux I__1917 (
            .O(N__9154),
            .I(N__9148));
    CascadeBuf I__1916 (
            .O(N__9151),
            .I(N__9145));
    CascadeBuf I__1915 (
            .O(N__9148),
            .I(N__9142));
    CascadeMux I__1914 (
            .O(N__9145),
            .I(N__9139));
    CascadeMux I__1913 (
            .O(N__9142),
            .I(N__9136));
    CascadeBuf I__1912 (
            .O(N__9139),
            .I(N__9133));
    CascadeBuf I__1911 (
            .O(N__9136),
            .I(N__9130));
    CascadeMux I__1910 (
            .O(N__9133),
            .I(N__9127));
    CascadeMux I__1909 (
            .O(N__9130),
            .I(N__9124));
    CascadeBuf I__1908 (
            .O(N__9127),
            .I(N__9121));
    CascadeBuf I__1907 (
            .O(N__9124),
            .I(N__9118));
    CascadeMux I__1906 (
            .O(N__9121),
            .I(N__9115));
    CascadeMux I__1905 (
            .O(N__9118),
            .I(N__9112));
    CascadeBuf I__1904 (
            .O(N__9115),
            .I(N__9109));
    CascadeBuf I__1903 (
            .O(N__9112),
            .I(N__9106));
    CascadeMux I__1902 (
            .O(N__9109),
            .I(N__9103));
    CascadeMux I__1901 (
            .O(N__9106),
            .I(N__9100));
    CascadeBuf I__1900 (
            .O(N__9103),
            .I(N__9097));
    CascadeBuf I__1899 (
            .O(N__9100),
            .I(N__9094));
    CascadeMux I__1898 (
            .O(N__9097),
            .I(N__9091));
    CascadeMux I__1897 (
            .O(N__9094),
            .I(N__9088));
    CascadeBuf I__1896 (
            .O(N__9091),
            .I(N__9085));
    CascadeBuf I__1895 (
            .O(N__9088),
            .I(N__9082));
    CascadeMux I__1894 (
            .O(N__9085),
            .I(N__9079));
    CascadeMux I__1893 (
            .O(N__9082),
            .I(N__9076));
    CascadeBuf I__1892 (
            .O(N__9079),
            .I(N__9073));
    CascadeBuf I__1891 (
            .O(N__9076),
            .I(N__9070));
    CascadeMux I__1890 (
            .O(N__9073),
            .I(N__9067));
    CascadeMux I__1889 (
            .O(N__9070),
            .I(N__9064));
    CascadeBuf I__1888 (
            .O(N__9067),
            .I(N__9061));
    CascadeBuf I__1887 (
            .O(N__9064),
            .I(N__9058));
    CascadeMux I__1886 (
            .O(N__9061),
            .I(N__9055));
    CascadeMux I__1885 (
            .O(N__9058),
            .I(N__9052));
    CascadeBuf I__1884 (
            .O(N__9055),
            .I(N__9049));
    CascadeBuf I__1883 (
            .O(N__9052),
            .I(N__9046));
    CascadeMux I__1882 (
            .O(N__9049),
            .I(N__9043));
    CascadeMux I__1881 (
            .O(N__9046),
            .I(N__9040));
    CascadeBuf I__1880 (
            .O(N__9043),
            .I(N__9037));
    CascadeBuf I__1879 (
            .O(N__9040),
            .I(N__9034));
    CascadeMux I__1878 (
            .O(N__9037),
            .I(N__9031));
    CascadeMux I__1877 (
            .O(N__9034),
            .I(N__9028));
    CascadeBuf I__1876 (
            .O(N__9031),
            .I(N__9025));
    InMux I__1875 (
            .O(N__9028),
            .I(N__9022));
    CascadeMux I__1874 (
            .O(N__9025),
            .I(N__9019));
    LocalMux I__1873 (
            .O(N__9022),
            .I(N__9016));
    CascadeBuf I__1872 (
            .O(N__9019),
            .I(N__9013));
    Span4Mux_s3_v I__1871 (
            .O(N__9016),
            .I(N__9010));
    CascadeMux I__1870 (
            .O(N__9013),
            .I(N__9007));
    Sp12to4 I__1869 (
            .O(N__9010),
            .I(N__9004));
    InMux I__1868 (
            .O(N__9007),
            .I(N__9001));
    Span12Mux_h I__1867 (
            .O(N__9004),
            .I(N__8998));
    LocalMux I__1866 (
            .O(N__9001),
            .I(N__8995));
    Span12Mux_h I__1865 (
            .O(N__8998),
            .I(N__8992));
    IoSpan4Mux I__1864 (
            .O(N__8995),
            .I(N__8989));
    Odrv12 I__1863 (
            .O(N__8992),
            .I(waddr_c_3));
    Odrv4 I__1862 (
            .O(N__8989),
            .I(waddr_c_3));
    CascadeMux I__1861 (
            .O(N__8984),
            .I(N__8981));
    CascadeBuf I__1860 (
            .O(N__8981),
            .I(N__8978));
    CascadeMux I__1859 (
            .O(N__8978),
            .I(N__8975));
    CascadeBuf I__1858 (
            .O(N__8975),
            .I(N__8972));
    CascadeMux I__1857 (
            .O(N__8972),
            .I(N__8969));
    CascadeBuf I__1856 (
            .O(N__8969),
            .I(N__8965));
    CascadeMux I__1855 (
            .O(N__8968),
            .I(N__8962));
    CascadeMux I__1854 (
            .O(N__8965),
            .I(N__8959));
    CascadeBuf I__1853 (
            .O(N__8962),
            .I(N__8956));
    CascadeBuf I__1852 (
            .O(N__8959),
            .I(N__8953));
    CascadeMux I__1851 (
            .O(N__8956),
            .I(N__8950));
    CascadeMux I__1850 (
            .O(N__8953),
            .I(N__8947));
    CascadeBuf I__1849 (
            .O(N__8950),
            .I(N__8944));
    CascadeBuf I__1848 (
            .O(N__8947),
            .I(N__8941));
    CascadeMux I__1847 (
            .O(N__8944),
            .I(N__8938));
    CascadeMux I__1846 (
            .O(N__8941),
            .I(N__8935));
    CascadeBuf I__1845 (
            .O(N__8938),
            .I(N__8932));
    CascadeBuf I__1844 (
            .O(N__8935),
            .I(N__8929));
    CascadeMux I__1843 (
            .O(N__8932),
            .I(N__8926));
    CascadeMux I__1842 (
            .O(N__8929),
            .I(N__8923));
    CascadeBuf I__1841 (
            .O(N__8926),
            .I(N__8920));
    CascadeBuf I__1840 (
            .O(N__8923),
            .I(N__8917));
    CascadeMux I__1839 (
            .O(N__8920),
            .I(N__8914));
    CascadeMux I__1838 (
            .O(N__8917),
            .I(N__8911));
    CascadeBuf I__1837 (
            .O(N__8914),
            .I(N__8908));
    CascadeBuf I__1836 (
            .O(N__8911),
            .I(N__8905));
    CascadeMux I__1835 (
            .O(N__8908),
            .I(N__8902));
    CascadeMux I__1834 (
            .O(N__8905),
            .I(N__8899));
    CascadeBuf I__1833 (
            .O(N__8902),
            .I(N__8896));
    CascadeBuf I__1832 (
            .O(N__8899),
            .I(N__8893));
    CascadeMux I__1831 (
            .O(N__8896),
            .I(N__8890));
    CascadeMux I__1830 (
            .O(N__8893),
            .I(N__8887));
    CascadeBuf I__1829 (
            .O(N__8890),
            .I(N__8884));
    CascadeBuf I__1828 (
            .O(N__8887),
            .I(N__8881));
    CascadeMux I__1827 (
            .O(N__8884),
            .I(N__8878));
    CascadeMux I__1826 (
            .O(N__8881),
            .I(N__8875));
    CascadeBuf I__1825 (
            .O(N__8878),
            .I(N__8872));
    CascadeBuf I__1824 (
            .O(N__8875),
            .I(N__8869));
    CascadeMux I__1823 (
            .O(N__8872),
            .I(N__8866));
    CascadeMux I__1822 (
            .O(N__8869),
            .I(N__8863));
    CascadeBuf I__1821 (
            .O(N__8866),
            .I(N__8860));
    CascadeBuf I__1820 (
            .O(N__8863),
            .I(N__8857));
    CascadeMux I__1819 (
            .O(N__8860),
            .I(N__8854));
    CascadeMux I__1818 (
            .O(N__8857),
            .I(N__8851));
    CascadeBuf I__1817 (
            .O(N__8854),
            .I(N__8848));
    CascadeBuf I__1816 (
            .O(N__8851),
            .I(N__8845));
    CascadeMux I__1815 (
            .O(N__8848),
            .I(N__8842));
    CascadeMux I__1814 (
            .O(N__8845),
            .I(N__8839));
    CascadeBuf I__1813 (
            .O(N__8842),
            .I(N__8836));
    CascadeBuf I__1812 (
            .O(N__8839),
            .I(N__8833));
    CascadeMux I__1811 (
            .O(N__8836),
            .I(N__8830));
    CascadeMux I__1810 (
            .O(N__8833),
            .I(N__8827));
    CascadeBuf I__1809 (
            .O(N__8830),
            .I(N__8824));
    CascadeBuf I__1808 (
            .O(N__8827),
            .I(N__8821));
    CascadeMux I__1807 (
            .O(N__8824),
            .I(N__8818));
    CascadeMux I__1806 (
            .O(N__8821),
            .I(N__8815));
    CascadeBuf I__1805 (
            .O(N__8818),
            .I(N__8812));
    InMux I__1804 (
            .O(N__8815),
            .I(N__8809));
    CascadeMux I__1803 (
            .O(N__8812),
            .I(N__8806));
    LocalMux I__1802 (
            .O(N__8809),
            .I(N__8803));
    CascadeBuf I__1801 (
            .O(N__8806),
            .I(N__8800));
    Span4Mux_s3_v I__1800 (
            .O(N__8803),
            .I(N__8797));
    CascadeMux I__1799 (
            .O(N__8800),
            .I(N__8794));
    Span4Mux_h I__1798 (
            .O(N__8797),
            .I(N__8791));
    CascadeBuf I__1797 (
            .O(N__8794),
            .I(N__8788));
    Sp12to4 I__1796 (
            .O(N__8791),
            .I(N__8785));
    CascadeMux I__1795 (
            .O(N__8788),
            .I(N__8782));
    Span12Mux_h I__1794 (
            .O(N__8785),
            .I(N__8779));
    InMux I__1793 (
            .O(N__8782),
            .I(N__8776));
    Odrv12 I__1792 (
            .O(N__8779),
            .I(waddr_c_6));
    LocalMux I__1791 (
            .O(N__8776),
            .I(waddr_c_6));
    ClkMux I__1790 (
            .O(N__8771),
            .I(N__8675));
    ClkMux I__1789 (
            .O(N__8770),
            .I(N__8675));
    ClkMux I__1788 (
            .O(N__8769),
            .I(N__8675));
    ClkMux I__1787 (
            .O(N__8768),
            .I(N__8675));
    ClkMux I__1786 (
            .O(N__8767),
            .I(N__8675));
    ClkMux I__1785 (
            .O(N__8766),
            .I(N__8675));
    ClkMux I__1784 (
            .O(N__8765),
            .I(N__8675));
    ClkMux I__1783 (
            .O(N__8764),
            .I(N__8675));
    ClkMux I__1782 (
            .O(N__8763),
            .I(N__8675));
    ClkMux I__1781 (
            .O(N__8762),
            .I(N__8675));
    ClkMux I__1780 (
            .O(N__8761),
            .I(N__8675));
    ClkMux I__1779 (
            .O(N__8760),
            .I(N__8675));
    ClkMux I__1778 (
            .O(N__8759),
            .I(N__8675));
    ClkMux I__1777 (
            .O(N__8758),
            .I(N__8675));
    ClkMux I__1776 (
            .O(N__8757),
            .I(N__8675));
    ClkMux I__1775 (
            .O(N__8756),
            .I(N__8675));
    ClkMux I__1774 (
            .O(N__8755),
            .I(N__8675));
    ClkMux I__1773 (
            .O(N__8754),
            .I(N__8675));
    ClkMux I__1772 (
            .O(N__8753),
            .I(N__8675));
    ClkMux I__1771 (
            .O(N__8752),
            .I(N__8675));
    ClkMux I__1770 (
            .O(N__8751),
            .I(N__8675));
    ClkMux I__1769 (
            .O(N__8750),
            .I(N__8675));
    ClkMux I__1768 (
            .O(N__8749),
            .I(N__8675));
    ClkMux I__1767 (
            .O(N__8748),
            .I(N__8675));
    ClkMux I__1766 (
            .O(N__8747),
            .I(N__8675));
    ClkMux I__1765 (
            .O(N__8746),
            .I(N__8675));
    ClkMux I__1764 (
            .O(N__8745),
            .I(N__8675));
    ClkMux I__1763 (
            .O(N__8744),
            .I(N__8675));
    ClkMux I__1762 (
            .O(N__8743),
            .I(N__8675));
    ClkMux I__1761 (
            .O(N__8742),
            .I(N__8675));
    ClkMux I__1760 (
            .O(N__8741),
            .I(N__8675));
    ClkMux I__1759 (
            .O(N__8740),
            .I(N__8675));
    GlobalMux I__1758 (
            .O(N__8675),
            .I(N__8672));
    gio2CtrlBuf I__1757 (
            .O(N__8672),
            .I(wclk_c_g));
    CascadeMux I__1756 (
            .O(N__8669),
            .I(N__8666));
    CascadeBuf I__1755 (
            .O(N__8666),
            .I(N__8663));
    CascadeMux I__1754 (
            .O(N__8663),
            .I(N__8659));
    CascadeMux I__1753 (
            .O(N__8662),
            .I(N__8656));
    CascadeBuf I__1752 (
            .O(N__8659),
            .I(N__8653));
    CascadeBuf I__1751 (
            .O(N__8656),
            .I(N__8650));
    CascadeMux I__1750 (
            .O(N__8653),
            .I(N__8647));
    CascadeMux I__1749 (
            .O(N__8650),
            .I(N__8644));
    CascadeBuf I__1748 (
            .O(N__8647),
            .I(N__8641));
    CascadeBuf I__1747 (
            .O(N__8644),
            .I(N__8638));
    CascadeMux I__1746 (
            .O(N__8641),
            .I(N__8635));
    CascadeMux I__1745 (
            .O(N__8638),
            .I(N__8632));
    CascadeBuf I__1744 (
            .O(N__8635),
            .I(N__8629));
    CascadeBuf I__1743 (
            .O(N__8632),
            .I(N__8626));
    CascadeMux I__1742 (
            .O(N__8629),
            .I(N__8623));
    CascadeMux I__1741 (
            .O(N__8626),
            .I(N__8620));
    CascadeBuf I__1740 (
            .O(N__8623),
            .I(N__8617));
    CascadeBuf I__1739 (
            .O(N__8620),
            .I(N__8614));
    CascadeMux I__1738 (
            .O(N__8617),
            .I(N__8611));
    CascadeMux I__1737 (
            .O(N__8614),
            .I(N__8608));
    CascadeBuf I__1736 (
            .O(N__8611),
            .I(N__8605));
    CascadeBuf I__1735 (
            .O(N__8608),
            .I(N__8602));
    CascadeMux I__1734 (
            .O(N__8605),
            .I(N__8599));
    CascadeMux I__1733 (
            .O(N__8602),
            .I(N__8596));
    CascadeBuf I__1732 (
            .O(N__8599),
            .I(N__8593));
    CascadeBuf I__1731 (
            .O(N__8596),
            .I(N__8590));
    CascadeMux I__1730 (
            .O(N__8593),
            .I(N__8587));
    CascadeMux I__1729 (
            .O(N__8590),
            .I(N__8584));
    CascadeBuf I__1728 (
            .O(N__8587),
            .I(N__8581));
    CascadeBuf I__1727 (
            .O(N__8584),
            .I(N__8578));
    CascadeMux I__1726 (
            .O(N__8581),
            .I(N__8575));
    CascadeMux I__1725 (
            .O(N__8578),
            .I(N__8572));
    CascadeBuf I__1724 (
            .O(N__8575),
            .I(N__8569));
    CascadeBuf I__1723 (
            .O(N__8572),
            .I(N__8566));
    CascadeMux I__1722 (
            .O(N__8569),
            .I(N__8563));
    CascadeMux I__1721 (
            .O(N__8566),
            .I(N__8560));
    CascadeBuf I__1720 (
            .O(N__8563),
            .I(N__8557));
    CascadeBuf I__1719 (
            .O(N__8560),
            .I(N__8554));
    CascadeMux I__1718 (
            .O(N__8557),
            .I(N__8551));
    CascadeMux I__1717 (
            .O(N__8554),
            .I(N__8548));
    CascadeBuf I__1716 (
            .O(N__8551),
            .I(N__8545));
    CascadeBuf I__1715 (
            .O(N__8548),
            .I(N__8542));
    CascadeMux I__1714 (
            .O(N__8545),
            .I(N__8539));
    CascadeMux I__1713 (
            .O(N__8542),
            .I(N__8536));
    CascadeBuf I__1712 (
            .O(N__8539),
            .I(N__8533));
    CascadeBuf I__1711 (
            .O(N__8536),
            .I(N__8530));
    CascadeMux I__1710 (
            .O(N__8533),
            .I(N__8527));
    CascadeMux I__1709 (
            .O(N__8530),
            .I(N__8524));
    CascadeBuf I__1708 (
            .O(N__8527),
            .I(N__8521));
    CascadeBuf I__1707 (
            .O(N__8524),
            .I(N__8518));
    CascadeMux I__1706 (
            .O(N__8521),
            .I(N__8515));
    CascadeMux I__1705 (
            .O(N__8518),
            .I(N__8512));
    CascadeBuf I__1704 (
            .O(N__8515),
            .I(N__8509));
    CascadeBuf I__1703 (
            .O(N__8512),
            .I(N__8506));
    CascadeMux I__1702 (
            .O(N__8509),
            .I(N__8503));
    CascadeMux I__1701 (
            .O(N__8506),
            .I(N__8500));
    CascadeBuf I__1700 (
            .O(N__8503),
            .I(N__8497));
    CascadeBuf I__1699 (
            .O(N__8500),
            .I(N__8494));
    CascadeMux I__1698 (
            .O(N__8497),
            .I(N__8491));
    CascadeMux I__1697 (
            .O(N__8494),
            .I(N__8488));
    InMux I__1696 (
            .O(N__8491),
            .I(N__8485));
    CascadeBuf I__1695 (
            .O(N__8488),
            .I(N__8482));
    LocalMux I__1694 (
            .O(N__8485),
            .I(N__8479));
    CascadeMux I__1693 (
            .O(N__8482),
            .I(N__8476));
    Span4Mux_h I__1692 (
            .O(N__8479),
            .I(N__8473));
    InMux I__1691 (
            .O(N__8476),
            .I(N__8470));
    Span4Mux_h I__1690 (
            .O(N__8473),
            .I(N__8467));
    LocalMux I__1689 (
            .O(N__8470),
            .I(N__8464));
    Sp12to4 I__1688 (
            .O(N__8467),
            .I(N__8461));
    Span4Mux_h I__1687 (
            .O(N__8464),
            .I(N__8458));
    Span12Mux_s11_v I__1686 (
            .O(N__8461),
            .I(N__8455));
    Sp12to4 I__1685 (
            .O(N__8458),
            .I(N__8452));
    Span12Mux_h I__1684 (
            .O(N__8455),
            .I(N__8447));
    Span12Mux_s11_v I__1683 (
            .O(N__8452),
            .I(N__8447));
    Odrv12 I__1682 (
            .O(N__8447),
            .I(raddr_c_2));
    CascadeMux I__1681 (
            .O(N__8444),
            .I(N__8441));
    CascadeBuf I__1680 (
            .O(N__8441),
            .I(N__8438));
    CascadeMux I__1679 (
            .O(N__8438),
            .I(N__8434));
    CascadeMux I__1678 (
            .O(N__8437),
            .I(N__8431));
    CascadeBuf I__1677 (
            .O(N__8434),
            .I(N__8428));
    CascadeBuf I__1676 (
            .O(N__8431),
            .I(N__8425));
    CascadeMux I__1675 (
            .O(N__8428),
            .I(N__8422));
    CascadeMux I__1674 (
            .O(N__8425),
            .I(N__8419));
    CascadeBuf I__1673 (
            .O(N__8422),
            .I(N__8416));
    CascadeBuf I__1672 (
            .O(N__8419),
            .I(N__8413));
    CascadeMux I__1671 (
            .O(N__8416),
            .I(N__8410));
    CascadeMux I__1670 (
            .O(N__8413),
            .I(N__8407));
    CascadeBuf I__1669 (
            .O(N__8410),
            .I(N__8404));
    CascadeBuf I__1668 (
            .O(N__8407),
            .I(N__8401));
    CascadeMux I__1667 (
            .O(N__8404),
            .I(N__8398));
    CascadeMux I__1666 (
            .O(N__8401),
            .I(N__8395));
    CascadeBuf I__1665 (
            .O(N__8398),
            .I(N__8392));
    CascadeBuf I__1664 (
            .O(N__8395),
            .I(N__8389));
    CascadeMux I__1663 (
            .O(N__8392),
            .I(N__8386));
    CascadeMux I__1662 (
            .O(N__8389),
            .I(N__8383));
    CascadeBuf I__1661 (
            .O(N__8386),
            .I(N__8380));
    CascadeBuf I__1660 (
            .O(N__8383),
            .I(N__8377));
    CascadeMux I__1659 (
            .O(N__8380),
            .I(N__8374));
    CascadeMux I__1658 (
            .O(N__8377),
            .I(N__8371));
    CascadeBuf I__1657 (
            .O(N__8374),
            .I(N__8368));
    CascadeBuf I__1656 (
            .O(N__8371),
            .I(N__8365));
    CascadeMux I__1655 (
            .O(N__8368),
            .I(N__8362));
    CascadeMux I__1654 (
            .O(N__8365),
            .I(N__8359));
    CascadeBuf I__1653 (
            .O(N__8362),
            .I(N__8356));
    CascadeBuf I__1652 (
            .O(N__8359),
            .I(N__8353));
    CascadeMux I__1651 (
            .O(N__8356),
            .I(N__8350));
    CascadeMux I__1650 (
            .O(N__8353),
            .I(N__8347));
    CascadeBuf I__1649 (
            .O(N__8350),
            .I(N__8344));
    CascadeBuf I__1648 (
            .O(N__8347),
            .I(N__8341));
    CascadeMux I__1647 (
            .O(N__8344),
            .I(N__8338));
    CascadeMux I__1646 (
            .O(N__8341),
            .I(N__8335));
    CascadeBuf I__1645 (
            .O(N__8338),
            .I(N__8332));
    CascadeBuf I__1644 (
            .O(N__8335),
            .I(N__8329));
    CascadeMux I__1643 (
            .O(N__8332),
            .I(N__8326));
    CascadeMux I__1642 (
            .O(N__8329),
            .I(N__8323));
    CascadeBuf I__1641 (
            .O(N__8326),
            .I(N__8320));
    CascadeBuf I__1640 (
            .O(N__8323),
            .I(N__8317));
    CascadeMux I__1639 (
            .O(N__8320),
            .I(N__8314));
    CascadeMux I__1638 (
            .O(N__8317),
            .I(N__8311));
    CascadeBuf I__1637 (
            .O(N__8314),
            .I(N__8308));
    CascadeBuf I__1636 (
            .O(N__8311),
            .I(N__8305));
    CascadeMux I__1635 (
            .O(N__8308),
            .I(N__8302));
    CascadeMux I__1634 (
            .O(N__8305),
            .I(N__8299));
    CascadeBuf I__1633 (
            .O(N__8302),
            .I(N__8296));
    CascadeBuf I__1632 (
            .O(N__8299),
            .I(N__8293));
    CascadeMux I__1631 (
            .O(N__8296),
            .I(N__8290));
    CascadeMux I__1630 (
            .O(N__8293),
            .I(N__8287));
    CascadeBuf I__1629 (
            .O(N__8290),
            .I(N__8284));
    CascadeBuf I__1628 (
            .O(N__8287),
            .I(N__8281));
    CascadeMux I__1627 (
            .O(N__8284),
            .I(N__8278));
    CascadeMux I__1626 (
            .O(N__8281),
            .I(N__8275));
    CascadeBuf I__1625 (
            .O(N__8278),
            .I(N__8272));
    CascadeBuf I__1624 (
            .O(N__8275),
            .I(N__8269));
    CascadeMux I__1623 (
            .O(N__8272),
            .I(N__8266));
    CascadeMux I__1622 (
            .O(N__8269),
            .I(N__8263));
    InMux I__1621 (
            .O(N__8266),
            .I(N__8260));
    CascadeBuf I__1620 (
            .O(N__8263),
            .I(N__8257));
    LocalMux I__1619 (
            .O(N__8260),
            .I(N__8254));
    CascadeMux I__1618 (
            .O(N__8257),
            .I(N__8251));
    Span4Mux_v I__1617 (
            .O(N__8254),
            .I(N__8248));
    InMux I__1616 (
            .O(N__8251),
            .I(N__8245));
    Sp12to4 I__1615 (
            .O(N__8248),
            .I(N__8242));
    LocalMux I__1614 (
            .O(N__8245),
            .I(N__8239));
    Span12Mux_h I__1613 (
            .O(N__8242),
            .I(N__8236));
    Span12Mux_s5_v I__1612 (
            .O(N__8239),
            .I(N__8233));
    Odrv12 I__1611 (
            .O(N__8236),
            .I(raddr_c_7));
    Odrv12 I__1610 (
            .O(N__8233),
            .I(raddr_c_7));
    CascadeMux I__1609 (
            .O(N__8228),
            .I(N__8225));
    CascadeBuf I__1608 (
            .O(N__8225),
            .I(N__8222));
    CascadeMux I__1607 (
            .O(N__8222),
            .I(N__8219));
    CascadeBuf I__1606 (
            .O(N__8219),
            .I(N__8216));
    CascadeMux I__1605 (
            .O(N__8216),
            .I(N__8213));
    CascadeBuf I__1604 (
            .O(N__8213),
            .I(N__8209));
    CascadeMux I__1603 (
            .O(N__8212),
            .I(N__8206));
    CascadeMux I__1602 (
            .O(N__8209),
            .I(N__8203));
    CascadeBuf I__1601 (
            .O(N__8206),
            .I(N__8200));
    CascadeBuf I__1600 (
            .O(N__8203),
            .I(N__8197));
    CascadeMux I__1599 (
            .O(N__8200),
            .I(N__8194));
    CascadeMux I__1598 (
            .O(N__8197),
            .I(N__8191));
    CascadeBuf I__1597 (
            .O(N__8194),
            .I(N__8188));
    CascadeBuf I__1596 (
            .O(N__8191),
            .I(N__8185));
    CascadeMux I__1595 (
            .O(N__8188),
            .I(N__8182));
    CascadeMux I__1594 (
            .O(N__8185),
            .I(N__8179));
    CascadeBuf I__1593 (
            .O(N__8182),
            .I(N__8176));
    CascadeBuf I__1592 (
            .O(N__8179),
            .I(N__8173));
    CascadeMux I__1591 (
            .O(N__8176),
            .I(N__8170));
    CascadeMux I__1590 (
            .O(N__8173),
            .I(N__8167));
    CascadeBuf I__1589 (
            .O(N__8170),
            .I(N__8164));
    CascadeBuf I__1588 (
            .O(N__8167),
            .I(N__8161));
    CascadeMux I__1587 (
            .O(N__8164),
            .I(N__8158));
    CascadeMux I__1586 (
            .O(N__8161),
            .I(N__8155));
    CascadeBuf I__1585 (
            .O(N__8158),
            .I(N__8152));
    CascadeBuf I__1584 (
            .O(N__8155),
            .I(N__8149));
    CascadeMux I__1583 (
            .O(N__8152),
            .I(N__8146));
    CascadeMux I__1582 (
            .O(N__8149),
            .I(N__8143));
    CascadeBuf I__1581 (
            .O(N__8146),
            .I(N__8140));
    CascadeBuf I__1580 (
            .O(N__8143),
            .I(N__8137));
    CascadeMux I__1579 (
            .O(N__8140),
            .I(N__8134));
    CascadeMux I__1578 (
            .O(N__8137),
            .I(N__8131));
    CascadeBuf I__1577 (
            .O(N__8134),
            .I(N__8128));
    CascadeBuf I__1576 (
            .O(N__8131),
            .I(N__8125));
    CascadeMux I__1575 (
            .O(N__8128),
            .I(N__8122));
    CascadeMux I__1574 (
            .O(N__8125),
            .I(N__8119));
    CascadeBuf I__1573 (
            .O(N__8122),
            .I(N__8116));
    CascadeBuf I__1572 (
            .O(N__8119),
            .I(N__8113));
    CascadeMux I__1571 (
            .O(N__8116),
            .I(N__8110));
    CascadeMux I__1570 (
            .O(N__8113),
            .I(N__8107));
    CascadeBuf I__1569 (
            .O(N__8110),
            .I(N__8104));
    CascadeBuf I__1568 (
            .O(N__8107),
            .I(N__8101));
    CascadeMux I__1567 (
            .O(N__8104),
            .I(N__8098));
    CascadeMux I__1566 (
            .O(N__8101),
            .I(N__8095));
    CascadeBuf I__1565 (
            .O(N__8098),
            .I(N__8092));
    CascadeBuf I__1564 (
            .O(N__8095),
            .I(N__8089));
    CascadeMux I__1563 (
            .O(N__8092),
            .I(N__8086));
    CascadeMux I__1562 (
            .O(N__8089),
            .I(N__8083));
    CascadeBuf I__1561 (
            .O(N__8086),
            .I(N__8080));
    CascadeBuf I__1560 (
            .O(N__8083),
            .I(N__8077));
    CascadeMux I__1559 (
            .O(N__8080),
            .I(N__8074));
    CascadeMux I__1558 (
            .O(N__8077),
            .I(N__8071));
    CascadeBuf I__1557 (
            .O(N__8074),
            .I(N__8068));
    CascadeBuf I__1556 (
            .O(N__8071),
            .I(N__8065));
    CascadeMux I__1555 (
            .O(N__8068),
            .I(N__8062));
    CascadeMux I__1554 (
            .O(N__8065),
            .I(N__8059));
    CascadeBuf I__1553 (
            .O(N__8062),
            .I(N__8056));
    InMux I__1552 (
            .O(N__8059),
            .I(N__8053));
    CascadeMux I__1551 (
            .O(N__8056),
            .I(N__8050));
    LocalMux I__1550 (
            .O(N__8053),
            .I(N__8047));
    CascadeBuf I__1549 (
            .O(N__8050),
            .I(N__8044));
    Span4Mux_s1_v I__1548 (
            .O(N__8047),
            .I(N__8041));
    CascadeMux I__1547 (
            .O(N__8044),
            .I(N__8038));
    Span4Mux_h I__1546 (
            .O(N__8041),
            .I(N__8035));
    CascadeBuf I__1545 (
            .O(N__8038),
            .I(N__8032));
    Sp12to4 I__1544 (
            .O(N__8035),
            .I(N__8029));
    CascadeMux I__1543 (
            .O(N__8032),
            .I(N__8026));
    Span12Mux_h I__1542 (
            .O(N__8029),
            .I(N__8023));
    InMux I__1541 (
            .O(N__8026),
            .I(N__8020));
    Odrv12 I__1540 (
            .O(N__8023),
            .I(waddr_c_5));
    LocalMux I__1539 (
            .O(N__8020),
            .I(waddr_c_5));
    InMux I__1538 (
            .O(N__8015),
            .I(N__8009));
    InMux I__1537 (
            .O(N__8014),
            .I(N__8006));
    InMux I__1536 (
            .O(N__8013),
            .I(N__7999));
    InMux I__1535 (
            .O(N__8012),
            .I(N__7996));
    LocalMux I__1534 (
            .O(N__8009),
            .I(N__7993));
    LocalMux I__1533 (
            .O(N__8006),
            .I(N__7990));
    InMux I__1532 (
            .O(N__8005),
            .I(N__7987));
    InMux I__1531 (
            .O(N__8004),
            .I(N__7984));
    InMux I__1530 (
            .O(N__8003),
            .I(N__7981));
    InMux I__1529 (
            .O(N__8002),
            .I(N__7978));
    LocalMux I__1528 (
            .O(N__7999),
            .I(N__7975));
    LocalMux I__1527 (
            .O(N__7996),
            .I(N__7972));
    Span12Mux_h I__1526 (
            .O(N__7993),
            .I(N__7967));
    Span12Mux_h I__1525 (
            .O(N__7990),
            .I(N__7967));
    LocalMux I__1524 (
            .O(N__7987),
            .I(N__7964));
    LocalMux I__1523 (
            .O(N__7984),
            .I(N__7961));
    LocalMux I__1522 (
            .O(N__7981),
            .I(N__7958));
    LocalMux I__1521 (
            .O(N__7978),
            .I(N__7955));
    Span4Mux_v I__1520 (
            .O(N__7975),
            .I(N__7952));
    Span4Mux_v I__1519 (
            .O(N__7972),
            .I(N__7949));
    Span12Mux_v I__1518 (
            .O(N__7967),
            .I(N__7946));
    Span12Mux_h I__1517 (
            .O(N__7964),
            .I(N__7941));
    Span12Mux_h I__1516 (
            .O(N__7961),
            .I(N__7941));
    Span12Mux_h I__1515 (
            .O(N__7958),
            .I(N__7936));
    Span12Mux_h I__1514 (
            .O(N__7955),
            .I(N__7936));
    Sp12to4 I__1513 (
            .O(N__7952),
            .I(N__7933));
    Sp12to4 I__1512 (
            .O(N__7949),
            .I(N__7930));
    Span12Mux_v I__1511 (
            .O(N__7946),
            .I(N__7927));
    Span12Mux_v I__1510 (
            .O(N__7941),
            .I(N__7924));
    Span12Mux_v I__1509 (
            .O(N__7936),
            .I(N__7917));
    Span12Mux_h I__1508 (
            .O(N__7933),
            .I(N__7917));
    Span12Mux_h I__1507 (
            .O(N__7930),
            .I(N__7917));
    Odrv12 I__1506 (
            .O(N__7927),
            .I(din_c_1));
    Odrv12 I__1505 (
            .O(N__7924),
            .I(din_c_1));
    Odrv12 I__1504 (
            .O(N__7917),
            .I(din_c_1));
    CascadeMux I__1503 (
            .O(N__7910),
            .I(N__7907));
    CascadeBuf I__1502 (
            .O(N__7907),
            .I(N__7904));
    CascadeMux I__1501 (
            .O(N__7904),
            .I(N__7900));
    CascadeMux I__1500 (
            .O(N__7903),
            .I(N__7897));
    CascadeBuf I__1499 (
            .O(N__7900),
            .I(N__7894));
    CascadeBuf I__1498 (
            .O(N__7897),
            .I(N__7891));
    CascadeMux I__1497 (
            .O(N__7894),
            .I(N__7888));
    CascadeMux I__1496 (
            .O(N__7891),
            .I(N__7885));
    CascadeBuf I__1495 (
            .O(N__7888),
            .I(N__7882));
    CascadeBuf I__1494 (
            .O(N__7885),
            .I(N__7879));
    CascadeMux I__1493 (
            .O(N__7882),
            .I(N__7876));
    CascadeMux I__1492 (
            .O(N__7879),
            .I(N__7873));
    CascadeBuf I__1491 (
            .O(N__7876),
            .I(N__7870));
    CascadeBuf I__1490 (
            .O(N__7873),
            .I(N__7867));
    CascadeMux I__1489 (
            .O(N__7870),
            .I(N__7864));
    CascadeMux I__1488 (
            .O(N__7867),
            .I(N__7861));
    CascadeBuf I__1487 (
            .O(N__7864),
            .I(N__7858));
    CascadeBuf I__1486 (
            .O(N__7861),
            .I(N__7855));
    CascadeMux I__1485 (
            .O(N__7858),
            .I(N__7852));
    CascadeMux I__1484 (
            .O(N__7855),
            .I(N__7849));
    CascadeBuf I__1483 (
            .O(N__7852),
            .I(N__7846));
    CascadeBuf I__1482 (
            .O(N__7849),
            .I(N__7843));
    CascadeMux I__1481 (
            .O(N__7846),
            .I(N__7840));
    CascadeMux I__1480 (
            .O(N__7843),
            .I(N__7837));
    CascadeBuf I__1479 (
            .O(N__7840),
            .I(N__7834));
    CascadeBuf I__1478 (
            .O(N__7837),
            .I(N__7831));
    CascadeMux I__1477 (
            .O(N__7834),
            .I(N__7828));
    CascadeMux I__1476 (
            .O(N__7831),
            .I(N__7825));
    CascadeBuf I__1475 (
            .O(N__7828),
            .I(N__7822));
    CascadeBuf I__1474 (
            .O(N__7825),
            .I(N__7819));
    CascadeMux I__1473 (
            .O(N__7822),
            .I(N__7816));
    CascadeMux I__1472 (
            .O(N__7819),
            .I(N__7813));
    CascadeBuf I__1471 (
            .O(N__7816),
            .I(N__7810));
    CascadeBuf I__1470 (
            .O(N__7813),
            .I(N__7807));
    CascadeMux I__1469 (
            .O(N__7810),
            .I(N__7804));
    CascadeMux I__1468 (
            .O(N__7807),
            .I(N__7801));
    CascadeBuf I__1467 (
            .O(N__7804),
            .I(N__7798));
    CascadeBuf I__1466 (
            .O(N__7801),
            .I(N__7795));
    CascadeMux I__1465 (
            .O(N__7798),
            .I(N__7792));
    CascadeMux I__1464 (
            .O(N__7795),
            .I(N__7789));
    CascadeBuf I__1463 (
            .O(N__7792),
            .I(N__7786));
    CascadeBuf I__1462 (
            .O(N__7789),
            .I(N__7783));
    CascadeMux I__1461 (
            .O(N__7786),
            .I(N__7780));
    CascadeMux I__1460 (
            .O(N__7783),
            .I(N__7777));
    CascadeBuf I__1459 (
            .O(N__7780),
            .I(N__7774));
    CascadeBuf I__1458 (
            .O(N__7777),
            .I(N__7771));
    CascadeMux I__1457 (
            .O(N__7774),
            .I(N__7768));
    CascadeMux I__1456 (
            .O(N__7771),
            .I(N__7765));
    CascadeBuf I__1455 (
            .O(N__7768),
            .I(N__7762));
    CascadeBuf I__1454 (
            .O(N__7765),
            .I(N__7759));
    CascadeMux I__1453 (
            .O(N__7762),
            .I(N__7756));
    CascadeMux I__1452 (
            .O(N__7759),
            .I(N__7753));
    CascadeBuf I__1451 (
            .O(N__7756),
            .I(N__7750));
    CascadeBuf I__1450 (
            .O(N__7753),
            .I(N__7747));
    CascadeMux I__1449 (
            .O(N__7750),
            .I(N__7744));
    CascadeMux I__1448 (
            .O(N__7747),
            .I(N__7741));
    CascadeBuf I__1447 (
            .O(N__7744),
            .I(N__7738));
    CascadeBuf I__1446 (
            .O(N__7741),
            .I(N__7735));
    CascadeMux I__1445 (
            .O(N__7738),
            .I(N__7732));
    CascadeMux I__1444 (
            .O(N__7735),
            .I(N__7729));
    InMux I__1443 (
            .O(N__7732),
            .I(N__7726));
    CascadeBuf I__1442 (
            .O(N__7729),
            .I(N__7723));
    LocalMux I__1441 (
            .O(N__7726),
            .I(N__7720));
    CascadeMux I__1440 (
            .O(N__7723),
            .I(N__7717));
    Span4Mux_v I__1439 (
            .O(N__7720),
            .I(N__7714));
    InMux I__1438 (
            .O(N__7717),
            .I(N__7711));
    Span4Mux_h I__1437 (
            .O(N__7714),
            .I(N__7708));
    LocalMux I__1436 (
            .O(N__7711),
            .I(N__7705));
    Sp12to4 I__1435 (
            .O(N__7708),
            .I(N__7702));
    Span4Mux_v I__1434 (
            .O(N__7705),
            .I(N__7699));
    Span12Mux_h I__1433 (
            .O(N__7702),
            .I(N__7694));
    Sp12to4 I__1432 (
            .O(N__7699),
            .I(N__7694));
    Odrv12 I__1431 (
            .O(N__7694),
            .I(raddr_c_8));
    CascadeMux I__1430 (
            .O(N__7691),
            .I(N__7688));
    CascadeBuf I__1429 (
            .O(N__7688),
            .I(N__7685));
    CascadeMux I__1428 (
            .O(N__7685),
            .I(N__7682));
    CascadeBuf I__1427 (
            .O(N__7682),
            .I(N__7678));
    CascadeMux I__1426 (
            .O(N__7681),
            .I(N__7675));
    CascadeMux I__1425 (
            .O(N__7678),
            .I(N__7672));
    CascadeBuf I__1424 (
            .O(N__7675),
            .I(N__7669));
    CascadeBuf I__1423 (
            .O(N__7672),
            .I(N__7666));
    CascadeMux I__1422 (
            .O(N__7669),
            .I(N__7663));
    CascadeMux I__1421 (
            .O(N__7666),
            .I(N__7660));
    CascadeBuf I__1420 (
            .O(N__7663),
            .I(N__7657));
    CascadeBuf I__1419 (
            .O(N__7660),
            .I(N__7654));
    CascadeMux I__1418 (
            .O(N__7657),
            .I(N__7651));
    CascadeMux I__1417 (
            .O(N__7654),
            .I(N__7648));
    CascadeBuf I__1416 (
            .O(N__7651),
            .I(N__7645));
    CascadeBuf I__1415 (
            .O(N__7648),
            .I(N__7642));
    CascadeMux I__1414 (
            .O(N__7645),
            .I(N__7639));
    CascadeMux I__1413 (
            .O(N__7642),
            .I(N__7636));
    CascadeBuf I__1412 (
            .O(N__7639),
            .I(N__7633));
    CascadeBuf I__1411 (
            .O(N__7636),
            .I(N__7630));
    CascadeMux I__1410 (
            .O(N__7633),
            .I(N__7627));
    CascadeMux I__1409 (
            .O(N__7630),
            .I(N__7624));
    CascadeBuf I__1408 (
            .O(N__7627),
            .I(N__7621));
    CascadeBuf I__1407 (
            .O(N__7624),
            .I(N__7618));
    CascadeMux I__1406 (
            .O(N__7621),
            .I(N__7615));
    CascadeMux I__1405 (
            .O(N__7618),
            .I(N__7612));
    CascadeBuf I__1404 (
            .O(N__7615),
            .I(N__7609));
    CascadeBuf I__1403 (
            .O(N__7612),
            .I(N__7606));
    CascadeMux I__1402 (
            .O(N__7609),
            .I(N__7603));
    CascadeMux I__1401 (
            .O(N__7606),
            .I(N__7600));
    CascadeBuf I__1400 (
            .O(N__7603),
            .I(N__7597));
    CascadeBuf I__1399 (
            .O(N__7600),
            .I(N__7594));
    CascadeMux I__1398 (
            .O(N__7597),
            .I(N__7591));
    CascadeMux I__1397 (
            .O(N__7594),
            .I(N__7588));
    CascadeBuf I__1396 (
            .O(N__7591),
            .I(N__7585));
    CascadeBuf I__1395 (
            .O(N__7588),
            .I(N__7582));
    CascadeMux I__1394 (
            .O(N__7585),
            .I(N__7579));
    CascadeMux I__1393 (
            .O(N__7582),
            .I(N__7576));
    CascadeBuf I__1392 (
            .O(N__7579),
            .I(N__7573));
    CascadeBuf I__1391 (
            .O(N__7576),
            .I(N__7570));
    CascadeMux I__1390 (
            .O(N__7573),
            .I(N__7567));
    CascadeMux I__1389 (
            .O(N__7570),
            .I(N__7564));
    CascadeBuf I__1388 (
            .O(N__7567),
            .I(N__7561));
    CascadeBuf I__1387 (
            .O(N__7564),
            .I(N__7558));
    CascadeMux I__1386 (
            .O(N__7561),
            .I(N__7555));
    CascadeMux I__1385 (
            .O(N__7558),
            .I(N__7552));
    CascadeBuf I__1384 (
            .O(N__7555),
            .I(N__7549));
    CascadeBuf I__1383 (
            .O(N__7552),
            .I(N__7546));
    CascadeMux I__1382 (
            .O(N__7549),
            .I(N__7543));
    CascadeMux I__1381 (
            .O(N__7546),
            .I(N__7540));
    CascadeBuf I__1380 (
            .O(N__7543),
            .I(N__7537));
    CascadeBuf I__1379 (
            .O(N__7540),
            .I(N__7534));
    CascadeMux I__1378 (
            .O(N__7537),
            .I(N__7531));
    CascadeMux I__1377 (
            .O(N__7534),
            .I(N__7528));
    CascadeBuf I__1376 (
            .O(N__7531),
            .I(N__7525));
    CascadeBuf I__1375 (
            .O(N__7528),
            .I(N__7522));
    CascadeMux I__1374 (
            .O(N__7525),
            .I(N__7519));
    CascadeMux I__1373 (
            .O(N__7522),
            .I(N__7516));
    CascadeBuf I__1372 (
            .O(N__7519),
            .I(N__7513));
    InMux I__1371 (
            .O(N__7516),
            .I(N__7510));
    CascadeMux I__1370 (
            .O(N__7513),
            .I(N__7507));
    LocalMux I__1369 (
            .O(N__7510),
            .I(N__7504));
    CascadeBuf I__1368 (
            .O(N__7507),
            .I(N__7501));
    Span4Mux_s3_v I__1367 (
            .O(N__7504),
            .I(N__7498));
    CascadeMux I__1366 (
            .O(N__7501),
            .I(N__7495));
    Sp12to4 I__1365 (
            .O(N__7498),
            .I(N__7492));
    InMux I__1364 (
            .O(N__7495),
            .I(N__7489));
    Span12Mux_h I__1363 (
            .O(N__7492),
            .I(N__7486));
    LocalMux I__1362 (
            .O(N__7489),
            .I(N__7483));
    Span12Mux_h I__1361 (
            .O(N__7486),
            .I(N__7480));
    Span4Mux_h I__1360 (
            .O(N__7483),
            .I(N__7477));
    Odrv12 I__1359 (
            .O(N__7480),
            .I(waddr_c_4));
    Odrv4 I__1358 (
            .O(N__7477),
            .I(waddr_c_4));
    CascadeMux I__1357 (
            .O(N__7472),
            .I(N__7469));
    CascadeBuf I__1356 (
            .O(N__7469),
            .I(N__7466));
    CascadeMux I__1355 (
            .O(N__7466),
            .I(N__7463));
    CascadeBuf I__1354 (
            .O(N__7463),
            .I(N__7459));
    CascadeMux I__1353 (
            .O(N__7462),
            .I(N__7456));
    CascadeMux I__1352 (
            .O(N__7459),
            .I(N__7453));
    CascadeBuf I__1351 (
            .O(N__7456),
            .I(N__7450));
    CascadeBuf I__1350 (
            .O(N__7453),
            .I(N__7447));
    CascadeMux I__1349 (
            .O(N__7450),
            .I(N__7444));
    CascadeMux I__1348 (
            .O(N__7447),
            .I(N__7441));
    CascadeBuf I__1347 (
            .O(N__7444),
            .I(N__7438));
    CascadeBuf I__1346 (
            .O(N__7441),
            .I(N__7435));
    CascadeMux I__1345 (
            .O(N__7438),
            .I(N__7432));
    CascadeMux I__1344 (
            .O(N__7435),
            .I(N__7429));
    CascadeBuf I__1343 (
            .O(N__7432),
            .I(N__7426));
    CascadeBuf I__1342 (
            .O(N__7429),
            .I(N__7423));
    CascadeMux I__1341 (
            .O(N__7426),
            .I(N__7420));
    CascadeMux I__1340 (
            .O(N__7423),
            .I(N__7417));
    CascadeBuf I__1339 (
            .O(N__7420),
            .I(N__7414));
    CascadeBuf I__1338 (
            .O(N__7417),
            .I(N__7411));
    CascadeMux I__1337 (
            .O(N__7414),
            .I(N__7408));
    CascadeMux I__1336 (
            .O(N__7411),
            .I(N__7405));
    CascadeBuf I__1335 (
            .O(N__7408),
            .I(N__7402));
    CascadeBuf I__1334 (
            .O(N__7405),
            .I(N__7399));
    CascadeMux I__1333 (
            .O(N__7402),
            .I(N__7396));
    CascadeMux I__1332 (
            .O(N__7399),
            .I(N__7393));
    CascadeBuf I__1331 (
            .O(N__7396),
            .I(N__7390));
    CascadeBuf I__1330 (
            .O(N__7393),
            .I(N__7387));
    CascadeMux I__1329 (
            .O(N__7390),
            .I(N__7384));
    CascadeMux I__1328 (
            .O(N__7387),
            .I(N__7381));
    CascadeBuf I__1327 (
            .O(N__7384),
            .I(N__7378));
    CascadeBuf I__1326 (
            .O(N__7381),
            .I(N__7375));
    CascadeMux I__1325 (
            .O(N__7378),
            .I(N__7372));
    CascadeMux I__1324 (
            .O(N__7375),
            .I(N__7369));
    CascadeBuf I__1323 (
            .O(N__7372),
            .I(N__7366));
    CascadeBuf I__1322 (
            .O(N__7369),
            .I(N__7363));
    CascadeMux I__1321 (
            .O(N__7366),
            .I(N__7360));
    CascadeMux I__1320 (
            .O(N__7363),
            .I(N__7357));
    CascadeBuf I__1319 (
            .O(N__7360),
            .I(N__7354));
    CascadeBuf I__1318 (
            .O(N__7357),
            .I(N__7351));
    CascadeMux I__1317 (
            .O(N__7354),
            .I(N__7348));
    CascadeMux I__1316 (
            .O(N__7351),
            .I(N__7345));
    CascadeBuf I__1315 (
            .O(N__7348),
            .I(N__7342));
    CascadeBuf I__1314 (
            .O(N__7345),
            .I(N__7339));
    CascadeMux I__1313 (
            .O(N__7342),
            .I(N__7336));
    CascadeMux I__1312 (
            .O(N__7339),
            .I(N__7333));
    CascadeBuf I__1311 (
            .O(N__7336),
            .I(N__7330));
    CascadeBuf I__1310 (
            .O(N__7333),
            .I(N__7327));
    CascadeMux I__1309 (
            .O(N__7330),
            .I(N__7324));
    CascadeMux I__1308 (
            .O(N__7327),
            .I(N__7321));
    CascadeBuf I__1307 (
            .O(N__7324),
            .I(N__7318));
    CascadeBuf I__1306 (
            .O(N__7321),
            .I(N__7315));
    CascadeMux I__1305 (
            .O(N__7318),
            .I(N__7312));
    CascadeMux I__1304 (
            .O(N__7315),
            .I(N__7309));
    CascadeBuf I__1303 (
            .O(N__7312),
            .I(N__7306));
    CascadeBuf I__1302 (
            .O(N__7309),
            .I(N__7303));
    CascadeMux I__1301 (
            .O(N__7306),
            .I(N__7300));
    CascadeMux I__1300 (
            .O(N__7303),
            .I(N__7297));
    CascadeBuf I__1299 (
            .O(N__7300),
            .I(N__7294));
    InMux I__1298 (
            .O(N__7297),
            .I(N__7291));
    CascadeMux I__1297 (
            .O(N__7294),
            .I(N__7288));
    LocalMux I__1296 (
            .O(N__7291),
            .I(N__7285));
    CascadeBuf I__1295 (
            .O(N__7288),
            .I(N__7282));
    Span4Mux_h I__1294 (
            .O(N__7285),
            .I(N__7279));
    CascadeMux I__1293 (
            .O(N__7282),
            .I(N__7276));
    Sp12to4 I__1292 (
            .O(N__7279),
            .I(N__7273));
    InMux I__1291 (
            .O(N__7276),
            .I(N__7270));
    Span12Mux_s11_v I__1290 (
            .O(N__7273),
            .I(N__7267));
    LocalMux I__1289 (
            .O(N__7270),
            .I(N__7264));
    Span12Mux_h I__1288 (
            .O(N__7267),
            .I(N__7261));
    Span12Mux_s11_v I__1287 (
            .O(N__7264),
            .I(N__7258));
    Odrv12 I__1286 (
            .O(N__7261),
            .I(raddr_c_10));
    Odrv12 I__1285 (
            .O(N__7258),
            .I(raddr_c_10));
    CascadeMux I__1284 (
            .O(N__7253),
            .I(N__7250));
    CascadeBuf I__1283 (
            .O(N__7250),
            .I(N__7246));
    CascadeMux I__1282 (
            .O(N__7249),
            .I(N__7243));
    CascadeMux I__1281 (
            .O(N__7246),
            .I(N__7240));
    CascadeBuf I__1280 (
            .O(N__7243),
            .I(N__7237));
    CascadeBuf I__1279 (
            .O(N__7240),
            .I(N__7234));
    CascadeMux I__1278 (
            .O(N__7237),
            .I(N__7231));
    CascadeMux I__1277 (
            .O(N__7234),
            .I(N__7228));
    CascadeBuf I__1276 (
            .O(N__7231),
            .I(N__7225));
    CascadeBuf I__1275 (
            .O(N__7228),
            .I(N__7222));
    CascadeMux I__1274 (
            .O(N__7225),
            .I(N__7219));
    CascadeMux I__1273 (
            .O(N__7222),
            .I(N__7216));
    CascadeBuf I__1272 (
            .O(N__7219),
            .I(N__7213));
    CascadeBuf I__1271 (
            .O(N__7216),
            .I(N__7210));
    CascadeMux I__1270 (
            .O(N__7213),
            .I(N__7207));
    CascadeMux I__1269 (
            .O(N__7210),
            .I(N__7204));
    CascadeBuf I__1268 (
            .O(N__7207),
            .I(N__7201));
    CascadeBuf I__1267 (
            .O(N__7204),
            .I(N__7198));
    CascadeMux I__1266 (
            .O(N__7201),
            .I(N__7195));
    CascadeMux I__1265 (
            .O(N__7198),
            .I(N__7192));
    CascadeBuf I__1264 (
            .O(N__7195),
            .I(N__7189));
    CascadeBuf I__1263 (
            .O(N__7192),
            .I(N__7186));
    CascadeMux I__1262 (
            .O(N__7189),
            .I(N__7183));
    CascadeMux I__1261 (
            .O(N__7186),
            .I(N__7180));
    CascadeBuf I__1260 (
            .O(N__7183),
            .I(N__7177));
    CascadeBuf I__1259 (
            .O(N__7180),
            .I(N__7174));
    CascadeMux I__1258 (
            .O(N__7177),
            .I(N__7171));
    CascadeMux I__1257 (
            .O(N__7174),
            .I(N__7168));
    CascadeBuf I__1256 (
            .O(N__7171),
            .I(N__7165));
    CascadeBuf I__1255 (
            .O(N__7168),
            .I(N__7162));
    CascadeMux I__1254 (
            .O(N__7165),
            .I(N__7159));
    CascadeMux I__1253 (
            .O(N__7162),
            .I(N__7156));
    CascadeBuf I__1252 (
            .O(N__7159),
            .I(N__7153));
    CascadeBuf I__1251 (
            .O(N__7156),
            .I(N__7150));
    CascadeMux I__1250 (
            .O(N__7153),
            .I(N__7147));
    CascadeMux I__1249 (
            .O(N__7150),
            .I(N__7144));
    CascadeBuf I__1248 (
            .O(N__7147),
            .I(N__7141));
    CascadeBuf I__1247 (
            .O(N__7144),
            .I(N__7138));
    CascadeMux I__1246 (
            .O(N__7141),
            .I(N__7135));
    CascadeMux I__1245 (
            .O(N__7138),
            .I(N__7132));
    CascadeBuf I__1244 (
            .O(N__7135),
            .I(N__7129));
    CascadeBuf I__1243 (
            .O(N__7132),
            .I(N__7126));
    CascadeMux I__1242 (
            .O(N__7129),
            .I(N__7123));
    CascadeMux I__1241 (
            .O(N__7126),
            .I(N__7120));
    CascadeBuf I__1240 (
            .O(N__7123),
            .I(N__7117));
    CascadeBuf I__1239 (
            .O(N__7120),
            .I(N__7114));
    CascadeMux I__1238 (
            .O(N__7117),
            .I(N__7111));
    CascadeMux I__1237 (
            .O(N__7114),
            .I(N__7108));
    CascadeBuf I__1236 (
            .O(N__7111),
            .I(N__7105));
    CascadeBuf I__1235 (
            .O(N__7108),
            .I(N__7102));
    CascadeMux I__1234 (
            .O(N__7105),
            .I(N__7099));
    CascadeMux I__1233 (
            .O(N__7102),
            .I(N__7096));
    CascadeBuf I__1232 (
            .O(N__7099),
            .I(N__7093));
    CascadeBuf I__1231 (
            .O(N__7096),
            .I(N__7090));
    CascadeMux I__1230 (
            .O(N__7093),
            .I(N__7087));
    CascadeMux I__1229 (
            .O(N__7090),
            .I(N__7084));
    CascadeBuf I__1228 (
            .O(N__7087),
            .I(N__7081));
    CascadeBuf I__1227 (
            .O(N__7084),
            .I(N__7078));
    CascadeMux I__1226 (
            .O(N__7081),
            .I(N__7075));
    CascadeMux I__1225 (
            .O(N__7078),
            .I(N__7072));
    CascadeBuf I__1224 (
            .O(N__7075),
            .I(N__7069));
    InMux I__1223 (
            .O(N__7072),
            .I(N__7066));
    CascadeMux I__1222 (
            .O(N__7069),
            .I(N__7063));
    LocalMux I__1221 (
            .O(N__7066),
            .I(N__7060));
    InMux I__1220 (
            .O(N__7063),
            .I(N__7057));
    Span4Mux_v I__1219 (
            .O(N__7060),
            .I(N__7054));
    LocalMux I__1218 (
            .O(N__7057),
            .I(N__7051));
    Span4Mux_h I__1217 (
            .O(N__7054),
            .I(N__7048));
    Span4Mux_s2_v I__1216 (
            .O(N__7051),
            .I(N__7045));
    Sp12to4 I__1215 (
            .O(N__7048),
            .I(N__7042));
    Span4Mux_v I__1214 (
            .O(N__7045),
            .I(N__7039));
    Span12Mux_s10_v I__1213 (
            .O(N__7042),
            .I(N__7036));
    Span4Mux_v I__1212 (
            .O(N__7039),
            .I(N__7033));
    Span12Mux_h I__1211 (
            .O(N__7036),
            .I(N__7028));
    Sp12to4 I__1210 (
            .O(N__7033),
            .I(N__7028));
    Odrv12 I__1209 (
            .O(N__7028),
            .I(raddr_c_4));
    CascadeMux I__1208 (
            .O(N__7025),
            .I(N__7022));
    CascadeBuf I__1207 (
            .O(N__7022),
            .I(N__7019));
    CascadeMux I__1206 (
            .O(N__7019),
            .I(N__7016));
    CascadeBuf I__1205 (
            .O(N__7016),
            .I(N__7012));
    CascadeMux I__1204 (
            .O(N__7015),
            .I(N__7009));
    CascadeMux I__1203 (
            .O(N__7012),
            .I(N__7006));
    CascadeBuf I__1202 (
            .O(N__7009),
            .I(N__7003));
    CascadeBuf I__1201 (
            .O(N__7006),
            .I(N__7000));
    CascadeMux I__1200 (
            .O(N__7003),
            .I(N__6997));
    CascadeMux I__1199 (
            .O(N__7000),
            .I(N__6994));
    CascadeBuf I__1198 (
            .O(N__6997),
            .I(N__6991));
    CascadeBuf I__1197 (
            .O(N__6994),
            .I(N__6988));
    CascadeMux I__1196 (
            .O(N__6991),
            .I(N__6985));
    CascadeMux I__1195 (
            .O(N__6988),
            .I(N__6982));
    CascadeBuf I__1194 (
            .O(N__6985),
            .I(N__6979));
    CascadeBuf I__1193 (
            .O(N__6982),
            .I(N__6976));
    CascadeMux I__1192 (
            .O(N__6979),
            .I(N__6973));
    CascadeMux I__1191 (
            .O(N__6976),
            .I(N__6970));
    CascadeBuf I__1190 (
            .O(N__6973),
            .I(N__6967));
    CascadeBuf I__1189 (
            .O(N__6970),
            .I(N__6964));
    CascadeMux I__1188 (
            .O(N__6967),
            .I(N__6961));
    CascadeMux I__1187 (
            .O(N__6964),
            .I(N__6958));
    CascadeBuf I__1186 (
            .O(N__6961),
            .I(N__6955));
    CascadeBuf I__1185 (
            .O(N__6958),
            .I(N__6952));
    CascadeMux I__1184 (
            .O(N__6955),
            .I(N__6949));
    CascadeMux I__1183 (
            .O(N__6952),
            .I(N__6946));
    CascadeBuf I__1182 (
            .O(N__6949),
            .I(N__6943));
    CascadeBuf I__1181 (
            .O(N__6946),
            .I(N__6940));
    CascadeMux I__1180 (
            .O(N__6943),
            .I(N__6937));
    CascadeMux I__1179 (
            .O(N__6940),
            .I(N__6934));
    CascadeBuf I__1178 (
            .O(N__6937),
            .I(N__6931));
    CascadeBuf I__1177 (
            .O(N__6934),
            .I(N__6928));
    CascadeMux I__1176 (
            .O(N__6931),
            .I(N__6925));
    CascadeMux I__1175 (
            .O(N__6928),
            .I(N__6922));
    CascadeBuf I__1174 (
            .O(N__6925),
            .I(N__6919));
    CascadeBuf I__1173 (
            .O(N__6922),
            .I(N__6916));
    CascadeMux I__1172 (
            .O(N__6919),
            .I(N__6913));
    CascadeMux I__1171 (
            .O(N__6916),
            .I(N__6910));
    CascadeBuf I__1170 (
            .O(N__6913),
            .I(N__6907));
    CascadeBuf I__1169 (
            .O(N__6910),
            .I(N__6904));
    CascadeMux I__1168 (
            .O(N__6907),
            .I(N__6901));
    CascadeMux I__1167 (
            .O(N__6904),
            .I(N__6898));
    CascadeBuf I__1166 (
            .O(N__6901),
            .I(N__6895));
    CascadeBuf I__1165 (
            .O(N__6898),
            .I(N__6892));
    CascadeMux I__1164 (
            .O(N__6895),
            .I(N__6889));
    CascadeMux I__1163 (
            .O(N__6892),
            .I(N__6886));
    CascadeBuf I__1162 (
            .O(N__6889),
            .I(N__6883));
    CascadeBuf I__1161 (
            .O(N__6886),
            .I(N__6880));
    CascadeMux I__1160 (
            .O(N__6883),
            .I(N__6877));
    CascadeMux I__1159 (
            .O(N__6880),
            .I(N__6874));
    CascadeBuf I__1158 (
            .O(N__6877),
            .I(N__6871));
    CascadeBuf I__1157 (
            .O(N__6874),
            .I(N__6868));
    CascadeMux I__1156 (
            .O(N__6871),
            .I(N__6865));
    CascadeMux I__1155 (
            .O(N__6868),
            .I(N__6862));
    CascadeBuf I__1154 (
            .O(N__6865),
            .I(N__6859));
    CascadeBuf I__1153 (
            .O(N__6862),
            .I(N__6856));
    CascadeMux I__1152 (
            .O(N__6859),
            .I(N__6853));
    CascadeMux I__1151 (
            .O(N__6856),
            .I(N__6850));
    CascadeBuf I__1150 (
            .O(N__6853),
            .I(N__6847));
    InMux I__1149 (
            .O(N__6850),
            .I(N__6844));
    CascadeMux I__1148 (
            .O(N__6847),
            .I(N__6841));
    LocalMux I__1147 (
            .O(N__6844),
            .I(N__6838));
    CascadeBuf I__1146 (
            .O(N__6841),
            .I(N__6835));
    Span4Mux_h I__1145 (
            .O(N__6838),
            .I(N__6832));
    CascadeMux I__1144 (
            .O(N__6835),
            .I(N__6829));
    Span4Mux_h I__1143 (
            .O(N__6832),
            .I(N__6826));
    InMux I__1142 (
            .O(N__6829),
            .I(N__6823));
    Span4Mux_h I__1141 (
            .O(N__6826),
            .I(N__6820));
    LocalMux I__1140 (
            .O(N__6823),
            .I(N__6817));
    Span4Mux_h I__1139 (
            .O(N__6820),
            .I(N__6812));
    Span4Mux_h I__1138 (
            .O(N__6817),
            .I(N__6812));
    Odrv4 I__1137 (
            .O(N__6812),
            .I(waddr_c_9));
    CascadeMux I__1136 (
            .O(N__6809),
            .I(N__6806));
    CascadeBuf I__1135 (
            .O(N__6806),
            .I(N__6803));
    CascadeMux I__1134 (
            .O(N__6803),
            .I(N__6800));
    CascadeBuf I__1133 (
            .O(N__6800),
            .I(N__6796));
    CascadeMux I__1132 (
            .O(N__6799),
            .I(N__6793));
    CascadeMux I__1131 (
            .O(N__6796),
            .I(N__6790));
    CascadeBuf I__1130 (
            .O(N__6793),
            .I(N__6787));
    CascadeBuf I__1129 (
            .O(N__6790),
            .I(N__6784));
    CascadeMux I__1128 (
            .O(N__6787),
            .I(N__6781));
    CascadeMux I__1127 (
            .O(N__6784),
            .I(N__6778));
    CascadeBuf I__1126 (
            .O(N__6781),
            .I(N__6775));
    CascadeBuf I__1125 (
            .O(N__6778),
            .I(N__6772));
    CascadeMux I__1124 (
            .O(N__6775),
            .I(N__6769));
    CascadeMux I__1123 (
            .O(N__6772),
            .I(N__6766));
    CascadeBuf I__1122 (
            .O(N__6769),
            .I(N__6763));
    CascadeBuf I__1121 (
            .O(N__6766),
            .I(N__6760));
    CascadeMux I__1120 (
            .O(N__6763),
            .I(N__6757));
    CascadeMux I__1119 (
            .O(N__6760),
            .I(N__6754));
    CascadeBuf I__1118 (
            .O(N__6757),
            .I(N__6751));
    CascadeBuf I__1117 (
            .O(N__6754),
            .I(N__6748));
    CascadeMux I__1116 (
            .O(N__6751),
            .I(N__6745));
    CascadeMux I__1115 (
            .O(N__6748),
            .I(N__6742));
    CascadeBuf I__1114 (
            .O(N__6745),
            .I(N__6739));
    CascadeBuf I__1113 (
            .O(N__6742),
            .I(N__6736));
    CascadeMux I__1112 (
            .O(N__6739),
            .I(N__6733));
    CascadeMux I__1111 (
            .O(N__6736),
            .I(N__6730));
    CascadeBuf I__1110 (
            .O(N__6733),
            .I(N__6727));
    CascadeBuf I__1109 (
            .O(N__6730),
            .I(N__6724));
    CascadeMux I__1108 (
            .O(N__6727),
            .I(N__6721));
    CascadeMux I__1107 (
            .O(N__6724),
            .I(N__6718));
    CascadeBuf I__1106 (
            .O(N__6721),
            .I(N__6715));
    CascadeBuf I__1105 (
            .O(N__6718),
            .I(N__6712));
    CascadeMux I__1104 (
            .O(N__6715),
            .I(N__6709));
    CascadeMux I__1103 (
            .O(N__6712),
            .I(N__6706));
    CascadeBuf I__1102 (
            .O(N__6709),
            .I(N__6703));
    CascadeBuf I__1101 (
            .O(N__6706),
            .I(N__6700));
    CascadeMux I__1100 (
            .O(N__6703),
            .I(N__6697));
    CascadeMux I__1099 (
            .O(N__6700),
            .I(N__6694));
    CascadeBuf I__1098 (
            .O(N__6697),
            .I(N__6691));
    CascadeBuf I__1097 (
            .O(N__6694),
            .I(N__6688));
    CascadeMux I__1096 (
            .O(N__6691),
            .I(N__6685));
    CascadeMux I__1095 (
            .O(N__6688),
            .I(N__6682));
    CascadeBuf I__1094 (
            .O(N__6685),
            .I(N__6679));
    CascadeBuf I__1093 (
            .O(N__6682),
            .I(N__6676));
    CascadeMux I__1092 (
            .O(N__6679),
            .I(N__6673));
    CascadeMux I__1091 (
            .O(N__6676),
            .I(N__6670));
    CascadeBuf I__1090 (
            .O(N__6673),
            .I(N__6667));
    CascadeBuf I__1089 (
            .O(N__6670),
            .I(N__6664));
    CascadeMux I__1088 (
            .O(N__6667),
            .I(N__6661));
    CascadeMux I__1087 (
            .O(N__6664),
            .I(N__6658));
    CascadeBuf I__1086 (
            .O(N__6661),
            .I(N__6655));
    CascadeBuf I__1085 (
            .O(N__6658),
            .I(N__6652));
    CascadeMux I__1084 (
            .O(N__6655),
            .I(N__6649));
    CascadeMux I__1083 (
            .O(N__6652),
            .I(N__6646));
    CascadeBuf I__1082 (
            .O(N__6649),
            .I(N__6643));
    CascadeBuf I__1081 (
            .O(N__6646),
            .I(N__6640));
    CascadeMux I__1080 (
            .O(N__6643),
            .I(N__6637));
    CascadeMux I__1079 (
            .O(N__6640),
            .I(N__6634));
    CascadeBuf I__1078 (
            .O(N__6637),
            .I(N__6631));
    InMux I__1077 (
            .O(N__6634),
            .I(N__6628));
    CascadeMux I__1076 (
            .O(N__6631),
            .I(N__6625));
    LocalMux I__1075 (
            .O(N__6628),
            .I(N__6622));
    CascadeBuf I__1074 (
            .O(N__6625),
            .I(N__6619));
    Span4Mux_s2_v I__1073 (
            .O(N__6622),
            .I(N__6616));
    CascadeMux I__1072 (
            .O(N__6619),
            .I(N__6613));
    Span4Mux_h I__1071 (
            .O(N__6616),
            .I(N__6610));
    InMux I__1070 (
            .O(N__6613),
            .I(N__6607));
    Sp12to4 I__1069 (
            .O(N__6610),
            .I(N__6604));
    LocalMux I__1068 (
            .O(N__6607),
            .I(N__6601));
    Span12Mux_h I__1067 (
            .O(N__6604),
            .I(N__6596));
    Span12Mux_s2_v I__1066 (
            .O(N__6601),
            .I(N__6596));
    Odrv12 I__1065 (
            .O(N__6596),
            .I(raddr_c_9));
    CascadeMux I__1064 (
            .O(N__6593),
            .I(N__6590));
    CascadeBuf I__1063 (
            .O(N__6590),
            .I(N__6587));
    CascadeMux I__1062 (
            .O(N__6587),
            .I(N__6584));
    CascadeBuf I__1061 (
            .O(N__6584),
            .I(N__6580));
    CascadeMux I__1060 (
            .O(N__6583),
            .I(N__6577));
    CascadeMux I__1059 (
            .O(N__6580),
            .I(N__6574));
    CascadeBuf I__1058 (
            .O(N__6577),
            .I(N__6571));
    CascadeBuf I__1057 (
            .O(N__6574),
            .I(N__6568));
    CascadeMux I__1056 (
            .O(N__6571),
            .I(N__6565));
    CascadeMux I__1055 (
            .O(N__6568),
            .I(N__6562));
    CascadeBuf I__1054 (
            .O(N__6565),
            .I(N__6559));
    CascadeBuf I__1053 (
            .O(N__6562),
            .I(N__6556));
    CascadeMux I__1052 (
            .O(N__6559),
            .I(N__6553));
    CascadeMux I__1051 (
            .O(N__6556),
            .I(N__6550));
    CascadeBuf I__1050 (
            .O(N__6553),
            .I(N__6547));
    CascadeBuf I__1049 (
            .O(N__6550),
            .I(N__6544));
    CascadeMux I__1048 (
            .O(N__6547),
            .I(N__6541));
    CascadeMux I__1047 (
            .O(N__6544),
            .I(N__6538));
    CascadeBuf I__1046 (
            .O(N__6541),
            .I(N__6535));
    CascadeBuf I__1045 (
            .O(N__6538),
            .I(N__6532));
    CascadeMux I__1044 (
            .O(N__6535),
            .I(N__6529));
    CascadeMux I__1043 (
            .O(N__6532),
            .I(N__6526));
    CascadeBuf I__1042 (
            .O(N__6529),
            .I(N__6523));
    CascadeBuf I__1041 (
            .O(N__6526),
            .I(N__6520));
    CascadeMux I__1040 (
            .O(N__6523),
            .I(N__6517));
    CascadeMux I__1039 (
            .O(N__6520),
            .I(N__6514));
    CascadeBuf I__1038 (
            .O(N__6517),
            .I(N__6511));
    CascadeBuf I__1037 (
            .O(N__6514),
            .I(N__6508));
    CascadeMux I__1036 (
            .O(N__6511),
            .I(N__6505));
    CascadeMux I__1035 (
            .O(N__6508),
            .I(N__6502));
    CascadeBuf I__1034 (
            .O(N__6505),
            .I(N__6499));
    CascadeBuf I__1033 (
            .O(N__6502),
            .I(N__6496));
    CascadeMux I__1032 (
            .O(N__6499),
            .I(N__6493));
    CascadeMux I__1031 (
            .O(N__6496),
            .I(N__6490));
    CascadeBuf I__1030 (
            .O(N__6493),
            .I(N__6487));
    CascadeBuf I__1029 (
            .O(N__6490),
            .I(N__6484));
    CascadeMux I__1028 (
            .O(N__6487),
            .I(N__6481));
    CascadeMux I__1027 (
            .O(N__6484),
            .I(N__6478));
    CascadeBuf I__1026 (
            .O(N__6481),
            .I(N__6475));
    CascadeBuf I__1025 (
            .O(N__6478),
            .I(N__6472));
    CascadeMux I__1024 (
            .O(N__6475),
            .I(N__6469));
    CascadeMux I__1023 (
            .O(N__6472),
            .I(N__6466));
    CascadeBuf I__1022 (
            .O(N__6469),
            .I(N__6463));
    CascadeBuf I__1021 (
            .O(N__6466),
            .I(N__6460));
    CascadeMux I__1020 (
            .O(N__6463),
            .I(N__6457));
    CascadeMux I__1019 (
            .O(N__6460),
            .I(N__6454));
    CascadeBuf I__1018 (
            .O(N__6457),
            .I(N__6451));
    CascadeBuf I__1017 (
            .O(N__6454),
            .I(N__6448));
    CascadeMux I__1016 (
            .O(N__6451),
            .I(N__6445));
    CascadeMux I__1015 (
            .O(N__6448),
            .I(N__6442));
    CascadeBuf I__1014 (
            .O(N__6445),
            .I(N__6439));
    CascadeBuf I__1013 (
            .O(N__6442),
            .I(N__6436));
    CascadeMux I__1012 (
            .O(N__6439),
            .I(N__6433));
    CascadeMux I__1011 (
            .O(N__6436),
            .I(N__6430));
    CascadeBuf I__1010 (
            .O(N__6433),
            .I(N__6427));
    CascadeBuf I__1009 (
            .O(N__6430),
            .I(N__6424));
    CascadeMux I__1008 (
            .O(N__6427),
            .I(N__6421));
    CascadeMux I__1007 (
            .O(N__6424),
            .I(N__6418));
    CascadeBuf I__1006 (
            .O(N__6421),
            .I(N__6415));
    InMux I__1005 (
            .O(N__6418),
            .I(N__6412));
    CascadeMux I__1004 (
            .O(N__6415),
            .I(N__6409));
    LocalMux I__1003 (
            .O(N__6412),
            .I(N__6406));
    CascadeBuf I__1002 (
            .O(N__6409),
            .I(N__6403));
    Span4Mux_h I__1001 (
            .O(N__6406),
            .I(N__6400));
    CascadeMux I__1000 (
            .O(N__6403),
            .I(N__6397));
    Span4Mux_h I__999 (
            .O(N__6400),
            .I(N__6394));
    InMux I__998 (
            .O(N__6397),
            .I(N__6391));
    Span4Mux_h I__997 (
            .O(N__6394),
            .I(N__6388));
    LocalMux I__996 (
            .O(N__6391),
            .I(N__6385));
    Span4Mux_h I__995 (
            .O(N__6388),
            .I(N__6380));
    Span4Mux_h I__994 (
            .O(N__6385),
            .I(N__6380));
    Odrv4 I__993 (
            .O(N__6380),
            .I(waddr_c_7));
    CascadeMux I__992 (
            .O(N__6377),
            .I(N__6374));
    CascadeBuf I__991 (
            .O(N__6374),
            .I(N__6371));
    CascadeMux I__990 (
            .O(N__6371),
            .I(N__6368));
    CascadeBuf I__989 (
            .O(N__6368),
            .I(N__6364));
    CascadeMux I__988 (
            .O(N__6367),
            .I(N__6361));
    CascadeMux I__987 (
            .O(N__6364),
            .I(N__6358));
    CascadeBuf I__986 (
            .O(N__6361),
            .I(N__6355));
    CascadeBuf I__985 (
            .O(N__6358),
            .I(N__6352));
    CascadeMux I__984 (
            .O(N__6355),
            .I(N__6349));
    CascadeMux I__983 (
            .O(N__6352),
            .I(N__6346));
    CascadeBuf I__982 (
            .O(N__6349),
            .I(N__6343));
    CascadeBuf I__981 (
            .O(N__6346),
            .I(N__6340));
    CascadeMux I__980 (
            .O(N__6343),
            .I(N__6337));
    CascadeMux I__979 (
            .O(N__6340),
            .I(N__6334));
    CascadeBuf I__978 (
            .O(N__6337),
            .I(N__6331));
    CascadeBuf I__977 (
            .O(N__6334),
            .I(N__6328));
    CascadeMux I__976 (
            .O(N__6331),
            .I(N__6325));
    CascadeMux I__975 (
            .O(N__6328),
            .I(N__6322));
    CascadeBuf I__974 (
            .O(N__6325),
            .I(N__6319));
    CascadeBuf I__973 (
            .O(N__6322),
            .I(N__6316));
    CascadeMux I__972 (
            .O(N__6319),
            .I(N__6313));
    CascadeMux I__971 (
            .O(N__6316),
            .I(N__6310));
    CascadeBuf I__970 (
            .O(N__6313),
            .I(N__6307));
    CascadeBuf I__969 (
            .O(N__6310),
            .I(N__6304));
    CascadeMux I__968 (
            .O(N__6307),
            .I(N__6301));
    CascadeMux I__967 (
            .O(N__6304),
            .I(N__6298));
    CascadeBuf I__966 (
            .O(N__6301),
            .I(N__6295));
    CascadeBuf I__965 (
            .O(N__6298),
            .I(N__6292));
    CascadeMux I__964 (
            .O(N__6295),
            .I(N__6289));
    CascadeMux I__963 (
            .O(N__6292),
            .I(N__6286));
    CascadeBuf I__962 (
            .O(N__6289),
            .I(N__6283));
    CascadeBuf I__961 (
            .O(N__6286),
            .I(N__6280));
    CascadeMux I__960 (
            .O(N__6283),
            .I(N__6277));
    CascadeMux I__959 (
            .O(N__6280),
            .I(N__6274));
    CascadeBuf I__958 (
            .O(N__6277),
            .I(N__6271));
    CascadeBuf I__957 (
            .O(N__6274),
            .I(N__6268));
    CascadeMux I__956 (
            .O(N__6271),
            .I(N__6265));
    CascadeMux I__955 (
            .O(N__6268),
            .I(N__6262));
    CascadeBuf I__954 (
            .O(N__6265),
            .I(N__6259));
    CascadeBuf I__953 (
            .O(N__6262),
            .I(N__6256));
    CascadeMux I__952 (
            .O(N__6259),
            .I(N__6253));
    CascadeMux I__951 (
            .O(N__6256),
            .I(N__6250));
    CascadeBuf I__950 (
            .O(N__6253),
            .I(N__6247));
    CascadeBuf I__949 (
            .O(N__6250),
            .I(N__6244));
    CascadeMux I__948 (
            .O(N__6247),
            .I(N__6241));
    CascadeMux I__947 (
            .O(N__6244),
            .I(N__6238));
    CascadeBuf I__946 (
            .O(N__6241),
            .I(N__6235));
    CascadeBuf I__945 (
            .O(N__6238),
            .I(N__6232));
    CascadeMux I__944 (
            .O(N__6235),
            .I(N__6229));
    CascadeMux I__943 (
            .O(N__6232),
            .I(N__6226));
    CascadeBuf I__942 (
            .O(N__6229),
            .I(N__6223));
    CascadeBuf I__941 (
            .O(N__6226),
            .I(N__6220));
    CascadeMux I__940 (
            .O(N__6223),
            .I(N__6217));
    CascadeMux I__939 (
            .O(N__6220),
            .I(N__6214));
    CascadeBuf I__938 (
            .O(N__6217),
            .I(N__6211));
    CascadeBuf I__937 (
            .O(N__6214),
            .I(N__6208));
    CascadeMux I__936 (
            .O(N__6211),
            .I(N__6205));
    CascadeMux I__935 (
            .O(N__6208),
            .I(N__6202));
    CascadeBuf I__934 (
            .O(N__6205),
            .I(N__6199));
    InMux I__933 (
            .O(N__6202),
            .I(N__6196));
    CascadeMux I__932 (
            .O(N__6199),
            .I(N__6193));
    LocalMux I__931 (
            .O(N__6196),
            .I(N__6190));
    CascadeBuf I__930 (
            .O(N__6193),
            .I(N__6187));
    Span4Mux_v I__929 (
            .O(N__6190),
            .I(N__6184));
    CascadeMux I__928 (
            .O(N__6187),
            .I(N__6181));
    Sp12to4 I__927 (
            .O(N__6184),
            .I(N__6178));
    InMux I__926 (
            .O(N__6181),
            .I(N__6175));
    Span12Mux_h I__925 (
            .O(N__6178),
            .I(N__6172));
    LocalMux I__924 (
            .O(N__6175),
            .I(N__6169));
    Span12Mux_v I__923 (
            .O(N__6172),
            .I(N__6166));
    Span12Mux_v I__922 (
            .O(N__6169),
            .I(N__6163));
    Odrv12 I__921 (
            .O(N__6166),
            .I(raddr_c_0));
    Odrv12 I__920 (
            .O(N__6163),
            .I(raddr_c_0));
    CascadeMux I__919 (
            .O(N__6158),
            .I(N__6155));
    CascadeBuf I__918 (
            .O(N__6155),
            .I(N__6152));
    CascadeMux I__917 (
            .O(N__6152),
            .I(N__6149));
    CascadeBuf I__916 (
            .O(N__6149),
            .I(N__6146));
    CascadeMux I__915 (
            .O(N__6146),
            .I(N__6142));
    CascadeMux I__914 (
            .O(N__6145),
            .I(N__6139));
    CascadeBuf I__913 (
            .O(N__6142),
            .I(N__6136));
    CascadeBuf I__912 (
            .O(N__6139),
            .I(N__6133));
    CascadeMux I__911 (
            .O(N__6136),
            .I(N__6130));
    CascadeMux I__910 (
            .O(N__6133),
            .I(N__6127));
    CascadeBuf I__909 (
            .O(N__6130),
            .I(N__6124));
    CascadeBuf I__908 (
            .O(N__6127),
            .I(N__6121));
    CascadeMux I__907 (
            .O(N__6124),
            .I(N__6118));
    CascadeMux I__906 (
            .O(N__6121),
            .I(N__6115));
    CascadeBuf I__905 (
            .O(N__6118),
            .I(N__6112));
    CascadeBuf I__904 (
            .O(N__6115),
            .I(N__6109));
    CascadeMux I__903 (
            .O(N__6112),
            .I(N__6106));
    CascadeMux I__902 (
            .O(N__6109),
            .I(N__6103));
    CascadeBuf I__901 (
            .O(N__6106),
            .I(N__6100));
    CascadeBuf I__900 (
            .O(N__6103),
            .I(N__6097));
    CascadeMux I__899 (
            .O(N__6100),
            .I(N__6094));
    CascadeMux I__898 (
            .O(N__6097),
            .I(N__6091));
    CascadeBuf I__897 (
            .O(N__6094),
            .I(N__6088));
    CascadeBuf I__896 (
            .O(N__6091),
            .I(N__6085));
    CascadeMux I__895 (
            .O(N__6088),
            .I(N__6082));
    CascadeMux I__894 (
            .O(N__6085),
            .I(N__6079));
    CascadeBuf I__893 (
            .O(N__6082),
            .I(N__6076));
    CascadeBuf I__892 (
            .O(N__6079),
            .I(N__6073));
    CascadeMux I__891 (
            .O(N__6076),
            .I(N__6070));
    CascadeMux I__890 (
            .O(N__6073),
            .I(N__6067));
    CascadeBuf I__889 (
            .O(N__6070),
            .I(N__6064));
    CascadeBuf I__888 (
            .O(N__6067),
            .I(N__6061));
    CascadeMux I__887 (
            .O(N__6064),
            .I(N__6058));
    CascadeMux I__886 (
            .O(N__6061),
            .I(N__6055));
    CascadeBuf I__885 (
            .O(N__6058),
            .I(N__6052));
    CascadeBuf I__884 (
            .O(N__6055),
            .I(N__6049));
    CascadeMux I__883 (
            .O(N__6052),
            .I(N__6046));
    CascadeMux I__882 (
            .O(N__6049),
            .I(N__6043));
    CascadeBuf I__881 (
            .O(N__6046),
            .I(N__6040));
    CascadeBuf I__880 (
            .O(N__6043),
            .I(N__6037));
    CascadeMux I__879 (
            .O(N__6040),
            .I(N__6034));
    CascadeMux I__878 (
            .O(N__6037),
            .I(N__6031));
    CascadeBuf I__877 (
            .O(N__6034),
            .I(N__6028));
    CascadeBuf I__876 (
            .O(N__6031),
            .I(N__6025));
    CascadeMux I__875 (
            .O(N__6028),
            .I(N__6022));
    CascadeMux I__874 (
            .O(N__6025),
            .I(N__6019));
    CascadeBuf I__873 (
            .O(N__6022),
            .I(N__6016));
    CascadeBuf I__872 (
            .O(N__6019),
            .I(N__6013));
    CascadeMux I__871 (
            .O(N__6016),
            .I(N__6010));
    CascadeMux I__870 (
            .O(N__6013),
            .I(N__6007));
    CascadeBuf I__869 (
            .O(N__6010),
            .I(N__6004));
    CascadeBuf I__868 (
            .O(N__6007),
            .I(N__6001));
    CascadeMux I__867 (
            .O(N__6004),
            .I(N__5998));
    CascadeMux I__866 (
            .O(N__6001),
            .I(N__5995));
    CascadeBuf I__865 (
            .O(N__5998),
            .I(N__5992));
    CascadeBuf I__864 (
            .O(N__5995),
            .I(N__5989));
    CascadeMux I__863 (
            .O(N__5992),
            .I(N__5986));
    CascadeMux I__862 (
            .O(N__5989),
            .I(N__5983));
    InMux I__861 (
            .O(N__5986),
            .I(N__5980));
    CascadeBuf I__860 (
            .O(N__5983),
            .I(N__5977));
    LocalMux I__859 (
            .O(N__5980),
            .I(N__5974));
    CascadeMux I__858 (
            .O(N__5977),
            .I(N__5971));
    Span4Mux_h I__857 (
            .O(N__5974),
            .I(N__5968));
    CascadeBuf I__856 (
            .O(N__5971),
            .I(N__5965));
    Span4Mux_h I__855 (
            .O(N__5968),
            .I(N__5962));
    CascadeMux I__854 (
            .O(N__5965),
            .I(N__5959));
    Span4Mux_h I__853 (
            .O(N__5962),
            .I(N__5956));
    InMux I__852 (
            .O(N__5959),
            .I(N__5953));
    Span4Mux_h I__851 (
            .O(N__5956),
            .I(N__5948));
    LocalMux I__850 (
            .O(N__5953),
            .I(N__5948));
    Span4Mux_h I__849 (
            .O(N__5948),
            .I(N__5945));
    Span4Mux_h I__848 (
            .O(N__5945),
            .I(N__5942));
    Odrv4 I__847 (
            .O(N__5942),
            .I(waddr_c_10));
    CascadeMux I__846 (
            .O(N__5939),
            .I(N__5936));
    CascadeBuf I__845 (
            .O(N__5936),
            .I(N__5933));
    CascadeMux I__844 (
            .O(N__5933),
            .I(N__5930));
    CascadeBuf I__843 (
            .O(N__5930),
            .I(N__5926));
    CascadeMux I__842 (
            .O(N__5929),
            .I(N__5923));
    CascadeMux I__841 (
            .O(N__5926),
            .I(N__5920));
    CascadeBuf I__840 (
            .O(N__5923),
            .I(N__5917));
    CascadeBuf I__839 (
            .O(N__5920),
            .I(N__5914));
    CascadeMux I__838 (
            .O(N__5917),
            .I(N__5911));
    CascadeMux I__837 (
            .O(N__5914),
            .I(N__5908));
    CascadeBuf I__836 (
            .O(N__5911),
            .I(N__5905));
    CascadeBuf I__835 (
            .O(N__5908),
            .I(N__5902));
    CascadeMux I__834 (
            .O(N__5905),
            .I(N__5899));
    CascadeMux I__833 (
            .O(N__5902),
            .I(N__5896));
    CascadeBuf I__832 (
            .O(N__5899),
            .I(N__5893));
    CascadeBuf I__831 (
            .O(N__5896),
            .I(N__5890));
    CascadeMux I__830 (
            .O(N__5893),
            .I(N__5887));
    CascadeMux I__829 (
            .O(N__5890),
            .I(N__5884));
    CascadeBuf I__828 (
            .O(N__5887),
            .I(N__5881));
    CascadeBuf I__827 (
            .O(N__5884),
            .I(N__5878));
    CascadeMux I__826 (
            .O(N__5881),
            .I(N__5875));
    CascadeMux I__825 (
            .O(N__5878),
            .I(N__5872));
    CascadeBuf I__824 (
            .O(N__5875),
            .I(N__5869));
    CascadeBuf I__823 (
            .O(N__5872),
            .I(N__5866));
    CascadeMux I__822 (
            .O(N__5869),
            .I(N__5863));
    CascadeMux I__821 (
            .O(N__5866),
            .I(N__5860));
    CascadeBuf I__820 (
            .O(N__5863),
            .I(N__5857));
    CascadeBuf I__819 (
            .O(N__5860),
            .I(N__5854));
    CascadeMux I__818 (
            .O(N__5857),
            .I(N__5851));
    CascadeMux I__817 (
            .O(N__5854),
            .I(N__5848));
    CascadeBuf I__816 (
            .O(N__5851),
            .I(N__5845));
    CascadeBuf I__815 (
            .O(N__5848),
            .I(N__5842));
    CascadeMux I__814 (
            .O(N__5845),
            .I(N__5839));
    CascadeMux I__813 (
            .O(N__5842),
            .I(N__5836));
    CascadeBuf I__812 (
            .O(N__5839),
            .I(N__5833));
    CascadeBuf I__811 (
            .O(N__5836),
            .I(N__5830));
    CascadeMux I__810 (
            .O(N__5833),
            .I(N__5827));
    CascadeMux I__809 (
            .O(N__5830),
            .I(N__5824));
    CascadeBuf I__808 (
            .O(N__5827),
            .I(N__5821));
    CascadeBuf I__807 (
            .O(N__5824),
            .I(N__5818));
    CascadeMux I__806 (
            .O(N__5821),
            .I(N__5815));
    CascadeMux I__805 (
            .O(N__5818),
            .I(N__5812));
    CascadeBuf I__804 (
            .O(N__5815),
            .I(N__5809));
    CascadeBuf I__803 (
            .O(N__5812),
            .I(N__5806));
    CascadeMux I__802 (
            .O(N__5809),
            .I(N__5803));
    CascadeMux I__801 (
            .O(N__5806),
            .I(N__5800));
    CascadeBuf I__800 (
            .O(N__5803),
            .I(N__5797));
    CascadeBuf I__799 (
            .O(N__5800),
            .I(N__5794));
    CascadeMux I__798 (
            .O(N__5797),
            .I(N__5791));
    CascadeMux I__797 (
            .O(N__5794),
            .I(N__5788));
    CascadeBuf I__796 (
            .O(N__5791),
            .I(N__5785));
    CascadeBuf I__795 (
            .O(N__5788),
            .I(N__5782));
    CascadeMux I__794 (
            .O(N__5785),
            .I(N__5779));
    CascadeMux I__793 (
            .O(N__5782),
            .I(N__5776));
    CascadeBuf I__792 (
            .O(N__5779),
            .I(N__5773));
    CascadeBuf I__791 (
            .O(N__5776),
            .I(N__5770));
    CascadeMux I__790 (
            .O(N__5773),
            .I(N__5767));
    CascadeMux I__789 (
            .O(N__5770),
            .I(N__5764));
    CascadeBuf I__788 (
            .O(N__5767),
            .I(N__5761));
    InMux I__787 (
            .O(N__5764),
            .I(N__5758));
    CascadeMux I__786 (
            .O(N__5761),
            .I(N__5755));
    LocalMux I__785 (
            .O(N__5758),
            .I(N__5752));
    CascadeBuf I__784 (
            .O(N__5755),
            .I(N__5749));
    Span4Mux_h I__783 (
            .O(N__5752),
            .I(N__5746));
    CascadeMux I__782 (
            .O(N__5749),
            .I(N__5743));
    Span4Mux_h I__781 (
            .O(N__5746),
            .I(N__5740));
    InMux I__780 (
            .O(N__5743),
            .I(N__5737));
    Span4Mux_h I__779 (
            .O(N__5740),
            .I(N__5734));
    LocalMux I__778 (
            .O(N__5737),
            .I(N__5731));
    Span4Mux_h I__777 (
            .O(N__5734),
            .I(N__5726));
    Span4Mux_h I__776 (
            .O(N__5731),
            .I(N__5726));
    Odrv4 I__775 (
            .O(N__5726),
            .I(waddr_c_8));
    CascadeMux I__774 (
            .O(N__5723),
            .I(N__5720));
    CascadeBuf I__773 (
            .O(N__5720),
            .I(N__5716));
    CascadeMux I__772 (
            .O(N__5719),
            .I(N__5713));
    CascadeMux I__771 (
            .O(N__5716),
            .I(N__5710));
    CascadeBuf I__770 (
            .O(N__5713),
            .I(N__5707));
    CascadeBuf I__769 (
            .O(N__5710),
            .I(N__5704));
    CascadeMux I__768 (
            .O(N__5707),
            .I(N__5701));
    CascadeMux I__767 (
            .O(N__5704),
            .I(N__5698));
    CascadeBuf I__766 (
            .O(N__5701),
            .I(N__5695));
    CascadeBuf I__765 (
            .O(N__5698),
            .I(N__5692));
    CascadeMux I__764 (
            .O(N__5695),
            .I(N__5689));
    CascadeMux I__763 (
            .O(N__5692),
            .I(N__5686));
    CascadeBuf I__762 (
            .O(N__5689),
            .I(N__5683));
    CascadeBuf I__761 (
            .O(N__5686),
            .I(N__5680));
    CascadeMux I__760 (
            .O(N__5683),
            .I(N__5677));
    CascadeMux I__759 (
            .O(N__5680),
            .I(N__5674));
    CascadeBuf I__758 (
            .O(N__5677),
            .I(N__5671));
    CascadeBuf I__757 (
            .O(N__5674),
            .I(N__5668));
    CascadeMux I__756 (
            .O(N__5671),
            .I(N__5665));
    CascadeMux I__755 (
            .O(N__5668),
            .I(N__5662));
    CascadeBuf I__754 (
            .O(N__5665),
            .I(N__5659));
    CascadeBuf I__753 (
            .O(N__5662),
            .I(N__5656));
    CascadeMux I__752 (
            .O(N__5659),
            .I(N__5653));
    CascadeMux I__751 (
            .O(N__5656),
            .I(N__5650));
    CascadeBuf I__750 (
            .O(N__5653),
            .I(N__5647));
    CascadeBuf I__749 (
            .O(N__5650),
            .I(N__5644));
    CascadeMux I__748 (
            .O(N__5647),
            .I(N__5641));
    CascadeMux I__747 (
            .O(N__5644),
            .I(N__5638));
    CascadeBuf I__746 (
            .O(N__5641),
            .I(N__5635));
    CascadeBuf I__745 (
            .O(N__5638),
            .I(N__5632));
    CascadeMux I__744 (
            .O(N__5635),
            .I(N__5629));
    CascadeMux I__743 (
            .O(N__5632),
            .I(N__5626));
    CascadeBuf I__742 (
            .O(N__5629),
            .I(N__5623));
    CascadeBuf I__741 (
            .O(N__5626),
            .I(N__5620));
    CascadeMux I__740 (
            .O(N__5623),
            .I(N__5617));
    CascadeMux I__739 (
            .O(N__5620),
            .I(N__5614));
    CascadeBuf I__738 (
            .O(N__5617),
            .I(N__5611));
    CascadeBuf I__737 (
            .O(N__5614),
            .I(N__5608));
    CascadeMux I__736 (
            .O(N__5611),
            .I(N__5605));
    CascadeMux I__735 (
            .O(N__5608),
            .I(N__5602));
    CascadeBuf I__734 (
            .O(N__5605),
            .I(N__5599));
    CascadeBuf I__733 (
            .O(N__5602),
            .I(N__5596));
    CascadeMux I__732 (
            .O(N__5599),
            .I(N__5593));
    CascadeMux I__731 (
            .O(N__5596),
            .I(N__5590));
    CascadeBuf I__730 (
            .O(N__5593),
            .I(N__5587));
    CascadeBuf I__729 (
            .O(N__5590),
            .I(N__5584));
    CascadeMux I__728 (
            .O(N__5587),
            .I(N__5581));
    CascadeMux I__727 (
            .O(N__5584),
            .I(N__5578));
    CascadeBuf I__726 (
            .O(N__5581),
            .I(N__5575));
    CascadeBuf I__725 (
            .O(N__5578),
            .I(N__5572));
    CascadeMux I__724 (
            .O(N__5575),
            .I(N__5569));
    CascadeMux I__723 (
            .O(N__5572),
            .I(N__5566));
    CascadeBuf I__722 (
            .O(N__5569),
            .I(N__5563));
    CascadeBuf I__721 (
            .O(N__5566),
            .I(N__5560));
    CascadeMux I__720 (
            .O(N__5563),
            .I(N__5557));
    CascadeMux I__719 (
            .O(N__5560),
            .I(N__5554));
    CascadeBuf I__718 (
            .O(N__5557),
            .I(N__5551));
    CascadeBuf I__717 (
            .O(N__5554),
            .I(N__5548));
    CascadeMux I__716 (
            .O(N__5551),
            .I(N__5545));
    CascadeMux I__715 (
            .O(N__5548),
            .I(N__5542));
    CascadeBuf I__714 (
            .O(N__5545),
            .I(N__5539));
    InMux I__713 (
            .O(N__5542),
            .I(N__5536));
    CascadeMux I__712 (
            .O(N__5539),
            .I(N__5533));
    LocalMux I__711 (
            .O(N__5536),
            .I(N__5530));
    InMux I__710 (
            .O(N__5533),
            .I(N__5527));
    Span4Mux_v I__709 (
            .O(N__5530),
            .I(N__5524));
    LocalMux I__708 (
            .O(N__5527),
            .I(N__5521));
    Span4Mux_h I__707 (
            .O(N__5524),
            .I(N__5518));
    Span4Mux_v I__706 (
            .O(N__5521),
            .I(N__5515));
    Sp12to4 I__705 (
            .O(N__5518),
            .I(N__5512));
    Span4Mux_v I__704 (
            .O(N__5515),
            .I(N__5509));
    Span12Mux_v I__703 (
            .O(N__5512),
            .I(N__5506));
    Span4Mux_v I__702 (
            .O(N__5509),
            .I(N__5503));
    Span12Mux_h I__701 (
            .O(N__5506),
            .I(N__5498));
    Sp12to4 I__700 (
            .O(N__5503),
            .I(N__5498));
    Odrv12 I__699 (
            .O(N__5498),
            .I(raddr_c_1));
    CascadeMux I__698 (
            .O(N__5495),
            .I(N__5492));
    CascadeBuf I__697 (
            .O(N__5492),
            .I(N__5488));
    CascadeMux I__696 (
            .O(N__5491),
            .I(N__5485));
    CascadeMux I__695 (
            .O(N__5488),
            .I(N__5482));
    CascadeBuf I__694 (
            .O(N__5485),
            .I(N__5479));
    CascadeBuf I__693 (
            .O(N__5482),
            .I(N__5476));
    CascadeMux I__692 (
            .O(N__5479),
            .I(N__5473));
    CascadeMux I__691 (
            .O(N__5476),
            .I(N__5470));
    CascadeBuf I__690 (
            .O(N__5473),
            .I(N__5467));
    CascadeBuf I__689 (
            .O(N__5470),
            .I(N__5464));
    CascadeMux I__688 (
            .O(N__5467),
            .I(N__5461));
    CascadeMux I__687 (
            .O(N__5464),
            .I(N__5458));
    CascadeBuf I__686 (
            .O(N__5461),
            .I(N__5455));
    CascadeBuf I__685 (
            .O(N__5458),
            .I(N__5452));
    CascadeMux I__684 (
            .O(N__5455),
            .I(N__5449));
    CascadeMux I__683 (
            .O(N__5452),
            .I(N__5446));
    CascadeBuf I__682 (
            .O(N__5449),
            .I(N__5443));
    CascadeBuf I__681 (
            .O(N__5446),
            .I(N__5440));
    CascadeMux I__680 (
            .O(N__5443),
            .I(N__5437));
    CascadeMux I__679 (
            .O(N__5440),
            .I(N__5434));
    CascadeBuf I__678 (
            .O(N__5437),
            .I(N__5431));
    CascadeBuf I__677 (
            .O(N__5434),
            .I(N__5428));
    CascadeMux I__676 (
            .O(N__5431),
            .I(N__5425));
    CascadeMux I__675 (
            .O(N__5428),
            .I(N__5422));
    CascadeBuf I__674 (
            .O(N__5425),
            .I(N__5419));
    CascadeBuf I__673 (
            .O(N__5422),
            .I(N__5416));
    CascadeMux I__672 (
            .O(N__5419),
            .I(N__5413));
    CascadeMux I__671 (
            .O(N__5416),
            .I(N__5410));
    CascadeBuf I__670 (
            .O(N__5413),
            .I(N__5407));
    CascadeBuf I__669 (
            .O(N__5410),
            .I(N__5404));
    CascadeMux I__668 (
            .O(N__5407),
            .I(N__5401));
    CascadeMux I__667 (
            .O(N__5404),
            .I(N__5398));
    CascadeBuf I__666 (
            .O(N__5401),
            .I(N__5395));
    CascadeBuf I__665 (
            .O(N__5398),
            .I(N__5392));
    CascadeMux I__664 (
            .O(N__5395),
            .I(N__5389));
    CascadeMux I__663 (
            .O(N__5392),
            .I(N__5386));
    CascadeBuf I__662 (
            .O(N__5389),
            .I(N__5383));
    CascadeBuf I__661 (
            .O(N__5386),
            .I(N__5380));
    CascadeMux I__660 (
            .O(N__5383),
            .I(N__5377));
    CascadeMux I__659 (
            .O(N__5380),
            .I(N__5374));
    CascadeBuf I__658 (
            .O(N__5377),
            .I(N__5371));
    CascadeBuf I__657 (
            .O(N__5374),
            .I(N__5368));
    CascadeMux I__656 (
            .O(N__5371),
            .I(N__5365));
    CascadeMux I__655 (
            .O(N__5368),
            .I(N__5362));
    CascadeBuf I__654 (
            .O(N__5365),
            .I(N__5359));
    CascadeBuf I__653 (
            .O(N__5362),
            .I(N__5356));
    CascadeMux I__652 (
            .O(N__5359),
            .I(N__5353));
    CascadeMux I__651 (
            .O(N__5356),
            .I(N__5350));
    CascadeBuf I__650 (
            .O(N__5353),
            .I(N__5347));
    CascadeBuf I__649 (
            .O(N__5350),
            .I(N__5344));
    CascadeMux I__648 (
            .O(N__5347),
            .I(N__5341));
    CascadeMux I__647 (
            .O(N__5344),
            .I(N__5338));
    CascadeBuf I__646 (
            .O(N__5341),
            .I(N__5335));
    CascadeBuf I__645 (
            .O(N__5338),
            .I(N__5332));
    CascadeMux I__644 (
            .O(N__5335),
            .I(N__5329));
    CascadeMux I__643 (
            .O(N__5332),
            .I(N__5326));
    CascadeBuf I__642 (
            .O(N__5329),
            .I(N__5323));
    CascadeBuf I__641 (
            .O(N__5326),
            .I(N__5320));
    CascadeMux I__640 (
            .O(N__5323),
            .I(N__5317));
    CascadeMux I__639 (
            .O(N__5320),
            .I(N__5314));
    CascadeBuf I__638 (
            .O(N__5317),
            .I(N__5311));
    InMux I__637 (
            .O(N__5314),
            .I(N__5308));
    CascadeMux I__636 (
            .O(N__5311),
            .I(N__5305));
    LocalMux I__635 (
            .O(N__5308),
            .I(N__5302));
    InMux I__634 (
            .O(N__5305),
            .I(N__5299));
    Span4Mux_h I__633 (
            .O(N__5302),
            .I(N__5296));
    LocalMux I__632 (
            .O(N__5299),
            .I(N__5293));
    Sp12to4 I__631 (
            .O(N__5296),
            .I(N__5290));
    Span4Mux_s3_v I__630 (
            .O(N__5293),
            .I(N__5287));
    Span12Mux_s7_v I__629 (
            .O(N__5290),
            .I(N__5284));
    Span4Mux_h I__628 (
            .O(N__5287),
            .I(N__5281));
    Span12Mux_h I__627 (
            .O(N__5284),
            .I(N__5278));
    Span4Mux_v I__626 (
            .O(N__5281),
            .I(N__5275));
    Odrv12 I__625 (
            .O(N__5278),
            .I(raddr_c_6));
    Odrv4 I__624 (
            .O(N__5275),
            .I(raddr_c_6));
    CascadeMux I__623 (
            .O(N__5270),
            .I(N__5267));
    CascadeBuf I__622 (
            .O(N__5267),
            .I(N__5264));
    CascadeMux I__621 (
            .O(N__5264),
            .I(N__5261));
    CascadeBuf I__620 (
            .O(N__5261),
            .I(N__5258));
    CascadeMux I__619 (
            .O(N__5258),
            .I(N__5254));
    CascadeMux I__618 (
            .O(N__5257),
            .I(N__5251));
    CascadeBuf I__617 (
            .O(N__5254),
            .I(N__5248));
    CascadeBuf I__616 (
            .O(N__5251),
            .I(N__5245));
    CascadeMux I__615 (
            .O(N__5248),
            .I(N__5242));
    CascadeMux I__614 (
            .O(N__5245),
            .I(N__5239));
    CascadeBuf I__613 (
            .O(N__5242),
            .I(N__5236));
    CascadeBuf I__612 (
            .O(N__5239),
            .I(N__5233));
    CascadeMux I__611 (
            .O(N__5236),
            .I(N__5230));
    CascadeMux I__610 (
            .O(N__5233),
            .I(N__5227));
    CascadeBuf I__609 (
            .O(N__5230),
            .I(N__5224));
    CascadeBuf I__608 (
            .O(N__5227),
            .I(N__5221));
    CascadeMux I__607 (
            .O(N__5224),
            .I(N__5218));
    CascadeMux I__606 (
            .O(N__5221),
            .I(N__5215));
    CascadeBuf I__605 (
            .O(N__5218),
            .I(N__5212));
    CascadeBuf I__604 (
            .O(N__5215),
            .I(N__5209));
    CascadeMux I__603 (
            .O(N__5212),
            .I(N__5206));
    CascadeMux I__602 (
            .O(N__5209),
            .I(N__5203));
    CascadeBuf I__601 (
            .O(N__5206),
            .I(N__5200));
    CascadeBuf I__600 (
            .O(N__5203),
            .I(N__5197));
    CascadeMux I__599 (
            .O(N__5200),
            .I(N__5194));
    CascadeMux I__598 (
            .O(N__5197),
            .I(N__5191));
    CascadeBuf I__597 (
            .O(N__5194),
            .I(N__5188));
    CascadeBuf I__596 (
            .O(N__5191),
            .I(N__5185));
    CascadeMux I__595 (
            .O(N__5188),
            .I(N__5182));
    CascadeMux I__594 (
            .O(N__5185),
            .I(N__5179));
    CascadeBuf I__593 (
            .O(N__5182),
            .I(N__5176));
    CascadeBuf I__592 (
            .O(N__5179),
            .I(N__5173));
    CascadeMux I__591 (
            .O(N__5176),
            .I(N__5170));
    CascadeMux I__590 (
            .O(N__5173),
            .I(N__5167));
    CascadeBuf I__589 (
            .O(N__5170),
            .I(N__5164));
    CascadeBuf I__588 (
            .O(N__5167),
            .I(N__5161));
    CascadeMux I__587 (
            .O(N__5164),
            .I(N__5158));
    CascadeMux I__586 (
            .O(N__5161),
            .I(N__5155));
    CascadeBuf I__585 (
            .O(N__5158),
            .I(N__5152));
    CascadeBuf I__584 (
            .O(N__5155),
            .I(N__5149));
    CascadeMux I__583 (
            .O(N__5152),
            .I(N__5146));
    CascadeMux I__582 (
            .O(N__5149),
            .I(N__5143));
    CascadeBuf I__581 (
            .O(N__5146),
            .I(N__5140));
    CascadeBuf I__580 (
            .O(N__5143),
            .I(N__5137));
    CascadeMux I__579 (
            .O(N__5140),
            .I(N__5134));
    CascadeMux I__578 (
            .O(N__5137),
            .I(N__5131));
    CascadeBuf I__577 (
            .O(N__5134),
            .I(N__5128));
    CascadeBuf I__576 (
            .O(N__5131),
            .I(N__5125));
    CascadeMux I__575 (
            .O(N__5128),
            .I(N__5122));
    CascadeMux I__574 (
            .O(N__5125),
            .I(N__5119));
    CascadeBuf I__573 (
            .O(N__5122),
            .I(N__5116));
    CascadeBuf I__572 (
            .O(N__5119),
            .I(N__5113));
    CascadeMux I__571 (
            .O(N__5116),
            .I(N__5110));
    CascadeMux I__570 (
            .O(N__5113),
            .I(N__5107));
    CascadeBuf I__569 (
            .O(N__5110),
            .I(N__5104));
    CascadeBuf I__568 (
            .O(N__5107),
            .I(N__5101));
    CascadeMux I__567 (
            .O(N__5104),
            .I(N__5098));
    CascadeMux I__566 (
            .O(N__5101),
            .I(N__5095));
    InMux I__565 (
            .O(N__5098),
            .I(N__5092));
    CascadeBuf I__564 (
            .O(N__5095),
            .I(N__5089));
    LocalMux I__563 (
            .O(N__5092),
            .I(N__5086));
    CascadeMux I__562 (
            .O(N__5089),
            .I(N__5083));
    Span4Mux_h I__561 (
            .O(N__5086),
            .I(N__5080));
    CascadeBuf I__560 (
            .O(N__5083),
            .I(N__5077));
    Span4Mux_h I__559 (
            .O(N__5080),
            .I(N__5074));
    CascadeMux I__558 (
            .O(N__5077),
            .I(N__5071));
    Span4Mux_h I__557 (
            .O(N__5074),
            .I(N__5068));
    InMux I__556 (
            .O(N__5071),
            .I(N__5065));
    Span4Mux_h I__555 (
            .O(N__5068),
            .I(N__5060));
    LocalMux I__554 (
            .O(N__5065),
            .I(N__5060));
    Span4Mux_h I__553 (
            .O(N__5060),
            .I(N__5057));
    IoSpan4Mux I__552 (
            .O(N__5057),
            .I(N__5054));
    Odrv4 I__551 (
            .O(N__5054),
            .I(waddr_c_2));
    InMux I__550 (
            .O(N__5051),
            .I(N__5047));
    InMux I__549 (
            .O(N__5050),
            .I(N__5044));
    LocalMux I__548 (
            .O(N__5047),
            .I(N__5041));
    LocalMux I__547 (
            .O(N__5044),
            .I(N__5037));
    Span4Mux_s2_v I__546 (
            .O(N__5041),
            .I(N__5033));
    InMux I__545 (
            .O(N__5040),
            .I(N__5030));
    Span4Mux_h I__544 (
            .O(N__5037),
            .I(N__5027));
    InMux I__543 (
            .O(N__5036),
            .I(N__5024));
    Span4Mux_v I__542 (
            .O(N__5033),
            .I(N__5019));
    LocalMux I__541 (
            .O(N__5030),
            .I(N__5019));
    Span4Mux_v I__540 (
            .O(N__5027),
            .I(N__5015));
    LocalMux I__539 (
            .O(N__5024),
            .I(N__5012));
    Span4Mux_v I__538 (
            .O(N__5019),
            .I(N__5008));
    InMux I__537 (
            .O(N__5018),
            .I(N__5005));
    Span4Mux_v I__536 (
            .O(N__5015),
            .I(N__5000));
    Span4Mux_h I__535 (
            .O(N__5012),
            .I(N__5000));
    InMux I__534 (
            .O(N__5011),
            .I(N__4997));
    Span4Mux_v I__533 (
            .O(N__5008),
            .I(N__4992));
    LocalMux I__532 (
            .O(N__5005),
            .I(N__4992));
    Span4Mux_v I__531 (
            .O(N__5000),
            .I(N__4988));
    LocalMux I__530 (
            .O(N__4997),
            .I(N__4985));
    Span4Mux_v I__529 (
            .O(N__4992),
            .I(N__4981));
    InMux I__528 (
            .O(N__4991),
            .I(N__4978));
    Span4Mux_v I__527 (
            .O(N__4988),
            .I(N__4973));
    Span4Mux_h I__526 (
            .O(N__4985),
            .I(N__4973));
    InMux I__525 (
            .O(N__4984),
            .I(N__4970));
    Span4Mux_v I__524 (
            .O(N__4981),
            .I(N__4965));
    LocalMux I__523 (
            .O(N__4978),
            .I(N__4965));
    Span4Mux_v I__522 (
            .O(N__4973),
            .I(N__4962));
    LocalMux I__521 (
            .O(N__4970),
            .I(N__4959));
    Span4Mux_v I__520 (
            .O(N__4965),
            .I(N__4956));
    Span4Mux_v I__519 (
            .O(N__4962),
            .I(N__4951));
    Span4Mux_h I__518 (
            .O(N__4959),
            .I(N__4951));
    Sp12to4 I__517 (
            .O(N__4956),
            .I(N__4948));
    Span4Mux_v I__516 (
            .O(N__4951),
            .I(N__4945));
    Span12Mux_h I__515 (
            .O(N__4948),
            .I(N__4942));
    Span4Mux_h I__514 (
            .O(N__4945),
            .I(N__4939));
    Odrv12 I__513 (
            .O(N__4942),
            .I(din_c_0));
    Odrv4 I__512 (
            .O(N__4939),
            .I(din_c_0));
    ClkMux I__511 (
            .O(N__4934),
            .I(N__4829));
    ClkMux I__510 (
            .O(N__4933),
            .I(N__4829));
    ClkMux I__509 (
            .O(N__4932),
            .I(N__4829));
    ClkMux I__508 (
            .O(N__4931),
            .I(N__4829));
    ClkMux I__507 (
            .O(N__4930),
            .I(N__4829));
    ClkMux I__506 (
            .O(N__4929),
            .I(N__4829));
    ClkMux I__505 (
            .O(N__4928),
            .I(N__4829));
    ClkMux I__504 (
            .O(N__4927),
            .I(N__4829));
    ClkMux I__503 (
            .O(N__4926),
            .I(N__4829));
    ClkMux I__502 (
            .O(N__4925),
            .I(N__4829));
    ClkMux I__501 (
            .O(N__4924),
            .I(N__4829));
    ClkMux I__500 (
            .O(N__4923),
            .I(N__4829));
    ClkMux I__499 (
            .O(N__4922),
            .I(N__4829));
    ClkMux I__498 (
            .O(N__4921),
            .I(N__4829));
    ClkMux I__497 (
            .O(N__4920),
            .I(N__4829));
    ClkMux I__496 (
            .O(N__4919),
            .I(N__4829));
    ClkMux I__495 (
            .O(N__4918),
            .I(N__4829));
    ClkMux I__494 (
            .O(N__4917),
            .I(N__4829));
    ClkMux I__493 (
            .O(N__4916),
            .I(N__4829));
    ClkMux I__492 (
            .O(N__4915),
            .I(N__4829));
    ClkMux I__491 (
            .O(N__4914),
            .I(N__4829));
    ClkMux I__490 (
            .O(N__4913),
            .I(N__4829));
    ClkMux I__489 (
            .O(N__4912),
            .I(N__4829));
    ClkMux I__488 (
            .O(N__4911),
            .I(N__4829));
    ClkMux I__487 (
            .O(N__4910),
            .I(N__4829));
    ClkMux I__486 (
            .O(N__4909),
            .I(N__4829));
    ClkMux I__485 (
            .O(N__4908),
            .I(N__4829));
    ClkMux I__484 (
            .O(N__4907),
            .I(N__4829));
    ClkMux I__483 (
            .O(N__4906),
            .I(N__4829));
    ClkMux I__482 (
            .O(N__4905),
            .I(N__4829));
    ClkMux I__481 (
            .O(N__4904),
            .I(N__4829));
    ClkMux I__480 (
            .O(N__4903),
            .I(N__4829));
    ClkMux I__479 (
            .O(N__4902),
            .I(N__4829));
    ClkMux I__478 (
            .O(N__4901),
            .I(N__4829));
    ClkMux I__477 (
            .O(N__4900),
            .I(N__4829));
    GlobalMux I__476 (
            .O(N__4829),
            .I(N__4826));
    gio2CtrlBuf I__475 (
            .O(N__4826),
            .I(rclk_c_g));
    CascadeMux I__474 (
            .O(N__4823),
            .I(N__4820));
    CascadeBuf I__473 (
            .O(N__4820),
            .I(N__4817));
    CascadeMux I__472 (
            .O(N__4817),
            .I(N__4814));
    CascadeBuf I__471 (
            .O(N__4814),
            .I(N__4811));
    CascadeMux I__470 (
            .O(N__4811),
            .I(N__4807));
    CascadeMux I__469 (
            .O(N__4810),
            .I(N__4804));
    CascadeBuf I__468 (
            .O(N__4807),
            .I(N__4801));
    CascadeBuf I__467 (
            .O(N__4804),
            .I(N__4798));
    CascadeMux I__466 (
            .O(N__4801),
            .I(N__4795));
    CascadeMux I__465 (
            .O(N__4798),
            .I(N__4792));
    CascadeBuf I__464 (
            .O(N__4795),
            .I(N__4789));
    CascadeBuf I__463 (
            .O(N__4792),
            .I(N__4786));
    CascadeMux I__462 (
            .O(N__4789),
            .I(N__4783));
    CascadeMux I__461 (
            .O(N__4786),
            .I(N__4780));
    CascadeBuf I__460 (
            .O(N__4783),
            .I(N__4777));
    CascadeBuf I__459 (
            .O(N__4780),
            .I(N__4774));
    CascadeMux I__458 (
            .O(N__4777),
            .I(N__4771));
    CascadeMux I__457 (
            .O(N__4774),
            .I(N__4768));
    CascadeBuf I__456 (
            .O(N__4771),
            .I(N__4765));
    CascadeBuf I__455 (
            .O(N__4768),
            .I(N__4762));
    CascadeMux I__454 (
            .O(N__4765),
            .I(N__4759));
    CascadeMux I__453 (
            .O(N__4762),
            .I(N__4756));
    CascadeBuf I__452 (
            .O(N__4759),
            .I(N__4753));
    CascadeBuf I__451 (
            .O(N__4756),
            .I(N__4750));
    CascadeMux I__450 (
            .O(N__4753),
            .I(N__4747));
    CascadeMux I__449 (
            .O(N__4750),
            .I(N__4744));
    CascadeBuf I__448 (
            .O(N__4747),
            .I(N__4741));
    CascadeBuf I__447 (
            .O(N__4744),
            .I(N__4738));
    CascadeMux I__446 (
            .O(N__4741),
            .I(N__4735));
    CascadeMux I__445 (
            .O(N__4738),
            .I(N__4732));
    CascadeBuf I__444 (
            .O(N__4735),
            .I(N__4729));
    CascadeBuf I__443 (
            .O(N__4732),
            .I(N__4726));
    CascadeMux I__442 (
            .O(N__4729),
            .I(N__4723));
    CascadeMux I__441 (
            .O(N__4726),
            .I(N__4720));
    CascadeBuf I__440 (
            .O(N__4723),
            .I(N__4717));
    CascadeBuf I__439 (
            .O(N__4720),
            .I(N__4714));
    CascadeMux I__438 (
            .O(N__4717),
            .I(N__4711));
    CascadeMux I__437 (
            .O(N__4714),
            .I(N__4708));
    CascadeBuf I__436 (
            .O(N__4711),
            .I(N__4705));
    CascadeBuf I__435 (
            .O(N__4708),
            .I(N__4702));
    CascadeMux I__434 (
            .O(N__4705),
            .I(N__4699));
    CascadeMux I__433 (
            .O(N__4702),
            .I(N__4696));
    CascadeBuf I__432 (
            .O(N__4699),
            .I(N__4693));
    CascadeBuf I__431 (
            .O(N__4696),
            .I(N__4690));
    CascadeMux I__430 (
            .O(N__4693),
            .I(N__4687));
    CascadeMux I__429 (
            .O(N__4690),
            .I(N__4684));
    CascadeBuf I__428 (
            .O(N__4687),
            .I(N__4681));
    CascadeBuf I__427 (
            .O(N__4684),
            .I(N__4678));
    CascadeMux I__426 (
            .O(N__4681),
            .I(N__4675));
    CascadeMux I__425 (
            .O(N__4678),
            .I(N__4672));
    CascadeBuf I__424 (
            .O(N__4675),
            .I(N__4669));
    CascadeBuf I__423 (
            .O(N__4672),
            .I(N__4666));
    CascadeMux I__422 (
            .O(N__4669),
            .I(N__4663));
    CascadeMux I__421 (
            .O(N__4666),
            .I(N__4660));
    CascadeBuf I__420 (
            .O(N__4663),
            .I(N__4657));
    CascadeBuf I__419 (
            .O(N__4660),
            .I(N__4654));
    CascadeMux I__418 (
            .O(N__4657),
            .I(N__4651));
    CascadeMux I__417 (
            .O(N__4654),
            .I(N__4648));
    InMux I__416 (
            .O(N__4651),
            .I(N__4645));
    CascadeBuf I__415 (
            .O(N__4648),
            .I(N__4642));
    LocalMux I__414 (
            .O(N__4645),
            .I(N__4639));
    CascadeMux I__413 (
            .O(N__4642),
            .I(N__4636));
    Span4Mux_s2_v I__412 (
            .O(N__4639),
            .I(N__4633));
    CascadeBuf I__411 (
            .O(N__4636),
            .I(N__4630));
    Span4Mux_h I__410 (
            .O(N__4633),
            .I(N__4627));
    CascadeMux I__409 (
            .O(N__4630),
            .I(N__4624));
    Span4Mux_v I__408 (
            .O(N__4627),
            .I(N__4621));
    InMux I__407 (
            .O(N__4624),
            .I(N__4618));
    Span4Mux_v I__406 (
            .O(N__4621),
            .I(N__4615));
    LocalMux I__405 (
            .O(N__4618),
            .I(N__4612));
    Sp12to4 I__404 (
            .O(N__4615),
            .I(N__4609));
    Sp12to4 I__403 (
            .O(N__4612),
            .I(N__4606));
    Span12Mux_h I__402 (
            .O(N__4609),
            .I(N__4601));
    Span12Mux_s10_v I__401 (
            .O(N__4606),
            .I(N__4601));
    Odrv12 I__400 (
            .O(N__4601),
            .I(raddr_c_3));
    CascadeMux I__399 (
            .O(N__4598),
            .I(N__4595));
    CascadeBuf I__398 (
            .O(N__4595),
            .I(N__4592));
    CascadeMux I__397 (
            .O(N__4592),
            .I(N__4589));
    CascadeBuf I__396 (
            .O(N__4589),
            .I(N__4586));
    CascadeMux I__395 (
            .O(N__4586),
            .I(N__4582));
    CascadeMux I__394 (
            .O(N__4585),
            .I(N__4579));
    CascadeBuf I__393 (
            .O(N__4582),
            .I(N__4576));
    CascadeBuf I__392 (
            .O(N__4579),
            .I(N__4573));
    CascadeMux I__391 (
            .O(N__4576),
            .I(N__4570));
    CascadeMux I__390 (
            .O(N__4573),
            .I(N__4567));
    CascadeBuf I__389 (
            .O(N__4570),
            .I(N__4564));
    CascadeBuf I__388 (
            .O(N__4567),
            .I(N__4561));
    CascadeMux I__387 (
            .O(N__4564),
            .I(N__4558));
    CascadeMux I__386 (
            .O(N__4561),
            .I(N__4555));
    CascadeBuf I__385 (
            .O(N__4558),
            .I(N__4552));
    CascadeBuf I__384 (
            .O(N__4555),
            .I(N__4549));
    CascadeMux I__383 (
            .O(N__4552),
            .I(N__4546));
    CascadeMux I__382 (
            .O(N__4549),
            .I(N__4543));
    CascadeBuf I__381 (
            .O(N__4546),
            .I(N__4540));
    CascadeBuf I__380 (
            .O(N__4543),
            .I(N__4537));
    CascadeMux I__379 (
            .O(N__4540),
            .I(N__4534));
    CascadeMux I__378 (
            .O(N__4537),
            .I(N__4531));
    CascadeBuf I__377 (
            .O(N__4534),
            .I(N__4528));
    CascadeBuf I__376 (
            .O(N__4531),
            .I(N__4525));
    CascadeMux I__375 (
            .O(N__4528),
            .I(N__4522));
    CascadeMux I__374 (
            .O(N__4525),
            .I(N__4519));
    CascadeBuf I__373 (
            .O(N__4522),
            .I(N__4516));
    CascadeBuf I__372 (
            .O(N__4519),
            .I(N__4513));
    CascadeMux I__371 (
            .O(N__4516),
            .I(N__4510));
    CascadeMux I__370 (
            .O(N__4513),
            .I(N__4507));
    CascadeBuf I__369 (
            .O(N__4510),
            .I(N__4504));
    CascadeBuf I__368 (
            .O(N__4507),
            .I(N__4501));
    CascadeMux I__367 (
            .O(N__4504),
            .I(N__4498));
    CascadeMux I__366 (
            .O(N__4501),
            .I(N__4495));
    CascadeBuf I__365 (
            .O(N__4498),
            .I(N__4492));
    CascadeBuf I__364 (
            .O(N__4495),
            .I(N__4489));
    CascadeMux I__363 (
            .O(N__4492),
            .I(N__4486));
    CascadeMux I__362 (
            .O(N__4489),
            .I(N__4483));
    CascadeBuf I__361 (
            .O(N__4486),
            .I(N__4480));
    CascadeBuf I__360 (
            .O(N__4483),
            .I(N__4477));
    CascadeMux I__359 (
            .O(N__4480),
            .I(N__4474));
    CascadeMux I__358 (
            .O(N__4477),
            .I(N__4471));
    CascadeBuf I__357 (
            .O(N__4474),
            .I(N__4468));
    CascadeBuf I__356 (
            .O(N__4471),
            .I(N__4465));
    CascadeMux I__355 (
            .O(N__4468),
            .I(N__4462));
    CascadeMux I__354 (
            .O(N__4465),
            .I(N__4459));
    CascadeBuf I__353 (
            .O(N__4462),
            .I(N__4456));
    CascadeBuf I__352 (
            .O(N__4459),
            .I(N__4453));
    CascadeMux I__351 (
            .O(N__4456),
            .I(N__4450));
    CascadeMux I__350 (
            .O(N__4453),
            .I(N__4447));
    CascadeBuf I__349 (
            .O(N__4450),
            .I(N__4444));
    CascadeBuf I__348 (
            .O(N__4447),
            .I(N__4441));
    CascadeMux I__347 (
            .O(N__4444),
            .I(N__4438));
    CascadeMux I__346 (
            .O(N__4441),
            .I(N__4435));
    CascadeBuf I__345 (
            .O(N__4438),
            .I(N__4432));
    CascadeBuf I__344 (
            .O(N__4435),
            .I(N__4429));
    CascadeMux I__343 (
            .O(N__4432),
            .I(N__4426));
    CascadeMux I__342 (
            .O(N__4429),
            .I(N__4423));
    InMux I__341 (
            .O(N__4426),
            .I(N__4420));
    CascadeBuf I__340 (
            .O(N__4423),
            .I(N__4417));
    LocalMux I__339 (
            .O(N__4420),
            .I(N__4414));
    CascadeMux I__338 (
            .O(N__4417),
            .I(N__4411));
    IoSpan4Mux I__337 (
            .O(N__4414),
            .I(N__4408));
    CascadeBuf I__336 (
            .O(N__4411),
            .I(N__4405));
    IoSpan4Mux I__335 (
            .O(N__4408),
            .I(N__4402));
    CascadeMux I__334 (
            .O(N__4405),
            .I(N__4399));
    IoSpan4Mux I__333 (
            .O(N__4402),
            .I(N__4396));
    InMux I__332 (
            .O(N__4399),
            .I(N__4393));
    IoSpan4Mux I__331 (
            .O(N__4396),
            .I(N__4390));
    LocalMux I__330 (
            .O(N__4393),
            .I(N__4387));
    IoSpan4Mux I__329 (
            .O(N__4390),
            .I(N__4382));
    IoSpan4Mux I__328 (
            .O(N__4387),
            .I(N__4382));
    IoSpan4Mux I__327 (
            .O(N__4382),
            .I(N__4379));
    Odrv4 I__326 (
            .O(N__4379),
            .I(waddr_c_1));
    InMux I__325 (
            .O(N__4376),
            .I(N__4373));
    LocalMux I__324 (
            .O(N__4373),
            .I(N__4369));
    InMux I__323 (
            .O(N__4372),
            .I(N__4365));
    Span4Mux_v I__322 (
            .O(N__4369),
            .I(N__4362));
    InMux I__321 (
            .O(N__4368),
            .I(N__4359));
    LocalMux I__320 (
            .O(N__4365),
            .I(N__4356));
    Span4Mux_v I__319 (
            .O(N__4362),
            .I(N__4350));
    LocalMux I__318 (
            .O(N__4359),
            .I(N__4350));
    Span4Mux_h I__317 (
            .O(N__4356),
            .I(N__4346));
    InMux I__316 (
            .O(N__4355),
            .I(N__4343));
    Span4Mux_v I__315 (
            .O(N__4350),
            .I(N__4340));
    InMux I__314 (
            .O(N__4349),
            .I(N__4337));
    Span4Mux_v I__313 (
            .O(N__4346),
            .I(N__4334));
    LocalMux I__312 (
            .O(N__4343),
            .I(N__4331));
    Span4Mux_v I__311 (
            .O(N__4340),
            .I(N__4325));
    LocalMux I__310 (
            .O(N__4337),
            .I(N__4325));
    Span4Mux_v I__309 (
            .O(N__4334),
            .I(N__4319));
    Span4Mux_h I__308 (
            .O(N__4331),
            .I(N__4319));
    InMux I__307 (
            .O(N__4330),
            .I(N__4316));
    Span4Mux_v I__306 (
            .O(N__4325),
            .I(N__4313));
    InMux I__305 (
            .O(N__4324),
            .I(N__4310));
    Span4Mux_v I__304 (
            .O(N__4319),
            .I(N__4307));
    LocalMux I__303 (
            .O(N__4316),
            .I(N__4304));
    Span4Mux_v I__302 (
            .O(N__4313),
            .I(N__4298));
    LocalMux I__301 (
            .O(N__4310),
            .I(N__4298));
    Span4Mux_v I__300 (
            .O(N__4307),
            .I(N__4293));
    Span4Mux_h I__299 (
            .O(N__4304),
            .I(N__4293));
    InMux I__298 (
            .O(N__4303),
            .I(N__4290));
    Span4Mux_v I__297 (
            .O(N__4298),
            .I(N__4287));
    Span4Mux_v I__296 (
            .O(N__4293),
            .I(N__4284));
    LocalMux I__295 (
            .O(N__4290),
            .I(N__4281));
    Sp12to4 I__294 (
            .O(N__4287),
            .I(N__4278));
    Span4Mux_v I__293 (
            .O(N__4284),
            .I(N__4273));
    Span4Mux_h I__292 (
            .O(N__4281),
            .I(N__4273));
    Span12Mux_h I__291 (
            .O(N__4278),
            .I(N__4270));
    IoSpan4Mux I__290 (
            .O(N__4273),
            .I(N__4267));
    Odrv12 I__289 (
            .O(N__4270),
            .I(din_c_4));
    Odrv4 I__288 (
            .O(N__4267),
            .I(din_c_4));
    InMux I__287 (
            .O(N__4262),
            .I(N__4258));
    InMux I__286 (
            .O(N__4261),
            .I(N__4255));
    LocalMux I__285 (
            .O(N__4258),
            .I(N__4252));
    LocalMux I__284 (
            .O(N__4255),
            .I(N__4248));
    Span4Mux_v I__283 (
            .O(N__4252),
            .I(N__4244));
    InMux I__282 (
            .O(N__4251),
            .I(N__4241));
    Span4Mux_v I__281 (
            .O(N__4248),
            .I(N__4237));
    InMux I__280 (
            .O(N__4247),
            .I(N__4234));
    Span4Mux_v I__279 (
            .O(N__4244),
            .I(N__4229));
    LocalMux I__278 (
            .O(N__4241),
            .I(N__4229));
    InMux I__277 (
            .O(N__4240),
            .I(N__4225));
    Span4Mux_v I__276 (
            .O(N__4237),
            .I(N__4220));
    LocalMux I__275 (
            .O(N__4234),
            .I(N__4220));
    Span4Mux_v I__274 (
            .O(N__4229),
            .I(N__4216));
    InMux I__273 (
            .O(N__4228),
            .I(N__4213));
    LocalMux I__272 (
            .O(N__4225),
            .I(N__4210));
    Span4Mux_v I__271 (
            .O(N__4220),
            .I(N__4207));
    InMux I__270 (
            .O(N__4219),
            .I(N__4204));
    Span4Mux_v I__269 (
            .O(N__4216),
            .I(N__4199));
    LocalMux I__268 (
            .O(N__4213),
            .I(N__4199));
    Span4Mux_s1_v I__267 (
            .O(N__4210),
            .I(N__4196));
    Span4Mux_v I__266 (
            .O(N__4207),
            .I(N__4191));
    LocalMux I__265 (
            .O(N__4204),
            .I(N__4191));
    Span4Mux_v I__264 (
            .O(N__4199),
            .I(N__4185));
    Span4Mux_v I__263 (
            .O(N__4196),
            .I(N__4185));
    Span4Mux_v I__262 (
            .O(N__4191),
            .I(N__4182));
    InMux I__261 (
            .O(N__4190),
            .I(N__4179));
    Sp12to4 I__260 (
            .O(N__4185),
            .I(N__4176));
    Span4Mux_v I__259 (
            .O(N__4182),
            .I(N__4171));
    LocalMux I__258 (
            .O(N__4179),
            .I(N__4171));
    Span12Mux_h I__257 (
            .O(N__4176),
            .I(N__4168));
    IoSpan4Mux I__256 (
            .O(N__4171),
            .I(N__4165));
    Span12Mux_h I__255 (
            .O(N__4168),
            .I(N__4162));
    IoSpan4Mux I__254 (
            .O(N__4165),
            .I(N__4159));
    Odrv12 I__253 (
            .O(N__4162),
            .I(din_c_6));
    Odrv4 I__252 (
            .O(N__4159),
            .I(din_c_6));
    InMux I__251 (
            .O(N__4154),
            .I(N__4151));
    LocalMux I__250 (
            .O(N__4151),
            .I(N__4148));
    Span4Mux_v I__249 (
            .O(N__4148),
            .I(N__4141));
    InMux I__248 (
            .O(N__4147),
            .I(N__4138));
    InMux I__247 (
            .O(N__4146),
            .I(N__4135));
    InMux I__246 (
            .O(N__4145),
            .I(N__4132));
    InMux I__245 (
            .O(N__4144),
            .I(N__4128));
    Span4Mux_v I__244 (
            .O(N__4141),
            .I(N__4123));
    LocalMux I__243 (
            .O(N__4138),
            .I(N__4123));
    LocalMux I__242 (
            .O(N__4135),
            .I(N__4119));
    LocalMux I__241 (
            .O(N__4132),
            .I(N__4116));
    InMux I__240 (
            .O(N__4131),
            .I(N__4113));
    LocalMux I__239 (
            .O(N__4128),
            .I(N__4110));
    Span4Mux_v I__238 (
            .O(N__4123),
            .I(N__4107));
    InMux I__237 (
            .O(N__4122),
            .I(N__4104));
    Span12Mux_v I__236 (
            .O(N__4119),
            .I(N__4100));
    Sp12to4 I__235 (
            .O(N__4116),
            .I(N__4095));
    LocalMux I__234 (
            .O(N__4113),
            .I(N__4095));
    Sp12to4 I__233 (
            .O(N__4110),
            .I(N__4092));
    Span4Mux_v I__232 (
            .O(N__4107),
            .I(N__4087));
    LocalMux I__231 (
            .O(N__4104),
            .I(N__4087));
    InMux I__230 (
            .O(N__4103),
            .I(N__4084));
    Span12Mux_h I__229 (
            .O(N__4100),
            .I(N__4081));
    Span12Mux_v I__228 (
            .O(N__4095),
            .I(N__4076));
    Span12Mux_s4_v I__227 (
            .O(N__4092),
            .I(N__4076));
    Span4Mux_v I__226 (
            .O(N__4087),
            .I(N__4073));
    LocalMux I__225 (
            .O(N__4084),
            .I(N__4070));
    Span12Mux_h I__224 (
            .O(N__4081),
            .I(N__4067));
    Span12Mux_h I__223 (
            .O(N__4076),
            .I(N__4064));
    Span4Mux_v I__222 (
            .O(N__4073),
            .I(N__4059));
    Span4Mux_v I__221 (
            .O(N__4070),
            .I(N__4059));
    Span12Mux_v I__220 (
            .O(N__4067),
            .I(N__4054));
    Span12Mux_h I__219 (
            .O(N__4064),
            .I(N__4054));
    Span4Mux_h I__218 (
            .O(N__4059),
            .I(N__4051));
    Odrv12 I__217 (
            .O(N__4054),
            .I(din_c_7));
    Odrv4 I__216 (
            .O(N__4051),
            .I(din_c_7));
    InMux I__215 (
            .O(N__4046),
            .I(N__4043));
    LocalMux I__214 (
            .O(N__4043),
            .I(N__4040));
    Span4Mux_v I__213 (
            .O(N__4040),
            .I(N__4036));
    InMux I__212 (
            .O(N__4039),
            .I(N__4033));
    Span4Mux_v I__211 (
            .O(N__4036),
            .I(N__4028));
    LocalMux I__210 (
            .O(N__4033),
            .I(N__4028));
    Span4Mux_v I__209 (
            .O(N__4028),
            .I(N__4024));
    InMux I__208 (
            .O(N__4027),
            .I(N__4021));
    Span4Mux_v I__207 (
            .O(N__4024),
            .I(N__4016));
    LocalMux I__206 (
            .O(N__4021),
            .I(N__4016));
    Span4Mux_v I__205 (
            .O(N__4016),
            .I(N__4011));
    InMux I__204 (
            .O(N__4015),
            .I(N__4008));
    InMux I__203 (
            .O(N__4014),
            .I(N__4004));
    Span4Mux_v I__202 (
            .O(N__4011),
            .I(N__3999));
    LocalMux I__201 (
            .O(N__4008),
            .I(N__3999));
    InMux I__200 (
            .O(N__4007),
            .I(N__3995));
    LocalMux I__199 (
            .O(N__4004),
            .I(N__3992));
    Span4Mux_v I__198 (
            .O(N__3999),
            .I(N__3989));
    InMux I__197 (
            .O(N__3998),
            .I(N__3986));
    LocalMux I__196 (
            .O(N__3995),
            .I(N__3983));
    Sp12to4 I__195 (
            .O(N__3992),
            .I(N__3979));
    Span4Mux_h I__194 (
            .O(N__3989),
            .I(N__3976));
    LocalMux I__193 (
            .O(N__3986),
            .I(N__3973));
    Span4Mux_v I__192 (
            .O(N__3983),
            .I(N__3970));
    InMux I__191 (
            .O(N__3982),
            .I(N__3967));
    Span12Mux_v I__190 (
            .O(N__3979),
            .I(N__3964));
    Sp12to4 I__189 (
            .O(N__3976),
            .I(N__3961));
    Sp12to4 I__188 (
            .O(N__3973),
            .I(N__3958));
    Span4Mux_v I__187 (
            .O(N__3970),
            .I(N__3953));
    LocalMux I__186 (
            .O(N__3967),
            .I(N__3953));
    Span12Mux_v I__185 (
            .O(N__3964),
            .I(N__3950));
    Span12Mux_h I__184 (
            .O(N__3961),
            .I(N__3947));
    Span12Mux_v I__183 (
            .O(N__3958),
            .I(N__3944));
    Span4Mux_v I__182 (
            .O(N__3953),
            .I(N__3941));
    Odrv12 I__181 (
            .O(N__3950),
            .I(din_c_3));
    Odrv12 I__180 (
            .O(N__3947),
            .I(din_c_3));
    Odrv12 I__179 (
            .O(N__3944),
            .I(din_c_3));
    Odrv4 I__178 (
            .O(N__3941),
            .I(din_c_3));
    InMux I__177 (
            .O(N__3932),
            .I(N__3929));
    LocalMux I__176 (
            .O(N__3929),
            .I(N__3926));
    Span4Mux_v I__175 (
            .O(N__3926),
            .I(N__3922));
    InMux I__174 (
            .O(N__3925),
            .I(N__3919));
    Span4Mux_v I__173 (
            .O(N__3922),
            .I(N__3914));
    LocalMux I__172 (
            .O(N__3919),
            .I(N__3914));
    Span4Mux_v I__171 (
            .O(N__3914),
            .I(N__3910));
    InMux I__170 (
            .O(N__3913),
            .I(N__3907));
    Span4Mux_v I__169 (
            .O(N__3910),
            .I(N__3901));
    LocalMux I__168 (
            .O(N__3907),
            .I(N__3901));
    InMux I__167 (
            .O(N__3906),
            .I(N__3898));
    Span4Mux_v I__166 (
            .O(N__3901),
            .I(N__3895));
    LocalMux I__165 (
            .O(N__3898),
            .I(N__3892));
    Span4Mux_v I__164 (
            .O(N__3895),
            .I(N__3885));
    Span4Mux_v I__163 (
            .O(N__3892),
            .I(N__3885));
    InMux I__162 (
            .O(N__3891),
            .I(N__3882));
    InMux I__161 (
            .O(N__3890),
            .I(N__3878));
    Span4Mux_h I__160 (
            .O(N__3885),
            .I(N__3875));
    LocalMux I__159 (
            .O(N__3882),
            .I(N__3872));
    InMux I__158 (
            .O(N__3881),
            .I(N__3869));
    LocalMux I__157 (
            .O(N__3878),
            .I(N__3865));
    Sp12to4 I__156 (
            .O(N__3875),
            .I(N__3862));
    Span12Mux_v I__155 (
            .O(N__3872),
            .I(N__3857));
    LocalMux I__154 (
            .O(N__3869),
            .I(N__3857));
    InMux I__153 (
            .O(N__3868),
            .I(N__3854));
    Span12Mux_v I__152 (
            .O(N__3865),
            .I(N__3851));
    Span12Mux_h I__151 (
            .O(N__3862),
            .I(N__3844));
    Span12Mux_v I__150 (
            .O(N__3857),
            .I(N__3844));
    LocalMux I__149 (
            .O(N__3854),
            .I(N__3844));
    Odrv12 I__148 (
            .O(N__3851),
            .I(din_c_2));
    Odrv12 I__147 (
            .O(N__3844),
            .I(din_c_2));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam waddr_ibuf_RNIO66O1_0_11_LC_7_17_0.C_ON=1'b0;
    defparam waddr_ibuf_RNIO66O1_0_11_LC_7_17_0.SEQ_MODE=4'b0000;
    defparam waddr_ibuf_RNIO66O1_0_11_LC_7_17_0.LUT_INIT=16'b0000000010000000;
    LogicCell40 waddr_ibuf_RNIO66O1_0_11_LC_7_17_0 (
            .in0(N__10057),
            .in1(N__10093),
            .in2(N__9977),
            .in3(N__10009),
            .lcout(mem_WE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam waddr_ibuf_RNIO66O1_11_LC_7_17_1.C_ON=1'b0;
    defparam waddr_ibuf_RNIO66O1_11_LC_7_17_1.SEQ_MODE=4'b0000;
    defparam waddr_ibuf_RNIO66O1_11_LC_7_17_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 waddr_ibuf_RNIO66O1_11_LC_7_17_1 (
            .in0(N__10094),
            .in1(N__10058),
            .in2(N__10025),
            .in3(N__9964),
            .lcout(mem_WE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam waddr_ibuf_RNIO66O1_1_11_LC_7_17_2.C_ON=1'b0;
    defparam waddr_ibuf_RNIO66O1_1_11_LC_7_17_2.SEQ_MODE=4'b0000;
    defparam waddr_ibuf_RNIO66O1_1_11_LC_7_17_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 waddr_ibuf_RNIO66O1_1_11_LC_7_17_2 (
            .in0(N__10059),
            .in1(N__10095),
            .in2(N__9978),
            .in3(N__10013),
            .lcout(mem_WE_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam waddr_ibuf_RNIO66O1_2_11_LC_7_17_3.C_ON=1'b0;
    defparam waddr_ibuf_RNIO66O1_2_11_LC_7_17_3.SEQ_MODE=4'b0000;
    defparam waddr_ibuf_RNIO66O1_2_11_LC_7_17_3.LUT_INIT=16'b0000000000001000;
    LogicCell40 waddr_ibuf_RNIO66O1_2_11_LC_7_17_3 (
            .in0(N__10096),
            .in1(N__10060),
            .in2(N__10026),
            .in3(N__9968),
            .lcout(mem_WE_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam waddr_ibuf_RNIO66O1_3_11_LC_7_17_4.C_ON=1'b0;
    defparam waddr_ibuf_RNIO66O1_3_11_LC_7_17_4.SEQ_MODE=4'b0000;
    defparam waddr_ibuf_RNIO66O1_3_11_LC_7_17_4.LUT_INIT=16'b0100000000000000;
    LogicCell40 waddr_ibuf_RNIO66O1_3_11_LC_7_17_4 (
            .in0(N__10061),
            .in1(N__10097),
            .in2(N__9979),
            .in3(N__10017),
            .lcout(mem_WE_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam waddr_ibuf_RNIO66O1_4_11_LC_7_17_5.C_ON=1'b0;
    defparam waddr_ibuf_RNIO66O1_4_11_LC_7_17_5.SEQ_MODE=4'b0000;
    defparam waddr_ibuf_RNIO66O1_4_11_LC_7_17_5.LUT_INIT=16'b0000001000000000;
    LogicCell40 waddr_ibuf_RNIO66O1_4_11_LC_7_17_5 (
            .in0(N__10098),
            .in1(N__10062),
            .in2(N__10027),
            .in3(N__9972),
            .lcout(mem_WE_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam waddr_ibuf_RNIO66O1_5_11_LC_7_17_6.C_ON=1'b0;
    defparam waddr_ibuf_RNIO66O1_5_11_LC_7_17_6.SEQ_MODE=4'b0000;
    defparam waddr_ibuf_RNIO66O1_5_11_LC_7_17_6.LUT_INIT=16'b0000010000000000;
    LogicCell40 waddr_ibuf_RNIO66O1_5_11_LC_7_17_6 (
            .in0(N__10063),
            .in1(N__10099),
            .in2(N__9980),
            .in3(N__10021),
            .lcout(mem_WE_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam waddr_ibuf_RNIO66O1_6_11_LC_7_17_7.C_ON=1'b0;
    defparam waddr_ibuf_RNIO66O1_6_11_LC_7_17_7.SEQ_MODE=4'b0000;
    defparam waddr_ibuf_RNIO66O1_6_11_LC_7_17_7.LUT_INIT=16'b0000000000000010;
    LogicCell40 waddr_ibuf_RNIO66O1_6_11_LC_7_17_7 (
            .in0(N__10100),
            .in1(N__10064),
            .in2(N__10028),
            .in3(N__9976),
            .lcout(mem_WE_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_0_LC_10_1_4.C_ON=1'b0;
    defparam dout_obuf_RNO_4_0_LC_10_1_4.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_0_LC_10_1_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_4_0_LC_10_1_4 (
            .in0(N__9896),
            .in1(N__12430),
            .in2(_gnd_net_),
            .in3(N__9878),
            .lcout(dout_obuf_RNO_4Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_1_LC_10_1_6.C_ON=1'b0;
    defparam dout_obuf_RNO_4_1_LC_10_1_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_1_LC_10_1_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_4_1_LC_10_1_6 (
            .in0(N__9866),
            .in1(N__12431),
            .in2(_gnd_net_),
            .in3(N__9851),
            .lcout(dout_obuf_RNO_4Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_7_LC_10_7_1.C_ON=1'b0;
    defparam dout_obuf_RNO_4_7_LC_10_7_1.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_7_LC_10_7_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 dout_obuf_RNO_4_7_LC_10_7_1 (
            .in0(N__9842),
            .in1(_gnd_net_),
            .in2(N__12364),
            .in3(N__9833),
            .lcout(dout_obuf_RNO_4Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_6_LC_10_7_6.C_ON=1'b0;
    defparam dout_obuf_RNO_4_6_LC_10_7_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_6_LC_10_7_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_4_6_LC_10_7_6 (
            .in0(N__11030),
            .in1(N__12345),
            .in2(_gnd_net_),
            .in3(N__11012),
            .lcout(dout_obuf_RNO_4Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_9_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_9_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_9_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_1_LC_10_9_3.C_ON=1'b0;
    defparam dout_obuf_RNO_2_1_LC_10_9_3.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_1_LC_10_9_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_2_1_LC_10_9_3 (
            .in0(N__10439),
            .in1(N__12414),
            .in2(_gnd_net_),
            .in3(N__10430),
            .lcout(dout_obuf_RNO_2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_0_LC_10_9_7.C_ON=1'b0;
    defparam dout_obuf_RNO_2_0_LC_10_9_7.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_0_LC_10_9_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_2_0_LC_10_9_7 (
            .in0(N__10415),
            .in1(N__12413),
            .in2(_gnd_net_),
            .in3(N__10403),
            .lcout(dout_obuf_RNO_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_1_LC_10_10_5.C_ON=1'b0;
    defparam dout_obuf_RNO_1_1_LC_10_10_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_1_LC_10_10_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_1_1_LC_10_10_5 (
            .in0(N__11414),
            .in1(N__12755),
            .in2(_gnd_net_),
            .in3(N__10385),
            .lcout(),
            .ltout(mem_N_162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_LC_10_10_6.C_ON=1'b0;
    defparam dout_obuf_RNO_1_LC_10_10_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_LC_10_10_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 dout_obuf_RNO_1_LC_10_10_6 (
            .in0(N__11162),
            .in1(_gnd_net_),
            .in2(N__10373),
            .in3(N__12584),
            .lcout(dout_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_0_LC_10_11_2.C_ON=1'b0;
    defparam dout_obuf_RNO_1_0_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_0_LC_10_11_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_1_0_LC_10_11_2 (
            .in0(N__12751),
            .in1(N__11372),
            .in2(_gnd_net_),
            .in3(N__10358),
            .lcout(),
            .ltout(mem_N_156_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_LC_10_11_3.C_ON=1'b0;
    defparam dout_obuf_RNO_0_LC_10_11_3.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_LC_10_11_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 dout_obuf_RNO_0_LC_10_11_3 (
            .in0(_gnd_net_),
            .in1(N__12559),
            .in2(N__10346),
            .in3(N__11147),
            .lcout(dout_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_1_LC_10_11_5.C_ON=1'b0;
    defparam dout_obuf_RNO_0_1_LC_10_11_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_1_LC_10_11_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_0_1_LC_10_11_5 (
            .in0(N__12011),
            .in1(N__12750),
            .in2(_gnd_net_),
            .in3(N__11171),
            .lcout(mem_N_160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_0_LC_10_11_6.C_ON=1'b0;
    defparam dout_obuf_RNO_0_0_LC_10_11_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_0_LC_10_11_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_0_0_LC_10_11_6 (
            .in0(N__11156),
            .in1(N__12749),
            .in2(_gnd_net_),
            .in3(N__11303),
            .lcout(mem_N_154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_2_LC_10_11_7.C_ON=1'b0;
    defparam dout_obuf_RNO_2_2_LC_10_11_7.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_2_LC_10_11_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_2_2_LC_10_11_7 (
            .in0(N__11141),
            .in1(N__12328),
            .in2(_gnd_net_),
            .in3(N__11129),
            .lcout(dout_obuf_RNO_2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_2_LC_10_12_5.C_ON=1'b0;
    defparam dout_obuf_RNO_0_2_LC_10_12_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_2_LC_10_12_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_0_2_LC_10_12_5 (
            .in0(N__11261),
            .in1(N__12730),
            .in2(_gnd_net_),
            .in3(N__11111),
            .lcout(),
            .ltout(mem_N_166_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_LC_10_12_6.C_ON=1'b0;
    defparam dout_obuf_RNO_2_LC_10_12_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_LC_10_12_6.LUT_INIT=16'b1111001111000000;
    LogicCell40 dout_obuf_RNO_2_LC_10_12_6 (
            .in0(_gnd_net_),
            .in1(N__12580),
            .in2(N__11105),
            .in3(N__11795),
            .lcout(dout_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_7_LC_10_15_0.C_ON=1'b0;
    defparam dout_obuf_RNO_1_7_LC_10_15_0.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_7_LC_10_15_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_1_7_LC_10_15_0 (
            .in0(N__12715),
            .in1(N__12047),
            .in2(_gnd_net_),
            .in3(N__11093),
            .lcout(mem_N_150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_7_LC_10_15_3.C_ON=1'b0;
    defparam dout_obuf_RNO_2_7_LC_10_15_3.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_7_LC_10_15_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_2_7_LC_10_15_3 (
            .in0(N__11084),
            .in1(N__12321),
            .in2(_gnd_net_),
            .in3(N__11075),
            .lcout(),
            .ltout(dout_obuf_RNO_2Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_7_LC_10_15_4.C_ON=1'b0;
    defparam dout_obuf_RNO_0_7_LC_10_15_4.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_7_LC_10_15_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 dout_obuf_RNO_0_7_LC_10_15_4 (
            .in0(_gnd_net_),
            .in1(N__12714),
            .in2(N__11060),
            .in3(N__11924),
            .lcout(),
            .ltout(mem_N_149_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_7_LC_10_15_5.C_ON=1'b0;
    defparam dout_obuf_RNO_7_LC_10_15_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_7_LC_10_15_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 dout_obuf_RNO_7_LC_10_15_5 (
            .in0(N__11057),
            .in1(_gnd_net_),
            .in2(N__11051),
            .in3(N__12560),
            .lcout(dout_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_1_LC_10_17_2.C_ON=1'b0;
    defparam dout_obuf_RNO_5_1_LC_10_17_2.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_1_LC_10_17_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 dout_obuf_RNO_5_1_LC_10_17_2 (
            .in0(N__11438),
            .in1(_gnd_net_),
            .in2(N__12400),
            .in3(N__11423),
            .lcout(dout_obuf_RNO_5Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_0_LC_10_17_3.C_ON=1'b0;
    defparam dout_obuf_RNO_5_0_LC_10_17_3.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_0_LC_10_17_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_5_0_LC_10_17_3 (
            .in0(N__11402),
            .in1(N__12384),
            .in2(_gnd_net_),
            .in3(N__11390),
            .lcout(dout_obuf_RNO_5Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_3_LC_10_17_6.C_ON=1'b0;
    defparam dout_obuf_RNO_5_3_LC_10_17_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_3_LC_10_17_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 dout_obuf_RNO_5_3_LC_10_17_6 (
            .in0(N__11363),
            .in1(_gnd_net_),
            .in2(N__12401),
            .in3(N__11351),
            .lcout(dout_obuf_RNO_5Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_0_LC_10_25_5.C_ON=1'b0;
    defparam dout_obuf_RNO_3_0_LC_10_25_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_0_LC_10_25_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_3_0_LC_10_25_5 (
            .in0(N__11333),
            .in1(N__12358),
            .in2(_gnd_net_),
            .in3(N__11321),
            .lcout(dout_obuf_RNO_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_2_LC_10_27_3.C_ON=1'b0;
    defparam dout_obuf_RNO_3_2_LC_10_27_3.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_2_LC_10_27_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_3_2_LC_10_27_3 (
            .in0(N__11291),
            .in1(N__12278),
            .in2(_gnd_net_),
            .in3(N__11279),
            .lcout(dout_obuf_RNO_3Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_3_LC_10_27_7.C_ON=1'b0;
    defparam dout_obuf_RNO_3_3_LC_10_27_7.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_3_LC_10_27_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_3_3_LC_10_27_7 (
            .in0(N__11246),
            .in1(N__12279),
            .in2(_gnd_net_),
            .in3(N__11237),
            .lcout(dout_obuf_RNO_3Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_2_LC_11_3_5.C_ON=1'b0;
    defparam dout_obuf_RNO_4_2_LC_11_3_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_2_LC_11_3_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_4_2_LC_11_3_5 (
            .in0(N__11222),
            .in1(N__12349),
            .in2(_gnd_net_),
            .in3(N__11210),
            .lcout(dout_obuf_RNO_4Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_3_LC_11_3_7.C_ON=1'b0;
    defparam dout_obuf_RNO_4_3_LC_11_3_7.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_3_LC_11_3_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_4_3_LC_11_3_7 (
            .in0(N__11192),
            .in1(N__12350),
            .in2(_gnd_net_),
            .in3(N__11183),
            .lcout(dout_obuf_RNO_4Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_5_LC_11_5_0.C_ON=1'b0;
    defparam dout_obuf_RNO_4_5_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_5_LC_11_5_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_4_5_LC_11_5_0 (
            .in0(N__11618),
            .in1(N__12424),
            .in2(_gnd_net_),
            .in3(N__11609),
            .lcout(dout_obuf_RNO_4Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_4_LC_11_5_4.C_ON=1'b0;
    defparam dout_obuf_RNO_4_4_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_4_LC_11_5_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_4_4_LC_11_5_4 (
            .in0(N__11597),
            .in1(N__12423),
            .in2(_gnd_net_),
            .in3(N__11579),
            .lcout(dout_obuf_RNO_4Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_4_LC_11_10_0.C_ON=1'b0;
    defparam dout_obuf_RNO_1_4_LC_11_10_0.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_4_LC_11_10_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_1_4_LC_11_10_0 (
            .in0(N__11669),
            .in1(N__12728),
            .in2(_gnd_net_),
            .in3(N__11567),
            .lcout(),
            .ltout(mem_N_180_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_4_LC_11_10_1.C_ON=1'b0;
    defparam dout_obuf_RNO_4_LC_11_10_1.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_4_LC_11_10_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 dout_obuf_RNO_4_LC_11_10_1 (
            .in0(N__12578),
            .in1(_gnd_net_),
            .in2(N__11555),
            .in3(N__11756),
            .lcout(dout_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_6_LC_11_10_4.C_ON=1'b0;
    defparam dout_obuf_RNO_1_6_LC_11_10_4.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_6_LC_11_10_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_1_6_LC_11_10_4 (
            .in0(N__12729),
            .in1(N__12080),
            .in2(_gnd_net_),
            .in3(N__11534),
            .lcout(),
            .ltout(mem_N_145_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_6_LC_11_10_5.C_ON=1'b0;
    defparam dout_obuf_RNO_6_LC_11_10_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_6_LC_11_10_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 dout_obuf_RNO_6_LC_11_10_5 (
            .in0(N__12579),
            .in1(_gnd_net_),
            .in2(N__11525),
            .in3(N__11711),
            .lcout(dout_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_3_LC_11_11_2.C_ON=1'b0;
    defparam dout_obuf_RNO_1_3_LC_11_11_2.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_3_LC_11_11_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 dout_obuf_RNO_1_3_LC_11_11_2 (
            .in0(N__12748),
            .in1(N__11504),
            .in2(_gnd_net_),
            .in3(N__11492),
            .lcout(mem_N_174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_3_LC_11_11_4.C_ON=1'b0;
    defparam dout_obuf_RNO_2_3_LC_11_11_4.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_3_LC_11_11_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_2_3_LC_11_11_4 (
            .in0(N__11480),
            .in1(N__12327),
            .in2(_gnd_net_),
            .in3(N__11471),
            .lcout(),
            .ltout(dout_obuf_RNO_2Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_3_LC_11_11_5.C_ON=1'b0;
    defparam dout_obuf_RNO_0_3_LC_11_11_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_3_LC_11_11_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 dout_obuf_RNO_0_3_LC_11_11_5 (
            .in0(N__11456),
            .in1(_gnd_net_),
            .in2(N__11441),
            .in3(N__12747),
            .lcout(),
            .ltout(mem_N_172_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_LC_11_11_6.C_ON=1'b0;
    defparam dout_obuf_RNO_3_LC_11_11_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_LC_11_11_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 dout_obuf_RNO_3_LC_11_11_6 (
            .in0(N__11828),
            .in1(_gnd_net_),
            .in2(N__11822),
            .in3(N__12558),
            .lcout(dout_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_2_LC_11_13_4.C_ON=1'b0;
    defparam dout_obuf_RNO_1_2_LC_11_13_4.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_2_LC_11_13_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_1_2_LC_11_13_4 (
            .in0(N__12712),
            .in1(N__11627),
            .in2(_gnd_net_),
            .in3(N__11807),
            .lcout(mem_N_168),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_4_LC_11_13_6.C_ON=1'b0;
    defparam dout_obuf_RNO_2_4_LC_11_13_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_4_LC_11_13_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_2_4_LC_11_13_6 (
            .in0(N__11789),
            .in1(N__12402),
            .in2(_gnd_net_),
            .in3(N__11771),
            .lcout(),
            .ltout(dout_obuf_RNO_2Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_4_LC_11_13_7.C_ON=1'b0;
    defparam dout_obuf_RNO_0_4_LC_11_13_7.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_4_LC_11_13_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 dout_obuf_RNO_0_4_LC_11_13_7 (
            .in0(N__12711),
            .in1(_gnd_net_),
            .in2(N__11759),
            .in3(N__11966),
            .lcout(mem_N_178),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_6_LC_11_15_0.C_ON=1'b0;
    defparam dout_obuf_RNO_2_6_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_6_LC_11_15_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_2_6_LC_11_15_0 (
            .in0(N__11744),
            .in1(N__12320),
            .in2(_gnd_net_),
            .in3(N__11726),
            .lcout(),
            .ltout(dout_obuf_RNO_2Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_6_LC_11_15_1.C_ON=1'b0;
    defparam dout_obuf_RNO_0_6_LC_11_15_1.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_6_LC_11_15_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 dout_obuf_RNO_0_6_LC_11_15_1 (
            .in0(N__12713),
            .in1(_gnd_net_),
            .in2(N__11714),
            .in3(N__11879),
            .lcout(mem_N_144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_4_LC_11_19_1.C_ON=1'b0;
    defparam dout_obuf_RNO_5_4_LC_11_19_1.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_4_LC_11_19_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_5_4_LC_11_19_1 (
            .in0(N__12314),
            .in1(N__11699),
            .in2(_gnd_net_),
            .in3(N__11687),
            .lcout(dout_obuf_RNO_5Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_2_LC_11_19_2.C_ON=1'b0;
    defparam dout_obuf_RNO_5_2_LC_11_19_2.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_2_LC_11_19_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_5_2_LC_11_19_2 (
            .in0(N__11657),
            .in1(N__12313),
            .in2(_gnd_net_),
            .in3(N__11639),
            .lcout(dout_obuf_RNO_5Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_6_LC_11_23_3.C_ON=1'b0;
    defparam dout_obuf_RNO_5_6_LC_11_23_3.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_6_LC_11_23_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_5_6_LC_11_23_3 (
            .in0(N__12289),
            .in1(N__12110),
            .in2(_gnd_net_),
            .in3(N__12098),
            .lcout(dout_obuf_RNO_5Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_7_LC_11_23_7.C_ON=1'b0;
    defparam dout_obuf_RNO_5_7_LC_11_23_7.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_7_LC_11_23_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_5_7_LC_11_23_7 (
            .in0(N__12290),
            .in1(N__12068),
            .in2(_gnd_net_),
            .in3(N__12059),
            .lcout(dout_obuf_RNO_5Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_1_LC_11_25_4.C_ON=1'b0;
    defparam dout_obuf_RNO_3_1_LC_11_25_4.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_1_LC_11_25_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_3_1_LC_11_25_4 (
            .in0(N__12032),
            .in1(N__12357),
            .in2(_gnd_net_),
            .in3(N__12023),
            .lcout(dout_obuf_RNO_3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_4_LC_11_29_3.C_ON=1'b0;
    defparam dout_obuf_RNO_3_4_LC_11_29_3.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_4_LC_11_29_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_3_4_LC_11_29_3 (
            .in0(N__12335),
            .in1(N__11996),
            .in2(_gnd_net_),
            .in3(N__11984),
            .lcout(dout_obuf_RNO_3Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_7_LC_11_31_6.C_ON=1'b0;
    defparam dout_obuf_RNO_3_7_LC_11_31_6.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_7_LC_11_31_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_3_7_LC_11_31_6 (
            .in0(N__12264),
            .in1(N__11945),
            .in2(_gnd_net_),
            .in3(N__11936),
            .lcout(dout_obuf_RNO_3Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_6_LC_11_31_7.C_ON=1'b0;
    defparam dout_obuf_RNO_3_6_LC_11_31_7.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_6_LC_11_31_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_3_6_LC_11_31_7 (
            .in0(N__11909),
            .in1(N__12263),
            .in2(_gnd_net_),
            .in3(N__11897),
            .lcout(dout_obuf_RNO_3Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_1_5_LC_13_13_2.C_ON=1'b0;
    defparam dout_obuf_RNO_1_5_LC_13_13_2.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_1_5_LC_13_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 dout_obuf_RNO_1_5_LC_13_13_2 (
            .in0(N__12440),
            .in1(N__12684),
            .in2(_gnd_net_),
            .in3(N__11861),
            .lcout(mem_N_140),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_2_5_LC_13_13_3.C_ON=1'b0;
    defparam dout_obuf_RNO_2_5_LC_13_13_3.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_2_5_LC_13_13_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_2_5_LC_13_13_3 (
            .in0(N__11849),
            .in1(N__12399),
            .in2(_gnd_net_),
            .in3(N__11837),
            .lcout(),
            .ltout(dout_obuf_RNO_2Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_0_5_LC_13_13_4.C_ON=1'b0;
    defparam dout_obuf_RNO_0_5_LC_13_13_4.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_0_5_LC_13_13_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 dout_obuf_RNO_0_5_LC_13_13_4 (
            .in0(N__12683),
            .in1(_gnd_net_),
            .in2(N__12593),
            .in3(N__12122),
            .lcout(mem_N_139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_LC_13_13_5.C_ON=1'b0;
    defparam dout_obuf_RNO_5_LC_13_13_5.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_LC_13_13_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 dout_obuf_RNO_5_LC_13_13_5 (
            .in0(N__12590),
            .in1(N__12566),
            .in2(_gnd_net_),
            .in3(N__12488),
            .lcout(dout_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_5_5_LC_13_21_0.C_ON=1'b0;
    defparam dout_obuf_RNO_5_5_LC_13_21_0.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_5_5_LC_13_21_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_5_5_LC_13_21_0 (
            .in0(N__12365),
            .in1(N__12461),
            .in2(_gnd_net_),
            .in3(N__12452),
            .lcout(dout_obuf_RNO_5Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dout_obuf_RNO_3_5_LC_13_29_0.C_ON=1'b0;
    defparam dout_obuf_RNO_3_5_LC_13_29_0.SEQ_MODE=4'b0000;
    defparam dout_obuf_RNO_3_5_LC_13_29_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 dout_obuf_RNO_3_5_LC_13_29_0 (
            .in0(N__12329),
            .in1(N__12143),
            .in2(_gnd_net_),
            .in3(N__12134),
            .lcout(dout_obuf_RNO_3Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // RAM
