// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Sep 14 01:22:08 2018
//
// Verilog Description of module main
//

module main (DEBUG, TVP_CLK, TVP_HSYNC, TVP_VSYNC, TVP_VIDEO, LED, 
            ADV_HSYNC, ADV_VSYNC, ADV_R, ADV_G, ADV_B, ADV_CLK, 
            ADV_SYNC_N, ADV_BLANK_N) /* synthesis syn_module_defined=1 */ ;   // ../main.v(1[8:12])
    output [7:0]DEBUG;   // ../main.v(2[19:24])
    input TVP_CLK;   // ../main.v(3[13:20])
    input TVP_HSYNC;   // ../main.v(4[13:22])
    input TVP_VSYNC;   // ../main.v(5[13:22])
    input [9:0]TVP_VIDEO;   // ../main.v(6[19:28])
    output LED;   // ../main.v(7[14:17])
    output ADV_HSYNC;   // ../main.v(8[14:23])
    output ADV_VSYNC;   // ../main.v(9[14:23])
    output [7:0]ADV_R;   // ../main.v(10[19:24])
    output [7:0]ADV_G;   // ../main.v(11[19:24])
    output [7:0]ADV_B;   // ../main.v(12[19:24])
    output ADV_CLK;   // ../main.v(13[14:21])
    output ADV_SYNC_N;   // ../main.v(14[14:24])
    output ADV_BLANK_N;   // ../main.v(15[14:25])
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    
    wire GND_net, VCC_net, DEBUG_c_7, DEBUG_c_6, DEBUG_c_5, DEBUG_c_4, 
        DEBUG_c_3, DEBUG_c_2, DEBUG_c_1, DEBUG_c_0, TVP_HSYNC_c, TVP_VSYNC_c, 
        TVP_VIDEO_c_9, TVP_VIDEO_c_8, TVP_VIDEO_c_7, TVP_VIDEO_c_6, 
        TVP_VIDEO_c_5, TVP_VIDEO_c_4, TVP_VIDEO_c_3, TVP_VIDEO_c_2, 
        LED_c, ADV_HSYNC_c, ADV_VSYNC_c, ADV_B_c, n1949, n1950, 
        n1951, n1952, n1953, n1954, n1955;
    wire [13:0]RX_ADDR;   // ../main.v(28[14:21])
    wire [13:0]TX_ADDR;   // ../main.v(45[14:21])
    wire [7:0]TX_DATA;   // ../main.v(46[13:20])
    
    wire VGA_VISIBLE, n3184, n25, n28;
    wire [8:0]Y;   // ../o_counter.v(48[19:20])
    
    wire n2147, n3009, n27, n26, n25_adj_573, n24, n23, n22, 
        n21, n20, n19, n18, n5;
    
    VCC i2 (.Y(VCC_net));
    RX receive_module (.n25(n25), .TVP_VSYNC_c(TVP_VSYNC_c), .RX_ADDR({RX_ADDR}), 
       .TVP_CLK_c(TVP_CLK_c), .GND_net(GND_net), .VCC_net(VCC_net), .TVP_HSYNC_c(TVP_HSYNC_c), 
       .\Y[1] (Y[1]), .n3184(n3184), .LED_c(LED_c), .\Y[0] (Y[0]), .n3009(n3009), 
       .n2147(n2147), .n5(n5)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(32[5] 42[25])
    TX transmit_module (.DEBUG_c_3(DEBUG_c_3), .GND_net(GND_net), .DEBUG_c_2(DEBUG_c_2), 
       .DEBUG_c_0(DEBUG_c_0), .n28(n28), .ADV_CLK_c(ADV_CLK_c), .ADV_VSYNC_c(ADV_VSYNC_c), 
       .DEBUG_c_5(DEBUG_c_5), .VGA_VISIBLE(VGA_VISIBLE), .n23(n23), .DEBUG_c_6(DEBUG_c_6), 
       .DEBUG_c_4(DEBUG_c_4), .n24(n24), .n18(n18), .n25(n25_adj_573), 
       .n19(n19), .n26(n26), .n20(n20), .DEBUG_c_1(DEBUG_c_1), .n27(n27), 
       .\TX_ADDR[11] (TX_ADDR[11]), .DEBUG_c_7(DEBUG_c_7), .n21(n21), 
       .n22(n22), .\TX_ADDR[12] (TX_ADDR[12]), .\TX_ADDR[13] (TX_ADDR[13]), 
       .VCC_net(VCC_net), .n2147(n2147), .ADV_HSYNC_c(ADV_HSYNC_c), .n5(n5), 
       .n3009(n3009), .\Y[1] (Y[1]), .\Y[0] (Y[0])) /* synthesis syn_module_defined=1 */ ;   // ../main.v(48[5] 59[27])
    SB_GB_IO TVP_CLK_pad (.PACKAGE_PIN(TVP_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(TVP_CLK_c));   // ../main.v(3[13:20])
    defparam TVP_CLK_pad.PIN_TYPE = 6'b000001;
    defparam TVP_CLK_pad.PULLUP = 1'b0;
    defparam TVP_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_VSYNC_pad (.PACKAGE_PIN(ADV_VSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_VSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_VSYNC_pad.PIN_TYPE = 6'b011001;
    defparam ADV_VSYNC_pad.PULLUP = 1'b0;
    defparam ADV_VSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_VSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_7 (.PACKAGE_PIN(ADV_R[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_7.PULLUP = 1'b0;
    defparam ADV_R_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_4 (.PACKAGE_PIN(DEBUG[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_4));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_4.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_4.PULLUP = 1'b0;
    defparam DEBUG_pad_4.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_8 (.PACKAGE_PIN(TVP_VIDEO[8]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_8));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_8.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_8.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_8.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_8.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_HSYNC_pad (.PACKAGE_PIN(TVP_HSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_HSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_HSYNC_pad.PIN_TYPE = 6'b000001;
    defparam TVP_HSYNC_pad.PULLUP = 1'b0;
    defparam TVP_HSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_HSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_7 (.PACKAGE_PIN(TVP_VIDEO[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_7));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_7.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_7.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_7.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_0 (.PACKAGE_PIN(DEBUG[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_0));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_0.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_0.PULLUP = 1'b0;
    defparam DEBUG_pad_0.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_1 (.PACKAGE_PIN(DEBUG[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_1));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_1.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_1.PULLUP = 1'b0;
    defparam DEBUG_pad_1.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_BLANK_N_pad (.PACKAGE_PIN(ADV_BLANK_N), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_BLANK_N_pad.PIN_TYPE = 6'b011001;
    defparam ADV_BLANK_N_pad.PULLUP = 1'b0;
    defparam ADV_BLANK_N_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_BLANK_N_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_2 (.PACKAGE_PIN(DEBUG[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_2));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_2.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_2.PULLUP = 1'b0;
    defparam DEBUG_pad_2.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_9 (.PACKAGE_PIN(TVP_VIDEO[9]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_9));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_9.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_9.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_9.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_9.IO_STANDARD = "SB_LVCMOS";
    SB_DFFNSR ADV_R__i8 (.Q(ADV_B_c), .C(ADV_CLK_c), .D(TX_DATA[7]), .R(VGA_VISIBLE));   // ../main.v(61[9] 65[5])
    SB_IO TVP_VIDEO_pad_6 (.PACKAGE_PIN(TVP_VIDEO[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_6));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_6.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_6.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_6.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_3 (.PACKAGE_PIN(DEBUG[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_3));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_3.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_3.PULLUP = 1'b0;
    defparam DEBUG_pad_3.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_5 (.PACKAGE_PIN(DEBUG[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_5));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_5.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_5.PULLUP = 1'b0;
    defparam DEBUG_pad_5.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_DFFNSR ADV_R__i7 (.Q(n1949), .C(ADV_CLK_c), .D(TX_DATA[6]), .R(VGA_VISIBLE));   // ../main.v(61[9] 65[5])
    SB_IO DEBUG_pad_6 (.PACKAGE_PIN(DEBUG[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_6));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_6.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_6.PULLUP = 1'b0;
    defparam DEBUG_pad_6.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_DFFNSR ADV_R__i6 (.Q(n1950), .C(ADV_CLK_c), .D(TX_DATA[5]), .R(VGA_VISIBLE));   // ../main.v(61[9] 65[5])
    SB_DFFNSR ADV_R__i5 (.Q(n1951), .C(ADV_CLK_c), .D(TX_DATA[4]), .R(VGA_VISIBLE));   // ../main.v(61[9] 65[5])
    SB_DFFNSR ADV_R__i4 (.Q(n1952), .C(ADV_CLK_c), .D(TX_DATA[3]), .R(VGA_VISIBLE));   // ../main.v(61[9] 65[5])
    SB_DFFNSR ADV_R__i3 (.Q(n1953), .C(ADV_CLK_c), .D(TX_DATA[2]), .R(VGA_VISIBLE));   // ../main.v(61[9] 65[5])
    SB_DFFNSR ADV_R__i2 (.Q(n1954), .C(ADV_CLK_c), .D(TX_DATA[1]), .R(VGA_VISIBLE));   // ../main.v(61[9] 65[5])
    SB_IO DEBUG_pad_7 (.PACKAGE_PIN(DEBUG[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_7));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_7.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_7.PULLUP = 1'b0;
    defparam DEBUG_pad_7.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_5 (.PACKAGE_PIN(TVP_VIDEO[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_5));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_5.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_5.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_5.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_DFFNSR ADV_R__i1 (.Q(n1955), .C(ADV_CLK_c), .D(TX_DATA[0]), .R(VGA_VISIBLE));   // ../main.v(61[9] 65[5])
    SB_IO TVP_VSYNC_pad (.PACKAGE_PIN(TVP_VSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VSYNC_pad.PIN_TYPE = 6'b000001;
    defparam TVP_VSYNC_pad.PULLUP = 1'b0;
    defparam TVP_VSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_VSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_SYNC_N_pad (.PACKAGE_PIN(ADV_SYNC_N), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_SYNC_N_pad.PIN_TYPE = 6'b011001;
    defparam ADV_SYNC_N_pad.PULLUP = 1'b0;
    defparam ADV_SYNC_N_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_SYNC_N_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_CLK_pad (.PACKAGE_PIN(ADV_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(ADV_CLK_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_CLK_pad.PIN_TYPE = 6'b011001;
    defparam ADV_CLK_pad.PULLUP = 1'b0;
    defparam ADV_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_0 (.PACKAGE_PIN(ADV_B[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1955));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_0.PULLUP = 1'b0;
    defparam ADV_B_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_1 (.PACKAGE_PIN(ADV_B[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1954));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_1.PULLUP = 1'b0;
    defparam ADV_B_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_2 (.PACKAGE_PIN(ADV_B[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1953));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_2.PULLUP = 1'b0;
    defparam ADV_B_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_3 (.PACKAGE_PIN(ADV_B[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1952));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_3.PULLUP = 1'b0;
    defparam ADV_B_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_4 (.PACKAGE_PIN(ADV_B[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1951));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_4.PULLUP = 1'b0;
    defparam ADV_B_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_5 (.PACKAGE_PIN(ADV_B[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1950));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_5.PULLUP = 1'b0;
    defparam ADV_B_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_6 (.PACKAGE_PIN(ADV_B[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1949));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_6.PULLUP = 1'b0;
    defparam ADV_B_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_7 (.PACKAGE_PIN(ADV_B[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_7.PULLUP = 1'b0;
    defparam ADV_B_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_0 (.PACKAGE_PIN(ADV_G[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1955));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_0.PULLUP = 1'b0;
    defparam ADV_G_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_1 (.PACKAGE_PIN(ADV_G[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1954));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_1.PULLUP = 1'b0;
    defparam ADV_G_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_2 (.PACKAGE_PIN(ADV_G[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1953));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_2.PULLUP = 1'b0;
    defparam ADV_G_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_3 (.PACKAGE_PIN(ADV_G[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1952));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_3.PULLUP = 1'b0;
    defparam ADV_G_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_4 (.PACKAGE_PIN(ADV_G[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1951));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_4.PULLUP = 1'b0;
    defparam ADV_G_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_5 (.PACKAGE_PIN(ADV_G[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1950));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_5.PULLUP = 1'b0;
    defparam ADV_G_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_6 (.PACKAGE_PIN(ADV_G[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1949));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_6.PULLUP = 1'b0;
    defparam ADV_G_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_7 (.PACKAGE_PIN(ADV_G[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_7.PULLUP = 1'b0;
    defparam ADV_G_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_0 (.PACKAGE_PIN(ADV_R[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1955));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_0.PULLUP = 1'b0;
    defparam ADV_R_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_1 (.PACKAGE_PIN(ADV_R[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1954));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_1.PULLUP = 1'b0;
    defparam ADV_R_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_2 (.PACKAGE_PIN(ADV_R[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1953));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_2.PULLUP = 1'b0;
    defparam ADV_R_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_3 (.PACKAGE_PIN(ADV_R[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1952));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_3.PULLUP = 1'b0;
    defparam ADV_R_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_4 (.PACKAGE_PIN(ADV_R[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1951));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_4.PULLUP = 1'b0;
    defparam ADV_R_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_5 (.PACKAGE_PIN(ADV_R[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1950));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_5.PULLUP = 1'b0;
    defparam ADV_R_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_6 (.PACKAGE_PIN(ADV_R[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1949));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_6.PULLUP = 1'b0;
    defparam ADV_R_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_4 (.PACKAGE_PIN(TVP_VIDEO[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_4));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_4.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_4.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_4.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_3 (.PACKAGE_PIN(TVP_VIDEO[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_3));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_3.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_3.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_3.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_2 (.PACKAGE_PIN(TVP_VIDEO[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_2));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_2.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_2.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_2.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_HSYNC_pad (.PACKAGE_PIN(ADV_HSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_HSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_HSYNC_pad.PIN_TYPE = 6'b011001;
    defparam ADV_HSYNC_pad.PULLUP = 1'b0;
    defparam ADV_HSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_HSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    GND i1 (.Y(GND_net));
    SB_LUT4 i27_1_lut_rep_20 (.I0(TVP_HSYNC_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3184));   // ../main.v(4[13:22])
    defparam i27_1_lut_rep_20.LUT_INIT = 16'h5555;
    TX_PLL tx_pll (.TVP_CLK_c(TVP_CLK_c), .VCC_net(VCC_net), .GND_net(GND_net), 
           .ADV_CLK_c(ADV_CLK_c)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(20[9] 24[25])
    RAM line_buffer (.TX_DATA({TX_DATA}), .ADV_CLK_c(ADV_CLK_c), .\TX_ADDR[12] (TX_ADDR[12]), 
        .n25(n25), .RX_ADDR({RX_ADDR}), .\TX_ADDR[13] (TX_ADDR[13]), .GND_net(GND_net), 
        .\TX_ADDR[11] (TX_ADDR[11]), .n28(n28), .n27(n27), .n26(n26), 
        .n25_adj_1(n25_adj_573), .n24(n24), .n23(n23), .n22(n22), .n21(n21), 
        .n20(n20), .n19(n19), .n18(n18), .TVP_VIDEO_c_8(TVP_VIDEO_c_8), 
        .TVP_VIDEO_c_9(TVP_VIDEO_c_9), .TVP_CLK_c(TVP_CLK_c), .VCC_net(VCC_net), 
        .TVP_VIDEO_c_6(TVP_VIDEO_c_6), .TVP_VIDEO_c_7(TVP_VIDEO_c_7), .TVP_VIDEO_c_4(TVP_VIDEO_c_4), 
        .TVP_VIDEO_c_5(TVP_VIDEO_c_5), .TVP_VIDEO_c_2(TVP_VIDEO_c_2), .TVP_VIDEO_c_3(TVP_VIDEO_c_3)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(68[6] 74[21])
    
endmodule
//
// Verilog Description of module RX
//

module RX (n25, TVP_VSYNC_c, RX_ADDR, TVP_CLK_c, GND_net, VCC_net, 
           TVP_HSYNC_c, \Y[1] , n3184, LED_c, \Y[0] , n3009, n2147, 
           n5) /* synthesis syn_module_defined=1 */ ;
    output n25;
    input TVP_VSYNC_c;
    output [13:0]RX_ADDR;
    input TVP_CLK_c;
    input GND_net;
    input VCC_net;
    input TVP_HSYNC_c;
    output \Y[1] ;
    input n3184;
    output LED_c;
    output \Y[0] ;
    output n3009;
    input n2147;
    output n5;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire [13:0]n122;
    
    wire n2323, n3181, n3185, n2730, n2735, n2736, n2739, n2728, 
        n2729, n2325, n2734, n2327, n2329, n2733, n2738, n2331, 
        n2731, n2727, n2737, n2732, n2333, n2335, n2337, n2339, 
        n2341, old_HS, n2152, old_VS, n252, n2321;
    
    SB_LUT4 i966_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[9]), 
            .I3(RX_ADDR[9]), .O(n2323));
    defparam i966_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFESR BRAM_ADDR__i12 (.Q(RX_ADDR[12]), .C(TVP_CLK_c), .E(n3181), 
            .D(n122[12]), .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(RX_ADDR[4]), .I2(GND_net), 
            .I3(n2730), .O(n122[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n2735), .I0(RX_ADDR[9]), .I1(GND_net), .CO(n2736));
    SB_DFFESR BRAM_ADDR__i11 (.Q(RX_ADDR[11]), .C(TVP_CLK_c), .E(n3181), 
            .D(n122[11]), .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(RX_ADDR[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n122[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(RX_ADDR[13]), .I2(GND_net), 
            .I3(n2739), .O(n122[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_4 (.CI(n2728), .I0(RX_ADDR[2]), .I1(GND_net), .CO(n2729));
    SB_LUT4 i968_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[8]), 
            .I3(RX_ADDR[8]), .O(n2325));
    defparam i968_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(RX_ADDR[8]), .I2(GND_net), 
            .I3(n2734), .O(n122[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i970_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[7]), 
            .I3(RX_ADDR[7]), .O(n2327));
    defparam i970_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i972_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[6]), 
            .I3(RX_ADDR[6]), .O(n2329));
    defparam i972_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_CARRY add_12_10 (.CI(n2734), .I0(RX_ADDR[8]), .I1(GND_net), .CO(n2735));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(RX_ADDR[7]), .I2(GND_net), 
            .I3(n2733), .O(n122[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(RX_ADDR[12]), .I2(GND_net), 
            .I3(n2738), .O(n122[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n2738), .I0(RX_ADDR[12]), .I1(GND_net), .CO(n2739));
    SB_LUT4 i974_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[5]), 
            .I3(RX_ADDR[5]), .O(n2331));
    defparam i974_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_CARRY add_12_6 (.CI(n2730), .I0(RX_ADDR[4]), .I1(GND_net), .CO(n2731));
    SB_CARRY add_12_2 (.CI(VCC_net), .I0(RX_ADDR[0]), .I1(GND_net), .CO(n2727));
    SB_CARRY add_12_9 (.CI(n2733), .I0(RX_ADDR[7]), .I1(GND_net), .CO(n2734));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(RX_ADDR[1]), .I2(GND_net), 
            .I3(n2727), .O(n122[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(RX_ADDR[11]), .I2(GND_net), 
            .I3(n2737), .O(n122[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(RX_ADDR[3]), .I2(GND_net), 
            .I3(n2729), .O(n122[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(RX_ADDR[6]), .I2(GND_net), 
            .I3(n2732), .O(n122[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_13 (.CI(n2737), .I0(RX_ADDR[11]), .I1(GND_net), .CO(n2738));
    SB_CARRY add_12_8 (.CI(n2732), .I0(RX_ADDR[6]), .I1(GND_net), .CO(n2733));
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(RX_ADDR[5]), .I2(GND_net), 
            .I3(n2731), .O(n122[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i976_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[0]), 
            .I3(RX_ADDR[0]), .O(n2333));
    defparam i976_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_CARRY add_12_3 (.CI(n2727), .I0(RX_ADDR[1]), .I1(GND_net), .CO(n2728));
    SB_CARRY add_12_7 (.CI(n2731), .I0(RX_ADDR[5]), .I1(GND_net), .CO(n2732));
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(RX_ADDR[10]), .I2(GND_net), 
            .I3(n2736), .O(n122[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n2736), .I0(RX_ADDR[10]), .I1(GND_net), .CO(n2737));
    SB_CARRY add_12_5 (.CI(n2729), .I0(RX_ADDR[3]), .I1(GND_net), .CO(n2730));
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(RX_ADDR[2]), .I2(GND_net), 
            .I3(n2728), .O(n122[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(RX_ADDR[9]), .I2(GND_net), 
            .I3(n2735), .O(n122[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i978_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[4]), 
            .I3(RX_ADDR[4]), .O(n2335));
    defparam i978_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i980_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[3]), 
            .I3(RX_ADDR[3]), .O(n2337));
    defparam i980_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i982_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[2]), 
            .I3(RX_ADDR[2]), .O(n2339));
    defparam i982_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i984_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[1]), 
            .I3(RX_ADDR[1]), .O(n2341));
    defparam i984_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i297_3_lut_3_lut_3_lut (.I0(TVP_VSYNC_c), .I1(old_HS), .I2(TVP_HSYNC_c), 
            .I3(GND_net), .O(n2152));   // ../main.v(5[13:22])
    defparam i297_3_lut_3_lut_3_lut.LUT_INIT = 16'h5d5d;
    SB_LUT4 i141_2_lut_2_lut (.I0(TVP_VSYNC_c), .I1(old_VS), .I2(GND_net), 
            .I3(GND_net), .O(n252));   // ../main.v(5[13:22])
    defparam i141_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i24_1_lut_rep_21 (.I0(TVP_VSYNC_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3185));   // ../main.v(5[13:22])
    defparam i24_1_lut_rep_21.LUT_INIT = 16'h5555;
    SB_LUT4 i1632_2_lut_rep_17 (.I0(n25), .I1(TVP_VSYNC_c), .I2(GND_net), 
            .I3(GND_net), .O(n3181));
    defparam i1632_2_lut_rep_17.LUT_INIT = 16'h7777;
    SB_DFFESR BRAM_ADDR__i13 (.Q(RX_ADDR[13]), .C(TVP_CLK_c), .E(n3181), 
            .D(n122[13]), .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i1 (.Q(RX_ADDR[1]), .C(TVP_CLK_c), .D(n2341), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i2 (.Q(RX_ADDR[2]), .C(TVP_CLK_c), .D(n2339), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i3 (.Q(RX_ADDR[3]), .C(TVP_CLK_c), .D(n2337), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i4 (.Q(RX_ADDR[4]), .C(TVP_CLK_c), .D(n2335), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i0 (.Q(RX_ADDR[0]), .C(TVP_CLK_c), .D(n2333), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i5 (.Q(RX_ADDR[5]), .C(TVP_CLK_c), .D(n2331), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i6 (.Q(RX_ADDR[6]), .C(TVP_CLK_c), .D(n2329), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i7 (.Q(RX_ADDR[7]), .C(TVP_CLK_c), .D(n2327), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i8 (.Q(RX_ADDR[8]), .C(TVP_CLK_c), .D(n2325), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i9 (.Q(RX_ADDR[9]), .C(TVP_CLK_c), .D(n2323), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_DFFSR BRAM_ADDR__i10 (.Q(RX_ADDR[10]), .C(TVP_CLK_c), .D(n2321), 
            .R(n3185));   // ../rx.v(50[12] 59[8])
    SB_LUT4 i964_3_lut_4_lut (.I0(n25), .I1(TVP_VSYNC_c), .I2(n122[10]), 
            .I3(RX_ADDR[10]), .O(n2321));
    defparam i964_3_lut_4_lut.LUT_INIT = 16'hf870;
    O_COUNTER rx_counter (.VCC_net(VCC_net), .GND_net(GND_net), .TVP_HSYNC_c(TVP_HSYNC_c), 
            .old_HS(old_HS), .TVP_CLK_c(TVP_CLK_c), .TVP_VSYNC_c(TVP_VSYNC_c), 
            .old_VS(old_VS), .\Y[1] (\Y[1] ), .n3184(n3184), .n252(n252), 
            .LED_c(LED_c), .\Y[0] (\Y[0] ), .n2152(n2152), .n3185(n3185), 
            .n25(n25), .n3009(n3009), .n2147(n2147), .n5(n5)) /* synthesis syn_module_defined=1 */ ;   // ../rx.v(40[15] 48[41])
    
endmodule
//
// Verilog Description of module O_COUNTER
//

module O_COUNTER (VCC_net, GND_net, TVP_HSYNC_c, old_HS, TVP_CLK_c, 
            TVP_VSYNC_c, old_VS, \Y[1] , n3184, n252, LED_c, \Y[0] , 
            n2152, n3185, n25, n3009, n2147, n5) /* synthesis syn_module_defined=1 */ ;
    input VCC_net;
    input GND_net;
    input TVP_HSYNC_c;
    output old_HS;
    input TVP_CLK_c;
    input TVP_VSYNC_c;
    output old_VS;
    output \Y[1] ;
    input n3184;
    input n252;
    output LED_c;
    output \Y[0] ;
    input n2152;
    input n3185;
    output n25;
    output n3009;
    input n2147;
    output n5;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire [9:0]n79;
    
    wire n2782;
    wire [9:0]n45;
    
    wire n2783, n2784;
    wire [9:0]X;   // ../o_counter.v(47[19:20])
    
    wire n2785, n2786, n2787, n2788;
    wire [8:0]n301;
    wire [8:0]Y;   // ../o_counter.v(48[19:20])
    
    wire n2765, n2764, n2763, n2762, n4, n2761, n2760, n2759, 
        n2758, n3166, PULSE_1HZ_N_92;
    wire [5:0]FRAME_COUNTER;   // ../o_counter.v(46[19:32])
    
    wire n10_adj_570;
    wire [5:0]n29;
    
    wire n2757, n2978, n2756, n2755, n2754, n2900, n2943, n2753, 
        n2975, n2986, n7, n4_adj_571, n31_adj_572, n2989, n6, 
        n2227, n2790, n2789;
    
    SB_CARRY X_284_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n79[0]), .CO(n2782));
    SB_LUT4 X_284_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n79[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_284_add_4_3 (.CI(n2782), .I0(GND_net), .I1(n79[1]), .CO(n2783));
    SB_LUT4 X_284_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(n79[1]), 
            .I3(n2782), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_284_add_4_4 (.CI(n2783), .I0(GND_net), .I1(n79[2]), .CO(n2784));
    SB_DFF old_HS_48 (.Q(old_HS), .C(TVP_CLK_c), .D(TVP_HSYNC_c));   // ../o_counter.v(51[16] 79[12])
    SB_LUT4 X_284_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(n79[2]), 
            .I3(n2783), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_284_add_4_5 (.CI(n2784), .I0(GND_net), .I1(X[3]), .CO(n2785));
    SB_DFF old_VS_49 (.Q(old_VS), .C(TVP_CLK_c), .D(TVP_VSYNC_c));   // ../o_counter.v(51[16] 79[12])
    SB_LUT4 X_284_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(X[3]), 
            .I3(n2784), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_284_add_4_6 (.CI(n2785), .I0(GND_net), .I1(X[4]), .CO(n2786));
    SB_LUT4 X_284_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(X[4]), 
            .I3(n2785), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_284_add_4_7 (.CI(n2786), .I0(GND_net), .I1(X[5]), .CO(n2787));
    SB_LUT4 X_284_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(X[5]), 
            .I3(n2786), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 X_284_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(X[6]), 
            .I3(n2787), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_284_add_4_8 (.CI(n2787), .I0(GND_net), .I1(X[6]), .CO(n2788));
    SB_LUT4 add_63_10_lut (.I0(GND_net), .I1(Y[8]), .I2(GND_net), .I3(n2765), 
            .O(n301[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_63_9_lut (.I0(GND_net), .I1(Y[7]), .I2(GND_net), .I3(n2764), 
            .O(n301[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_63_9 (.CI(n2764), .I0(Y[7]), .I1(GND_net), .CO(n2765));
    SB_LUT4 add_63_8_lut (.I0(GND_net), .I1(Y[6]), .I2(GND_net), .I3(n2763), 
            .O(n301[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_63_8 (.CI(n2763), .I0(Y[6]), .I1(GND_net), .CO(n2764));
    SB_LUT4 add_63_7_lut (.I0(GND_net), .I1(Y[5]), .I2(GND_net), .I3(n2762), 
            .O(n301[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_63_7 (.CI(n2762), .I0(Y[5]), .I1(GND_net), .CO(n2763));
    SB_LUT4 i1_2_lut (.I0(Y[4]), .I1(Y[3]), .I2(GND_net), .I3(GND_net), 
            .O(n4));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_63_6_lut (.I0(GND_net), .I1(Y[4]), .I2(GND_net), .I3(n2761), 
            .O(n301[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_63_6 (.CI(n2761), .I0(Y[4]), .I1(GND_net), .CO(n2762));
    SB_LUT4 add_63_5_lut (.I0(GND_net), .I1(Y[3]), .I2(GND_net), .I3(n2760), 
            .O(n301[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_63_5 (.CI(n2760), .I0(Y[3]), .I1(GND_net), .CO(n2761));
    SB_LUT4 add_63_4_lut (.I0(GND_net), .I1(Y[2]), .I2(GND_net), .I3(n2759), 
            .O(n301[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_63_4 (.CI(n2759), .I0(Y[2]), .I1(GND_net), .CO(n2760));
    SB_LUT4 add_63_3_lut (.I0(GND_net), .I1(\Y[1] ), .I2(GND_net), .I3(n2758), 
            .O(n301[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_rep_2_2_lut (.I0(Y[6]), .I1(Y[5]), .I2(GND_net), .I3(GND_net), 
            .O(n3166));
    defparam i1_rep_2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFSR X_284__i0 (.Q(n79[0]), .C(TVP_CLK_c), .D(n45[0]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_DFFE PULSE_1HZ_46 (.Q(LED_c), .C(TVP_CLK_c), .E(n252), .D(PULSE_1HZ_N_92));   // ../o_counter.v(51[16] 79[12])
    SB_LUT4 i4_4_lut (.I0(FRAME_COUNTER[2]), .I1(FRAME_COUNTER[3]), .I2(FRAME_COUNTER[4]), 
            .I3(FRAME_COUNTER[1]), .O(n10_adj_570));
    defparam i4_4_lut.LUT_INIT = 16'hbfff;
    SB_CARRY add_63_3 (.CI(n2758), .I0(\Y[1] ), .I1(GND_net), .CO(n2759));
    SB_LUT4 add_63_2_lut (.I0(GND_net), .I1(\Y[0] ), .I2(GND_net), .I3(VCC_net), 
            .O(n301[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_63_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_63_2 (.CI(VCC_net), .I0(\Y[0] ), .I1(GND_net), .CO(n2758));
    SB_LUT4 FRAME_COUNTER_285_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[5]), 
            .I3(n2757), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_285_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut (.I0(Y[2]), .I1(Y[3]), .I2(\Y[0] ), .I3(\Y[1] ), 
            .O(n2978));
    defparam i2_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 FRAME_COUNTER_285_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[4]), 
            .I3(n2756), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_285_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_285_add_4_6 (.CI(n2756), .I0(GND_net), .I1(FRAME_COUNTER[4]), 
            .CO(n2757));
    SB_LUT4 FRAME_COUNTER_285_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[3]), 
            .I3(n2755), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_285_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_285_add_4_5 (.CI(n2755), .I0(GND_net), .I1(FRAME_COUNTER[3]), 
            .CO(n2756));
    SB_LUT4 FRAME_COUNTER_285_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[2]), 
            .I3(n2754), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_285_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1499_3_lut (.I0(X[6]), .I1(X[7]), .I2(n2900), .I3(GND_net), 
            .O(n2943));
    defparam i1499_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY FRAME_COUNTER_285_add_4_4 (.CI(n2754), .I0(GND_net), .I1(FRAME_COUNTER[2]), 
            .CO(n2755));
    SB_LUT4 FRAME_COUNTER_285_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[1]), 
            .I3(n2753), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_285_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_285_add_4_3 (.CI(n2753), .I0(GND_net), .I1(FRAME_COUNTER[1]), 
            .CO(n2754));
    SB_LUT4 FRAME_COUNTER_285_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[0]), 
            .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_285_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_285_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(FRAME_COUNTER[0]), 
            .CO(n2753));
    SB_LUT4 i2_3_lut (.I0(X[6]), .I1(X[7]), .I2(n2900), .I3(GND_net), 
            .O(n2975));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_17 (.I0(Y[2]), .I1(n4), .I2(\Y[1] ), .I3(\Y[0] ), 
            .O(n2986));
    defparam i2_4_lut_adj_17.LUT_INIT = 16'hccc8;
    SB_LUT4 i2_2_lut (.I0(Y[6]), .I1(Y[7]), .I2(GND_net), .I3(GND_net), 
            .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(Y[8]), .I1(n2978), .I2(n3166), .I3(Y[4]), 
            .O(n4_adj_571));   // ../o_counter.v(81[28:148])
    defparam i1_4_lut.LUT_INIT = 16'ha8a0;
    SB_DFFESR Y__i0 (.Q(\Y[0] ), .C(TVP_CLK_c), .E(n2152), .D(n301[0]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_LUT4 i38_4_lut (.I0(X[8]), .I1(n2975), .I2(X[9]), .I3(n2943), 
            .O(n31_adj_572));   // ../o_counter.v(81[28:148])
    defparam i38_4_lut.LUT_INIT = 16'he0e5;
    SB_LUT4 i4_4_lut_adj_18 (.I0(n7), .I1(Y[8]), .I2(Y[5]), .I3(n2986), 
            .O(n2989));
    defparam i4_4_lut_adj_18.LUT_INIT = 16'hfffe;
    SB_DFFSR X_284__i1 (.Q(n79[1]), .C(TVP_CLK_c), .D(n45[1]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_LUT4 i2_3_lut_adj_19 (.I0(X[4]), .I1(X[5]), .I2(X[3]), .I3(GND_net), 
            .O(n2900));   // ../o_counter.v(81[61:90])
    defparam i2_3_lut_adj_19.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_20 (.I0(n2989), .I1(n31_adj_572), .I2(Y[7]), 
            .I3(n4_adj_571), .O(n25));   // ../o_counter.v(81[28:148])
    defparam i2_4_lut_adj_20.LUT_INIT = 16'hfddd;
    SB_LUT4 i1_2_lut_adj_21 (.I0(Y[4]), .I1(Y[7]), .I2(GND_net), .I3(GND_net), 
            .O(n6));
    defparam i1_2_lut_adj_21.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_22 (.I0(Y[8]), .I1(Y[3]), .I2(Y[2]), .I3(n6), 
            .O(n3009));
    defparam i4_4_lut_adj_22.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut (.I0(n2147), .I1(Y[6]), .I2(Y[5]), .I3(GND_net), 
            .O(n5));
    defparam i1_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFFESR Y__i8 (.Q(Y[8]), .C(TVP_CLK_c), .E(n2152), .D(n301[8]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_DFFESR Y__i7 (.Q(Y[7]), .C(TVP_CLK_c), .E(n2152), .D(n301[7]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_DFFESR Y__i6 (.Q(Y[6]), .C(TVP_CLK_c), .E(n2152), .D(n301[6]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_DFFESR Y__i5 (.Q(Y[5]), .C(TVP_CLK_c), .E(n2152), .D(n301[5]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_DFFESR Y__i4 (.Q(Y[4]), .C(TVP_CLK_c), .E(n2152), .D(n301[4]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_DFFESR Y__i3 (.Q(Y[3]), .C(TVP_CLK_c), .E(n2152), .D(n301[3]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_DFFESR Y__i2 (.Q(Y[2]), .C(TVP_CLK_c), .E(n2152), .D(n301[2]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_DFFESR Y__i1 (.Q(\Y[1] ), .C(TVP_CLK_c), .E(n2152), .D(n301[1]), 
            .R(n3185));   // ../o_counter.v(51[16] 79[12])
    SB_DFFESR FRAME_COUNTER_285__i2 (.Q(FRAME_COUNTER[2]), .C(TVP_CLK_c), 
            .E(n252), .D(n29[2]), .R(n2227));   // ../o_counter.v(71[46:63])
    SB_DFFESR FRAME_COUNTER_285__i3 (.Q(FRAME_COUNTER[3]), .C(TVP_CLK_c), 
            .E(n252), .D(n29[3]), .R(n2227));   // ../o_counter.v(71[46:63])
    SB_DFFESR FRAME_COUNTER_285__i0 (.Q(FRAME_COUNTER[0]), .C(TVP_CLK_c), 
            .E(n252), .D(n29[0]), .R(n2227));   // ../o_counter.v(71[46:63])
    SB_DFFESR FRAME_COUNTER_285__i4 (.Q(FRAME_COUNTER[4]), .C(TVP_CLK_c), 
            .E(n252), .D(n29[4]), .R(n2227));   // ../o_counter.v(71[46:63])
    SB_DFFESR FRAME_COUNTER_285__i5 (.Q(FRAME_COUNTER[5]), .C(TVP_CLK_c), 
            .E(n252), .D(n29[5]), .R(n2227));   // ../o_counter.v(71[46:63])
    SB_DFFESR FRAME_COUNTER_285__i1 (.Q(FRAME_COUNTER[1]), .C(TVP_CLK_c), 
            .E(n252), .D(n29[1]), .R(n2227));   // ../o_counter.v(71[46:63])
    SB_DFFSR X_284__i2 (.Q(n79[2]), .C(TVP_CLK_c), .D(n45[2]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_DFFSR X_284__i3 (.Q(X[3]), .C(TVP_CLK_c), .D(n45[3]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_DFFSR X_284__i4 (.Q(X[4]), .C(TVP_CLK_c), .D(n45[4]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_DFFSR X_284__i5 (.Q(X[5]), .C(TVP_CLK_c), .D(n45[5]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_DFFSR X_284__i6 (.Q(X[6]), .C(TVP_CLK_c), .D(n45[6]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_DFFSR X_284__i7 (.Q(X[7]), .C(TVP_CLK_c), .D(n45[7]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_DFFSR X_284__i8 (.Q(X[8]), .C(TVP_CLK_c), .D(n45[8]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_DFFSR X_284__i9 (.Q(X[9]), .C(TVP_CLK_c), .D(n45[9]), .R(n3184));   // ../o_counter.v(61[26:31])
    SB_LUT4 X_284_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(X[9]), 
            .I3(n2790), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 X_284_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(X[8]), 
            .I3(n2789), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_284_add_4_10 (.CI(n2789), .I0(GND_net), .I1(X[8]), .CO(n2790));
    SB_LUT4 X_284_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(X[7]), 
            .I3(n2788), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam X_284_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_284_add_4_9 (.CI(n2788), .I0(GND_net), .I1(X[7]), .CO(n2789));
    SB_LUT4 i873_2_lut_4_lut (.I0(FRAME_COUNTER[5]), .I1(n10_adj_570), .I2(FRAME_COUNTER[0]), 
            .I3(n252), .O(n2227));
    defparam i873_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_4_lut (.I0(FRAME_COUNTER[5]), .I1(n10_adj_570), .I2(FRAME_COUNTER[0]), 
            .I3(LED_c), .O(PULSE_1HZ_N_92));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdf20;
    
endmodule
//
// Verilog Description of module TX
//

module TX (DEBUG_c_3, GND_net, DEBUG_c_2, DEBUG_c_0, n28, ADV_CLK_c, 
           ADV_VSYNC_c, DEBUG_c_5, VGA_VISIBLE, n23, DEBUG_c_6, DEBUG_c_4, 
           n24, n18, n25, n19, n26, n20, DEBUG_c_1, n27, \TX_ADDR[11] , 
           DEBUG_c_7, n21, n22, \TX_ADDR[12] , \TX_ADDR[13] , VCC_net, 
           n2147, ADV_HSYNC_c, n5, n3009, \Y[1] , \Y[0] ) /* synthesis syn_module_defined=1 */ ;
    output DEBUG_c_3;
    input GND_net;
    output DEBUG_c_2;
    output DEBUG_c_0;
    output n28;
    input ADV_CLK_c;
    output ADV_VSYNC_c;
    output DEBUG_c_5;
    output VGA_VISIBLE;
    output n23;
    output DEBUG_c_6;
    output DEBUG_c_4;
    output n24;
    output n18;
    output n25;
    output n19;
    output n26;
    output n20;
    output DEBUG_c_1;
    output n27;
    output \TX_ADDR[11] ;
    output DEBUG_c_7;
    output n21;
    output n22;
    output \TX_ADDR[12] ;
    output \TX_ADDR[13] ;
    input VCC_net;
    output n2147;
    output ADV_HSYNC_c;
    input n5;
    input n3009;
    input \Y[1] ;
    input \Y[0] ;
    
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    
    wire n2742, n2743;
    wire [13:0]n374;
    
    wire n2741;
    wire [15:0]X_DELTA_PATTERN;   // ../tx.v(59[16:31])
    
    wire n2740, n2745;
    wire [13:0]TX_ADDR;   // ../main.v(45[14:21])
    
    wire n2746, n2744, n2748, n2749, n2200, n2747, n2752, n2751, 
        n2750;
    
    SB_CARRY add_15_5 (.CI(n2742), .I0(DEBUG_c_3), .I1(GND_net), .CO(n2743));
    SB_LUT4 add_15_4_lut (.I0(GND_net), .I1(DEBUG_c_2), .I2(GND_net), 
            .I3(n2741), .O(n374[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_15_2 (.CI(GND_net), .I0(DEBUG_c_0), .I1(X_DELTA_PATTERN[0]), 
            .CO(n2740));
    SB_DFF BRAM_ADDR__i1 (.Q(DEBUG_c_0), .C(ADV_CLK_c), .D(n28));   // ../tx.v(65[12] 88[8])
    SB_LUT4 i1057_4_lut (.I0(n374[5]), .I1(ADV_VSYNC_c), .I2(DEBUG_c_5), 
            .I3(VGA_VISIBLE), .O(n23));   // ../tx.v(65[12] 88[8])
    defparam i1057_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_15_8_lut (.I0(GND_net), .I1(DEBUG_c_6), .I2(GND_net), 
            .I3(n2745), .O(n374[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1058_4_lut (.I0(n374[4]), .I1(ADV_VSYNC_c), .I2(DEBUG_c_4), 
            .I3(VGA_VISIBLE), .O(n24));   // ../tx.v(65[12] 88[8])
    defparam i1058_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1052_4_lut (.I0(n374[10]), .I1(ADV_VSYNC_c), .I2(TX_ADDR[10]), 
            .I3(VGA_VISIBLE), .O(n18));   // ../tx.v(65[12] 88[8])
    defparam i1052_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1059_4_lut (.I0(n374[3]), .I1(ADV_VSYNC_c), .I2(DEBUG_c_3), 
            .I3(VGA_VISIBLE), .O(n25));   // ../tx.v(65[12] 88[8])
    defparam i1059_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1053_4_lut (.I0(n374[9]), .I1(ADV_VSYNC_c), .I2(TX_ADDR[9]), 
            .I3(VGA_VISIBLE), .O(n19));   // ../tx.v(65[12] 88[8])
    defparam i1053_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_15_8 (.CI(n2745), .I0(DEBUG_c_6), .I1(GND_net), .CO(n2746));
    SB_LUT4 i1060_4_lut (.I0(n374[2]), .I1(ADV_VSYNC_c), .I2(DEBUG_c_2), 
            .I3(VGA_VISIBLE), .O(n26));   // ../tx.v(65[12] 88[8])
    defparam i1060_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_15_7_lut (.I0(GND_net), .I1(DEBUG_c_5), .I2(GND_net), 
            .I3(n2744), .O(n374[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1054_4_lut (.I0(n374[8]), .I1(ADV_VSYNC_c), .I2(TX_ADDR[8]), 
            .I3(VGA_VISIBLE), .O(n20));   // ../tx.v(65[12] 88[8])
    defparam i1054_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1096_4_lut (.I0(n374[0]), .I1(ADV_VSYNC_c), .I2(DEBUG_c_0), 
            .I3(VGA_VISIBLE), .O(n28));   // ../tx.v(65[12] 88[8])
    defparam i1096_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1061_4_lut (.I0(n374[1]), .I1(ADV_VSYNC_c), .I2(DEBUG_c_1), 
            .I3(VGA_VISIBLE), .O(n27));   // ../tx.v(65[12] 88[8])
    defparam i1061_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_15_11 (.CI(n2748), .I0(TX_ADDR[9]), .I1(GND_net), .CO(n2749));
    SB_CARRY add_15_7 (.CI(n2744), .I0(DEBUG_c_5), .I1(GND_net), .CO(n2745));
    SB_CARRY add_15_4 (.CI(n2741), .I0(DEBUG_c_2), .I1(GND_net), .CO(n2742));
    SB_DFFESS X_DELTA_PATTERN_i0 (.Q(X_DELTA_PATTERN[0]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[1]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESR BRAM_ADDR__rep_1_i0 (.Q(\TX_ADDR[11] ), .C(ADV_CLK_c), .E(n2200), 
            .D(n374[11]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_LUT4 add_15_10_lut (.I0(GND_net), .I1(TX_ADDR[8]), .I2(GND_net), 
            .I3(n2747), .O(n374[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_15_6_lut (.I0(GND_net), .I1(DEBUG_c_4), .I2(GND_net), 
            .I3(n2743), .O(n374[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_15_3_lut (.I0(GND_net), .I1(DEBUG_c_1), .I2(GND_net), 
            .I3(n2740), .O(n374[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1055_4_lut (.I0(n374[7]), .I1(ADV_VSYNC_c), .I2(DEBUG_c_7), 
            .I3(VGA_VISIBLE), .O(n21));   // ../tx.v(65[12] 88[8])
    defparam i1055_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1056_4_lut (.I0(n374[6]), .I1(ADV_VSYNC_c), .I2(DEBUG_c_6), 
            .I3(VGA_VISIBLE), .O(n22));   // ../tx.v(65[12] 88[8])
    defparam i1056_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_15_10 (.CI(n2747), .I0(TX_ADDR[8]), .I1(GND_net), .CO(n2748));
    SB_LUT4 add_15_9_lut (.I0(GND_net), .I1(DEBUG_c_7), .I2(GND_net), 
            .I3(n2746), .O(n374[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_15_9 (.CI(n2746), .I0(DEBUG_c_7), .I1(GND_net), .CO(n2747));
    SB_CARRY add_15_3 (.CI(n2740), .I0(DEBUG_c_1), .I1(GND_net), .CO(n2741));
    SB_LUT4 i1_2_lut (.I0(VGA_VISIBLE), .I1(ADV_VSYNC_c), .I2(GND_net), 
            .I3(GND_net), .O(n2200));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFESR X_DELTA_PATTERN_i1 (.Q(X_DELTA_PATTERN[1]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[2]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_CARRY add_15_6 (.CI(n2743), .I0(DEBUG_c_4), .I1(GND_net), .CO(n2744));
    SB_LUT4 add_15_5_lut (.I0(GND_net), .I1(DEBUG_c_3), .I2(GND_net), 
            .I3(n2742), .O(n374[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_15_2_lut (.I0(GND_net), .I1(DEBUG_c_0), .I2(X_DELTA_PATTERN[0]), 
            .I3(GND_net), .O(n374[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR X_DELTA_PATTERN_i3 (.Q(X_DELTA_PATTERN[3]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[4]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESR X_DELTA_PATTERN_i5 (.Q(X_DELTA_PATTERN[5]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[6]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESR X_DELTA_PATTERN_i8 (.Q(X_DELTA_PATTERN[8]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[9]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESR X_DELTA_PATTERN_i10 (.Q(X_DELTA_PATTERN[10]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[11]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESR X_DELTA_PATTERN_i12 (.Q(X_DELTA_PATTERN[12]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[13]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESR X_DELTA_PATTERN_i14 (.Q(X_DELTA_PATTERN[14]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[15]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i2 (.Q(DEBUG_c_1), .C(ADV_CLK_c), .D(n27));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i3 (.Q(DEBUG_c_2), .C(ADV_CLK_c), .D(n26));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i4 (.Q(DEBUG_c_3), .C(ADV_CLK_c), .D(n25));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i5 (.Q(DEBUG_c_4), .C(ADV_CLK_c), .D(n24));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i6 (.Q(DEBUG_c_5), .C(ADV_CLK_c), .D(n23));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i7 (.Q(DEBUG_c_6), .C(ADV_CLK_c), .D(n22));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i8 (.Q(DEBUG_c_7), .C(ADV_CLK_c), .D(n21));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i9 (.Q(TX_ADDR[8]), .C(ADV_CLK_c), .D(n20));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i10 (.Q(TX_ADDR[9]), .C(ADV_CLK_c), .D(n19));   // ../tx.v(65[12] 88[8])
    SB_DFF BRAM_ADDR__i11 (.Q(TX_ADDR[10]), .C(ADV_CLK_c), .D(n18));   // ../tx.v(65[12] 88[8])
    SB_DFFESR BRAM_ADDR__rep_1_i1 (.Q(\TX_ADDR[12] ), .C(ADV_CLK_c), .E(n2200), 
            .D(n374[12]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESR BRAM_ADDR__rep_1_i2 (.Q(\TX_ADDR[13] ), .C(ADV_CLK_c), .E(n2200), 
            .D(n374[13]), .R(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESS X_DELTA_PATTERN_i15 (.Q(X_DELTA_PATTERN[15]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[0]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESS X_DELTA_PATTERN_i13 (.Q(X_DELTA_PATTERN[13]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[14]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESS X_DELTA_PATTERN_i11 (.Q(X_DELTA_PATTERN[11]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[12]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_LUT4 add_15_15_lut (.I0(GND_net), .I1(\TX_ADDR[13] ), .I2(GND_net), 
            .I3(n2752), .O(n374[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_15_14_lut (.I0(GND_net), .I1(\TX_ADDR[12] ), .I2(GND_net), 
            .I3(n2751), .O(n374[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_15_14 (.CI(n2751), .I0(\TX_ADDR[12] ), .I1(GND_net), 
            .CO(n2752));
    SB_LUT4 add_15_13_lut (.I0(GND_net), .I1(\TX_ADDR[11] ), .I2(GND_net), 
            .I3(n2750), .O(n374[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_15_13 (.CI(n2750), .I0(\TX_ADDR[11] ), .I1(GND_net), 
            .CO(n2751));
    SB_DFFESS X_DELTA_PATTERN_i9 (.Q(X_DELTA_PATTERN[9]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[10]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_LUT4 add_15_12_lut (.I0(GND_net), .I1(TX_ADDR[10]), .I2(GND_net), 
            .I3(n2749), .O(n374[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS X_DELTA_PATTERN_i7 (.Q(X_DELTA_PATTERN[7]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[8]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESS X_DELTA_PATTERN_i6 (.Q(X_DELTA_PATTERN[6]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[7]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_CARRY add_15_12 (.CI(n2749), .I0(TX_ADDR[10]), .I1(GND_net), .CO(n2750));
    SB_DFFESS X_DELTA_PATTERN_i4 (.Q(X_DELTA_PATTERN[4]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[5]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_DFFESS X_DELTA_PATTERN_i2 (.Q(X_DELTA_PATTERN[2]), .C(ADV_CLK_c), 
            .E(n2200), .D(X_DELTA_PATTERN[3]), .S(ADV_VSYNC_c));   // ../tx.v(65[12] 88[8])
    SB_LUT4 add_15_11_lut (.I0(GND_net), .I1(TX_ADDR[9]), .I2(GND_net), 
            .I3(n2748), .O(n374[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_15_11_lut.LUT_INIT = 16'hC33C;
    VGA_CONTROL video_signal_controller (.GND_net(GND_net), .VCC_net(VCC_net), 
            .ADV_CLK_c(ADV_CLK_c), .n2147(n2147), .ADV_VSYNC_c(ADV_VSYNC_c), 
            .ADV_HSYNC_c(ADV_HSYNC_c), .n5(n5), .n3009(n3009), .\Y[1] (\Y[1] ), 
            .\Y[0] (\Y[0] ), .VGA_VISIBLE(VGA_VISIBLE)) /* synthesis syn_module_defined=1 */ ;   // ../tx.v(41[17] 53[67])
    
endmodule
//
// Verilog Description of module VGA_CONTROL
//

module VGA_CONTROL (GND_net, VCC_net, ADV_CLK_c, n2147, ADV_VSYNC_c, 
            ADV_HSYNC_c, n5, n3009, \Y[1] , \Y[0] , VGA_VISIBLE) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input ADV_CLK_c;
    output n2147;
    output ADV_VSYNC_c;
    output ADV_HSYNC_c;
    input n5;
    input n3009;
    input \Y[1] ;
    input \Y[0] ;
    output VGA_VISIBLE;
    
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    
    wire n2776;
    wire [11:0]VGA_Y;   // ../vga_control.v(52[23:28])
    
    wire n2777;
    wire [6:0]n33;
    wire [10:0]n49;
    wire [11:0]VGA_X;   // ../vga_control.v(52[16:21])
    
    wire VGA_VS_N_552, VGA_HS_N_549, n2775, n2774, n2773, n2772, 
        n2771, n2770, n2769, n2768, n6, n3183, VGA_VISIBLE_N_558, 
        n2767, n2766, n2778, n2779, n2780, n2781, n2972, n12, 
        n3014, n3186, n3022, n3182, n8, n18, n2484, n2262;
    
    SB_CARRY VGA_Y_286_287_add_4_3 (.CI(n2776), .I0(GND_net), .I1(VGA_Y[1]), 
            .CO(n2777));
    SB_LUT4 VGA_Y_286_287_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_286_287_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR VGA_X_288_289__i1 (.Q(VGA_X[0]), .C(ADV_CLK_c), .D(n49[0]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_CARRY VGA_Y_286_287_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(VGA_Y[0]), 
            .CO(n2776));
    SB_DFF VGA_VS_49 (.Q(ADV_VSYNC_c), .C(ADV_CLK_c), .D(VGA_VS_N_552));   // ../vga_control.v(67[12] 90[8])
    SB_DFF VGA_HS_48 (.Q(ADV_HSYNC_c), .C(ADV_CLK_c), .D(VGA_HS_N_549));   // ../vga_control.v(67[12] 90[8])
    SB_LUT4 VGA_X_288_289_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[10]), 
            .I3(n2775), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 VGA_X_288_289_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[9]), 
            .I3(n2774), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_11 (.CI(n2774), .I0(GND_net), .I1(VGA_X[9]), 
            .CO(n2775));
    SB_LUT4 VGA_X_288_289_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[8]), 
            .I3(n2773), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_10 (.CI(n2773), .I0(GND_net), .I1(VGA_X[8]), 
            .CO(n2774));
    SB_LUT4 VGA_X_288_289_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[7]), 
            .I3(n2772), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_9 (.CI(n2772), .I0(GND_net), .I1(VGA_X[7]), 
            .CO(n2773));
    SB_LUT4 VGA_X_288_289_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[6]), 
            .I3(n2771), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_8 (.CI(n2771), .I0(GND_net), .I1(VGA_X[6]), 
            .CO(n2772));
    SB_LUT4 VGA_X_288_289_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[5]), 
            .I3(n2770), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_7 (.CI(n2770), .I0(GND_net), .I1(VGA_X[5]), 
            .CO(n2771));
    SB_LUT4 VGA_X_288_289_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[4]), 
            .I3(n2769), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_6 (.CI(n2769), .I0(GND_net), .I1(VGA_X[4]), 
            .CO(n2770));
    SB_LUT4 VGA_X_288_289_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[3]), 
            .I3(n2768), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i508_2_lut (.I0(VGA_Y[1]), .I1(VGA_Y[2]), .I2(GND_net), .I3(GND_net), 
            .O(n6));
    defparam i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY VGA_X_288_289_add_4_5 (.CI(n2768), .I0(GND_net), .I1(VGA_X[3]), 
            .CO(n2769));
    SB_LUT4 i1_4_lut (.I0(n6), .I1(n3183), .I2(VGA_Y[4]), .I3(VGA_Y[3]), 
            .O(VGA_VISIBLE_N_558));
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 VGA_X_288_289_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[2]), 
            .I3(n2767), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_4 (.CI(n2767), .I0(GND_net), .I1(VGA_X[2]), 
            .CO(n2768));
    SB_LUT4 VGA_X_288_289_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[1]), 
            .I3(n2766), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_3 (.CI(n2766), .I0(GND_net), .I1(VGA_X[1]), 
            .CO(n2767));
    SB_LUT4 VGA_X_288_289_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_288_289_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_288_289_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(VGA_X[0]), 
            .CO(n2766));
    SB_LUT4 VGA_Y_286_287_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[1]), 
            .I3(n2776), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_286_287_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_286_287_add_4_4 (.CI(n2777), .I0(GND_net), .I1(VGA_Y[2]), 
            .CO(n2778));
    SB_LUT4 VGA_Y_286_287_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[2]), 
            .I3(n2777), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_286_287_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_286_287_add_4_5 (.CI(n2778), .I0(GND_net), .I1(VGA_Y[3]), 
            .CO(n2779));
    SB_LUT4 VGA_Y_286_287_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[3]), 
            .I3(n2778), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_286_287_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_286_287_add_4_6 (.CI(n2779), .I0(GND_net), .I1(VGA_Y[4]), 
            .CO(n2780));
    SB_LUT4 VGA_Y_286_287_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[4]), 
            .I3(n2779), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_286_287_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_286_287_add_4_7 (.CI(n2780), .I0(GND_net), .I1(VGA_Y[5]), 
            .CO(n2781));
    SB_LUT4 i2_3_lut (.I0(VGA_X[5]), .I1(VGA_X[6]), .I2(VGA_X[4]), .I3(GND_net), 
            .O(n2972));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i541_3_lut (.I0(VGA_X[3]), .I1(VGA_X[5]), .I2(VGA_X[4]), .I3(GND_net), 
            .O(n12));
    defparam i541_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1570_4_lut (.I0(n2972), .I1(VGA_X[9]), .I2(VGA_X[7]), .I3(VGA_X[10]), 
            .O(n3014));
    defparam i1570_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i1629_4_lut (.I0(n3186), .I1(n3014), .I2(VGA_X[8]), .I3(n12), 
            .O(VGA_HS_N_549));   // ../vga_control.v(69[19:88])
    defparam i1629_4_lut.LUT_INIT = 16'hfcfd;
    SB_LUT4 i4_4_lut (.I0(VGA_Y[0]), .I1(n3022), .I2(VGA_Y[2]), .I3(VGA_Y[1]), 
            .O(VGA_VS_N_552));
    defparam i4_4_lut.LUT_INIT = 16'h0302;
    SB_DFFSR VGA_X_288_289__i2 (.Q(VGA_X[1]), .C(ADV_CLK_c), .D(n49[1]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_LUT4 i1_2_lut_rep_18_3_lut (.I0(VGA_X[7]), .I1(VGA_X[6]), .I2(VGA_X[5]), 
            .I3(GND_net), .O(n3182));
    defparam i1_2_lut_rep_18_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_3_lut (.I0(VGA_X[4]), .I1(VGA_X[3]), .I2(VGA_X[2]), .I3(GND_net), 
            .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_DFFSR VGA_X_288_289__i3 (.Q(VGA_X[2]), .C(ADV_CLK_c), .D(n49[2]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_DFFSR VGA_X_288_289__i4 (.Q(VGA_X[3]), .C(ADV_CLK_c), .D(n49[3]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_DFFSR VGA_X_288_289__i5 (.Q(VGA_X[4]), .C(ADV_CLK_c), .D(n49[4]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_DFFSR VGA_X_288_289__i6 (.Q(VGA_X[5]), .C(ADV_CLK_c), .D(n49[5]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_DFFSR VGA_X_288_289__i7 (.Q(VGA_X[6]), .C(ADV_CLK_c), .D(n49[6]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_DFFSR VGA_X_288_289__i8 (.Q(VGA_X[7]), .C(ADV_CLK_c), .D(n49[7]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_DFFSR VGA_X_288_289__i9 (.Q(VGA_X[8]), .C(ADV_CLK_c), .D(n49[8]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_DFFSR VGA_X_288_289__i10 (.Q(VGA_X[9]), .C(ADV_CLK_c), .D(n49[9]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_DFFSR VGA_X_288_289__i11 (.Q(VGA_X[10]), .C(ADV_CLK_c), .D(n49[10]), 
            .R(n2147));   // ../vga_control.v(75[26:35])
    SB_LUT4 i511_2_lut_3_lut_4_lut (.I0(VGA_X[7]), .I1(VGA_X[6]), .I2(VGA_X[8]), 
            .I3(VGA_X[5]), .O(n18));
    defparam i511_2_lut_3_lut_4_lut.LUT_INIT = 16'hf0e0;
    SB_LUT4 i1_2_lut_rep_22 (.I0(VGA_X[7]), .I1(VGA_X[6]), .I2(GND_net), 
            .I3(GND_net), .O(n3186));
    defparam i1_2_lut_rep_22.LUT_INIT = 16'heeee;
    SB_LUT4 i1127_4_lut (.I0(VGA_X[0]), .I1(n3182), .I2(n8), .I3(VGA_X[1]), 
            .O(n2484));
    defparam i1127_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1642_4_lut (.I0(n5), .I1(n3009), .I2(\Y[1] ), .I3(\Y[0] ), 
            .O(n2262));
    defparam i1642_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1145_4_lut (.I0(n2484), .I1(VGA_X[10]), .I2(VGA_X[9]), .I3(VGA_X[8]), 
            .O(n2147));
    defparam i1145_4_lut.LUT_INIT = 16'hc8c0;
    SB_DFFESR VGA_Y_286_287__i1 (.Q(VGA_Y[0]), .C(ADV_CLK_c), .E(n2147), 
            .D(n33[0]), .R(n2262));   // ../vga_control.v(81[30:39])
    SB_LUT4 VGA_Y_286_287_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[5]), 
            .I3(n2780), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_286_287_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR VGA_Y_286_287__i7 (.Q(VGA_Y[6]), .C(ADV_CLK_c), .E(n2147), 
            .D(n33[6]), .R(n2262));   // ../vga_control.v(81[30:39])
    SB_LUT4 VGA_Y_286_287_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[6]), 
            .I3(n2781), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_286_287_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1578_3_lut_4_lut (.I0(VGA_Y[6]), .I1(VGA_Y[5]), .I2(VGA_Y[3]), 
            .I3(VGA_Y[4]), .O(n3022));
    defparam i1578_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR VGA_Y_286_287__i6 (.Q(VGA_Y[5]), .C(ADV_CLK_c), .E(n2147), 
            .D(n33[5]), .R(n2262));   // ../vga_control.v(81[30:39])
    SB_DFFESR VGA_Y_286_287__i5 (.Q(VGA_Y[4]), .C(ADV_CLK_c), .E(n2147), 
            .D(n33[4]), .R(n2262));   // ../vga_control.v(81[30:39])
    SB_DFFESR VGA_Y_286_287__i4 (.Q(VGA_Y[3]), .C(ADV_CLK_c), .E(n2147), 
            .D(n33[3]), .R(n2262));   // ../vga_control.v(81[30:39])
    SB_DFFESR VGA_Y_286_287__i3 (.Q(VGA_Y[2]), .C(ADV_CLK_c), .E(n2147), 
            .D(n33[2]), .R(n2262));   // ../vga_control.v(81[30:39])
    SB_DFFESR VGA_Y_286_287__i2 (.Q(VGA_Y[1]), .C(ADV_CLK_c), .E(n2147), 
            .D(n33[1]), .R(n2262));   // ../vga_control.v(81[30:39])
    SB_LUT4 i1_2_lut_rep_19 (.I0(VGA_Y[6]), .I1(VGA_Y[5]), .I2(GND_net), 
            .I3(GND_net), .O(n3183));
    defparam i1_2_lut_rep_19.LUT_INIT = 16'heeee;
    SB_LUT4 i1636_4_lut_4_lut (.I0(n18), .I1(VGA_VISIBLE_N_558), .I2(VGA_X[10]), 
            .I3(VGA_X[9]), .O(VGA_VISIBLE));   // ../vga_control.v(54[26:180])
    defparam i1636_4_lut_4_lut.LUT_INIT = 16'hf3b7;
    
endmodule
//
// Verilog Description of module TX_PLL
//

module TX_PLL (TVP_CLK_c, VCC_net, GND_net, ADV_CLK_c) /* synthesis syn_module_defined=1 */ ;
    input TVP_CLK_c;
    input VCC_net;
    input GND_net;
    output ADV_CLK_c;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    
    SB_PLL40_CORE TX_PLL_inst (.REFERENCECLK(TVP_CLK_c), .PLLOUTCORE(ADV_CLK_c), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=13, LSE_LCOL=9, LSE_RCOL=25, LSE_LLINE=20, LSE_RLINE=24 */ ;   // ../main.v(20[9] 24[25])
    defparam TX_PLL_inst.FEEDBACK_PATH = "SIMPLE";
    defparam TX_PLL_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam TX_PLL_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam TX_PLL_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam TX_PLL_inst.FDA_FEEDBACK = 4'b0000;
    defparam TX_PLL_inst.FDA_RELATIVE = 4'b0000;
    defparam TX_PLL_inst.PLLOUT_SELECT = "GENCLK";
    defparam TX_PLL_inst.DIVR = 4'b0000;
    defparam TX_PLL_inst.DIVF = 7'b0100110;
    defparam TX_PLL_inst.DIVQ = 3'b100;
    defparam TX_PLL_inst.FILTER_RANGE = 3'b010;
    defparam TX_PLL_inst.ENABLE_ICEGATE = 1'b0;
    defparam TX_PLL_inst.TEST_MODE = 1'b0;
    defparam TX_PLL_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module RAM
//

module RAM (TX_DATA, ADV_CLK_c, \TX_ADDR[12] , n25, RX_ADDR, \TX_ADDR[13] , 
            GND_net, \TX_ADDR[11] , n28, n27, n26, n25_adj_1, n24, 
            n23, n22, n21, n20, n19, n18, TVP_VIDEO_c_8, TVP_VIDEO_c_9, 
            TVP_CLK_c, VCC_net, TVP_VIDEO_c_6, TVP_VIDEO_c_7, TVP_VIDEO_c_4, 
            TVP_VIDEO_c_5, TVP_VIDEO_c_2, TVP_VIDEO_c_3) /* synthesis syn_module_defined=1 */ ;
    output [7:0]TX_DATA;
    input ADV_CLK_c;
    input \TX_ADDR[12] ;
    input n25;
    input [13:0]RX_ADDR;
    input \TX_ADDR[13] ;
    input GND_net;
    input \TX_ADDR[11] ;
    input n28;
    input n27;
    input n26;
    input n25_adj_1;
    input n24;
    input n23;
    input n22;
    input n21;
    input n20;
    input n19;
    input n18;
    input TVP_VIDEO_c_8;
    input TVP_VIDEO_c_9;
    input TVP_CLK_c;
    input VCC_net;
    input TVP_VIDEO_c_6;
    input TVP_VIDEO_c_7;
    input TVP_VIDEO_c_4;
    input TVP_VIDEO_c_5;
    input TVP_VIDEO_c_2;
    input TVP_VIDEO_c_3;
    
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire [7:0]dout_7__N_561;
    
    wire n3107, n624, n616, n3110, n730, n3116, n3122, n750, 
        n758, n3101, n718, n726, n3161, n629, n621, n3164, n749, 
        n757, n3155, n693, n685, n3158, n686, n687, n697, n619, 
        n620, n632, n617, n618, n717, n725, n3149, n615, n628, 
        n3152, n684, n719, n729, n682, n683, n680, n681, n716, 
        n630, n633, n714, n715, n712, n713, n627, n751, n761, 
        n625, n626, n623, n748, n694, n695, n698, n746, n747, 
        n744, n745, n692, n727, n690, n691, n688, n689, n724, 
        n759, n762, n722, n723, n720, n721, n756, n622, n754, 
        n755, n752, n753, n3143, n3146, n3137, n3140, n3024, 
        n3025, n3131, n3046, n3045, n3027, n3028, n3125, n3043, 
        n3042, n3119, n3113, n3104, n3030, n3031, n3095, n3040, 
        n3039, n3089, n3092;
    
    SB_DFF dout_i0 (.Q(TX_DATA[0]), .C(ADV_CLK_c), .D(dout_7__N_561[0]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 n3107_bdd_4_lut (.I0(n3107), .I1(n624), .I2(n616), .I3(\TX_ADDR[12] ), 
            .O(n3110));
    defparam n3107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n25), .I1(RX_ADDR[13]), .I2(RX_ADDR[12]), 
            .I3(RX_ADDR[11]), .O(n730));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i115911_i1_3_lut (.I0(n3116), .I1(n3122), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_561[0]));
    defparam i115911_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1661 (.I0(\TX_ADDR[11] ), .I1(n750), .I2(n758), 
            .I3(\TX_ADDR[12] ), .O(n3101));
    defparam TX_ADDR_11__bdd_4_lut_1661.LUT_INIT = 16'he4aa;
    SB_LUT4 TX_ADDR_11__bdd_4_lut (.I0(\TX_ADDR[11] ), .I1(n718), .I2(n726), 
            .I3(\TX_ADDR[12] ), .O(n3161));
    defparam TX_ADDR_11__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n3161_bdd_4_lut (.I0(n3161), .I1(n629), .I2(n621), .I3(\TX_ADDR[12] ), 
            .O(n3164));
    defparam n3161_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1706 (.I0(\TX_ADDR[11] ), .I1(n749), .I2(n757), 
            .I3(\TX_ADDR[12] ), .O(n3155));
    defparam TX_ADDR_11__bdd_4_lut_1706.LUT_INIT = 16'he4aa;
    SB_LUT4 n3155_bdd_4_lut (.I0(n3155), .I1(n693), .I2(n685), .I3(\TX_ADDR[12] ), 
            .O(n3158));
    defparam n3155_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_RAM2048x2 mem0 (.RDATA({n687, n686}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n697), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem0.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem8 (.RDATA({n620, n619}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n632), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem8.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem9 (.RDATA({n618, n617}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n632), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem9.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1701 (.I0(\TX_ADDR[11] ), .I1(n717), .I2(n725), 
            .I3(\TX_ADDR[12] ), .O(n3149));
    defparam TX_ADDR_11__bdd_4_lut_1701.LUT_INIT = 16'he4aa;
    SB_RAM2048x2 mem10 (.RDATA({n616, n615}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n632), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem10.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 n3149_bdd_4_lut (.I0(n3149), .I1(n628), .I2(n620), .I3(\TX_ADDR[12] ), 
            .O(n3152));
    defparam n3149_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_RAM2048x2 mem11 (.RDATA({n685, n684}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n697), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem11.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem1 (.RDATA({n719, n718}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n729), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem1.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem12 (.RDATA({n683, n682}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n697), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem13 (.RDATA({n681, n680}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n697), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem13.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem14 (.RDATA({n717, n716}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n729), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem14.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem2 (.RDATA({n630, n629}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n633), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem2.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem15 (.RDATA({n715, n714}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n729), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem15.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem16 (.RDATA({n713, n712}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n729), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem16.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem17 (.RDATA({n628, n627}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n633), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem17.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem3 (.RDATA({n751, n750}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n761), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem3.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem18 (.RDATA({n626, n625}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n633), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem18.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem19 (.RDATA({n624, n623}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n633), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem19.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem20 (.RDATA({n749, n748}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n761), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem20.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem4 (.RDATA({n695, n694}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n698), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem4.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem21 (.RDATA({n747, n746}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n761), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem21.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem22 (.RDATA({n745, n744}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n761), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem22.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem23 (.RDATA({n693, n692}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n698), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem23.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem5 (.RDATA({n727, n726}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n730), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem5.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem24 (.RDATA({n691, n690}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n698), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem24.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem25 (.RDATA({n689, n688}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n698), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem25.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem26 (.RDATA({n725, n724}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n730), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem26.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem6 (.RDATA({n759, n758}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n762), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem6.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem27 (.RDATA({n723, n722}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n730), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem27.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem28 (.RDATA({n721, n720}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n730), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem28.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem29 (.RDATA({n757, n756}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n762), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem29.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem7 (.RDATA({n622, n621}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n632), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem7.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem30 (.RDATA({n755, n754}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n762), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem30.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem31 (.RDATA({n753, n752}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25_adj_1, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n762), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem31.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1696 (.I0(\TX_ADDR[11] ), .I1(n746), .I2(n754), 
            .I3(\TX_ADDR[12] ), .O(n3143));
    defparam TX_ADDR_11__bdd_4_lut_1696.LUT_INIT = 16'he4aa;
    SB_LUT4 n3143_bdd_4_lut (.I0(n3143), .I1(n690), .I2(n682), .I3(\TX_ADDR[12] ), 
            .O(n3146));
    defparam n3143_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1691 (.I0(\TX_ADDR[11] ), .I1(n745), .I2(n753), 
            .I3(\TX_ADDR[12] ), .O(n3137));
    defparam TX_ADDR_11__bdd_4_lut_1691.LUT_INIT = 16'he4aa;
    SB_LUT4 n3137_bdd_4_lut (.I0(n3137), .I1(n689), .I2(n681), .I3(\TX_ADDR[12] ), 
            .O(n3140));
    defparam n3137_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_12__bdd_4_lut (.I0(\TX_ADDR[12] ), .I1(n3024), .I2(n3025), 
            .I3(\TX_ADDR[13] ), .O(n3131));
    defparam TX_ADDR_12__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n3131_bdd_4_lut (.I0(n3131), .I1(n3046), .I2(n3045), .I3(\TX_ADDR[13] ), 
            .O(dout_7__N_561[4]));
    defparam n3131_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_12__bdd_4_lut_1681 (.I0(\TX_ADDR[12] ), .I1(n3027), 
            .I2(n3028), .I3(\TX_ADDR[13] ), .O(n3125));
    defparam TX_ADDR_12__bdd_4_lut_1681.LUT_INIT = 16'he4aa;
    SB_LUT4 n3125_bdd_4_lut (.I0(n3125), .I1(n3043), .I2(n3042), .I3(\TX_ADDR[13] ), 
            .O(dout_7__N_561[7]));
    defparam n3125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1686 (.I0(\TX_ADDR[11] ), .I1(n744), .I2(n752), 
            .I3(\TX_ADDR[12] ), .O(n3119));
    defparam TX_ADDR_11__bdd_4_lut_1686.LUT_INIT = 16'he4aa;
    SB_LUT4 n3119_bdd_4_lut (.I0(n3119), .I1(n688), .I2(n680), .I3(\TX_ADDR[12] ), 
            .O(n3122));
    defparam n3119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1671 (.I0(\TX_ADDR[11] ), .I1(n712), .I2(n720), 
            .I3(\TX_ADDR[12] ), .O(n3113));
    defparam TX_ADDR_11__bdd_4_lut_1671.LUT_INIT = 16'he4aa;
    SB_LUT4 n3113_bdd_4_lut (.I0(n3113), .I1(n623), .I2(n615), .I3(\TX_ADDR[12] ), 
            .O(n3116));
    defparam n3113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1666 (.I0(\TX_ADDR[11] ), .I1(n713), .I2(n721), 
            .I3(\TX_ADDR[12] ), .O(n3107));
    defparam TX_ADDR_11__bdd_4_lut_1666.LUT_INIT = 16'he4aa;
    SB_DFF dout_i1 (.Q(TX_DATA[1]), .C(ADV_CLK_c), .D(dout_7__N_561[1]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i2 (.Q(TX_DATA[2]), .C(ADV_CLK_c), .D(dout_7__N_561[2]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 n3101_bdd_4_lut (.I0(n3101), .I1(n694), .I2(n686), .I3(\TX_ADDR[12] ), 
            .O(n3104));
    defparam n3101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF dout_i3 (.Q(TX_DATA[3]), .C(ADV_CLK_c), .D(dout_7__N_561[3]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i4 (.Q(TX_DATA[4]), .C(ADV_CLK_c), .D(dout_7__N_561[4]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i5 (.Q(TX_DATA[5]), .C(ADV_CLK_c), .D(dout_7__N_561[5]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i6 (.Q(TX_DATA[6]), .C(ADV_CLK_c), .D(dout_7__N_561[6]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i7 (.Q(TX_DATA[7]), .C(ADV_CLK_c), .D(dout_7__N_561[7]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 TX_ADDR_12__bdd_4_lut_1676 (.I0(\TX_ADDR[12] ), .I1(n3030), 
            .I2(n3031), .I3(\TX_ADDR[13] ), .O(n3095));
    defparam TX_ADDR_12__bdd_4_lut_1676.LUT_INIT = 16'he4aa;
    SB_LUT4 n3095_bdd_4_lut (.I0(n3095), .I1(n3040), .I2(n3039), .I3(\TX_ADDR[13] ), 
            .O(dout_7__N_561[3]));
    defparam n3095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1595_3_lut (.I0(n618), .I1(n626), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3039));
    defparam i1595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_11 (.I0(n25), .I1(RX_ADDR[13]), .I2(RX_ADDR[12]), 
            .I3(RX_ADDR[11]), .O(n762));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_11.LUT_INIT = 16'h4000;
    SB_LUT4 i1596_3_lut (.I0(n715), .I1(n723), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3040));
    defparam i1596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1587_3_lut (.I0(n747), .I1(n755), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3031));
    defparam i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_12 (.I0(RX_ADDR[12]), .I1(RX_ADDR[11]), 
            .I2(RX_ADDR[13]), .I3(n25), .O(n697));
    defparam i1_2_lut_3_lut_4_lut_adj_12.LUT_INIT = 16'h0010;
    SB_LUT4 i1639_2_lut_3_lut_4_lut (.I0(RX_ADDR[12]), .I1(RX_ADDR[11]), 
            .I2(RX_ADDR[13]), .I3(n25), .O(n632));
    defparam i1639_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_1656 (.I0(\TX_ADDR[11] ), .I1(n714), .I2(n722), 
            .I3(\TX_ADDR[12] ), .O(n3089));
    defparam TX_ADDR_11__bdd_4_lut_1656.LUT_INIT = 16'he4aa;
    SB_LUT4 i1586_3_lut (.I0(n683), .I1(n691), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3030));
    defparam i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i119529_i1_3_lut (.I0(n3164), .I1(n3104), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_561[6]));
    defparam i119529_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n3089_bdd_4_lut (.I0(n3089), .I1(n625), .I2(n617), .I3(\TX_ADDR[12] ), 
            .O(n3092));
    defparam n3089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i118926_i1_3_lut (.I0(n3152), .I1(n3158), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_561[5]));
    defparam i118926_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i117117_i1_3_lut (.I0(n3092), .I1(n3146), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_561[2]));
    defparam i117117_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.I0(n25), .I1(RX_ADDR[13]), .I2(RX_ADDR[12]), 
            .I3(RX_ADDR[11]), .O(n698));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_13.LUT_INIT = 16'h0400;
    SB_LUT4 i116514_i1_3_lut (.I0(n3110), .I1(n3140), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_561[1]));
    defparam i116514_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_14 (.I0(RX_ADDR[12]), .I1(RX_ADDR[11]), 
            .I2(RX_ADDR[13]), .I3(n25), .O(n761));
    defparam i1_2_lut_3_lut_4_lut_adj_14.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_15 (.I0(RX_ADDR[12]), .I1(RX_ADDR[11]), 
            .I2(RX_ADDR[13]), .I3(n25), .O(n729));
    defparam i1_2_lut_3_lut_4_lut_adj_15.LUT_INIT = 16'h0002;
    SB_LUT4 i1598_3_lut (.I0(n622), .I1(n630), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3042));
    defparam i1598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1599_3_lut (.I0(n719), .I1(n727), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3043));
    defparam i1599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1584_3_lut (.I0(n751), .I1(n759), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3028));
    defparam i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1583_3_lut (.I0(n687), .I1(n695), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3027));
    defparam i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1601_3_lut (.I0(n619), .I1(n627), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3045));
    defparam i1601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1602_3_lut (.I0(n716), .I1(n724), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3046));
    defparam i1602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1581_3_lut (.I0(n748), .I1(n756), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3025));
    defparam i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1580_3_lut (.I0(n684), .I1(n692), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3024));
    defparam i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_16 (.I0(n25), .I1(RX_ADDR[13]), .I2(RX_ADDR[12]), 
            .I3(RX_ADDR[11]), .O(n633));
    defparam i1_2_lut_3_lut_4_lut_adj_16.LUT_INIT = 16'h0100;
    
endmodule
