-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 23 2018 02:41:33

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    TVP_VIDEO : in std_logic_vector(9 downto 0);
    ADV_B : out std_logic_vector(7 downto 0);
    ADV_G : out std_logic_vector(7 downto 0);
    ADV_R : out std_logic_vector(7 downto 0);
    DEBUG : inout std_logic_vector(7 downto 0);
    TVP_CLK : in std_logic;
    ADV_CLK : out std_logic;
    TVP_HSYNC : in std_logic;
    ADV_HSYNC : out std_logic;
    TVP_VSYNC : in std_logic;
    ADV_VSYNC : out std_logic;
    ADV_BLANK_N : out std_logic;
    LED : out std_logic;
    ADV_SYNC_N : out std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__10324\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \CLK_100MHz\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_38\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_79\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_40\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_39\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_41\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_82\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_81\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_80\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_86\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_90\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_89\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_85\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_88\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_87\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_84\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_83\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_92\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_91\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_97\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_98\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_93\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_96\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_95\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_94\ : std_logic;
signal \ADV_R_c_2\ : std_logic;
signal \ADV_R_c_0\ : std_logic;
signal \ADV_R_c_6\ : std_logic;
signal \INVADV_R__i3C_net\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_61\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_65\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_62\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_64\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_63\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_60\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_59\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_76\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_75\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_78\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_77\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_37\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_69\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_70\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_36\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_35\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_74\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_73\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_72\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_71\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_45\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_58\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_57\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_48\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_56\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_47\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_46\ : std_logic;
signal \transmit_module.n868\ : std_logic;
signal \transmit_module.video_signal_controller.SYNC_BUFF1\ : std_logic;
signal \DEBUG_c_7\ : std_logic;
signal \transmit_module.video_signal_controller.SYNC_BUFF2\ : std_logic;
signal \transmit_module.video_signal_controller.n2067_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n4\ : std_logic;
signal \transmit_module.video_signal_controller.SYNC_EN_SMOOTH\ : std_logic;
signal \transmit_module.video_signal_controller.n1983\ : std_logic;
signal \transmit_module.video_signal_controller.n2004_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n9\ : std_logic;
signal \transmit_module.video_signal_controller.n11\ : std_logic;
signal \transmit_module.video_signal_controller.n2121\ : std_logic;
signal \transmit_module.video_signal_controller.n7_cascade_\ : std_logic;
signal \bfn_3_21_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n1854\ : std_logic;
signal \transmit_module.video_signal_controller.n1855\ : std_logic;
signal \transmit_module.video_signal_controller.n1856\ : std_logic;
signal \transmit_module.video_signal_controller.n1857\ : std_logic;
signal \transmit_module.video_signal_controller.n1858\ : std_logic;
signal \transmit_module.video_signal_controller.n1859\ : std_logic;
signal \transmit_module.video_signal_controller.n1860\ : std_logic;
signal \transmit_module.video_signal_controller.n1861\ : std_logic;
signal \bfn_3_22_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n1862\ : std_logic;
signal \transmit_module.video_signal_controller.n1863\ : std_logic;
signal \transmit_module.video_signal_controller.n1864\ : std_logic;
signal \transmit_module.video_signal_controller.n1582\ : std_logic;
signal \ADV_G_c_6\ : std_logic;
signal \ADV_R_c_1\ : std_logic;
signal \INVADV_G__i7C_net\ : std_logic;
signal \receive_module.BRAM_ADDR_0\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal \receive_module.BRAM_ADDR_1\ : std_logic;
signal \receive_module.n1810\ : std_logic;
signal \receive_module.BRAM_ADDR_2\ : std_logic;
signal \receive_module.n1811\ : std_logic;
signal \receive_module.BRAM_ADDR_3\ : std_logic;
signal \receive_module.n1812\ : std_logic;
signal \receive_module.BRAM_ADDR_4\ : std_logic;
signal \receive_module.n1813\ : std_logic;
signal \receive_module.BRAM_ADDR_5\ : std_logic;
signal \receive_module.n1814\ : std_logic;
signal \receive_module.BRAM_ADDR_6\ : std_logic;
signal \receive_module.n1815\ : std_logic;
signal \receive_module.BRAM_ADDR_7\ : std_logic;
signal \receive_module.n1816\ : std_logic;
signal \receive_module.n1817\ : std_logic;
signal \receive_module.BRAM_ADDR_8\ : std_logic;
signal \bfn_4_8_0_\ : std_logic;
signal \receive_module.BRAM_ADDR_9\ : std_logic;
signal \receive_module.n1818\ : std_logic;
signal \receive_module.BRAM_ADDR_10\ : std_logic;
signal \receive_module.n1819\ : std_logic;
signal \receive_module.BRAM_ADDR_11\ : std_logic;
signal \receive_module.n1820\ : std_logic;
signal \receive_module.BRAM_ADDR_12\ : std_logic;
signal \receive_module.n1821\ : std_logic;
signal \receive_module.n1822\ : std_logic;
signal \DEBUG_c_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_34\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_68\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_67\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_66\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_53\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_55\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_54\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_44\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_49\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_43\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_42\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_52\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_51\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_50\ : std_logic;
signal \transmit_module.n2159\ : std_logic;
signal \transmit_module.video_signal_controller.n2079_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2117_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2154\ : std_logic;
signal \transmit_module.video_signal_controller.n12\ : std_logic;
signal \transmit_module.video_signal_controller.n2146_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n1769_cascade_\ : std_logic;
signal \transmit_module.n2147\ : std_logic;
signal \transmit_module.video_signal_controller.n18_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n8_adj_572\ : std_logic;
signal \ADV_R_c_5\ : std_logic;
signal \ADV_R_c_3\ : std_logic;
signal \ADV_B_c_5\ : std_logic;
signal \ADV_G_c_0\ : std_logic;
signal \ADV_R_c_4\ : std_logic;
signal \INVADV_R__i6C_net\ : std_logic;
signal \transmit_module.video_signal_controller.n2076\ : std_logic;
signal \transmit_module.video_signal_controller.n2011_cascade_\ : std_logic;
signal \transmit_module.n1997_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n18\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_9\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_8\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_11\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_10\ : std_logic;
signal \transmit_module.video_signal_controller.n679\ : std_logic;
signal \transmit_module.video_signal_controller.n679_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2151\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_552\ : std_logic;
signal \VGA_Y_5\ : std_logic;
signal \transmit_module.video_signal_controller.n2149_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2152\ : std_logic;
signal \transmit_module.video_signal_controller.n2006\ : std_logic;
signal \transmit_module.video_signal_controller.n8\ : std_logic;
signal \transmit_module.video_signal_controller.n2140\ : std_logic;
signal \ADV_G_c_3\ : std_logic;
signal \VGA_Y_3\ : std_logic;
signal \ADV_B_c_3\ : std_logic;
signal \INVADV_G__i4C_net\ : std_logic;
signal \DEBUG_c_5\ : std_logic;
signal \receive_module.rx_counter.n28_cascade_\ : std_logic;
signal \DEBUG_c_4\ : std_logic;
signal \DEBUG_c_4_cascade_\ : std_logic;
signal \receive_module.n788\ : std_logic;
signal \receive_module.rx_counter.n2083\ : std_logic;
signal \receive_module.rx_counter.n2033\ : std_logic;
signal \receive_module.rx_counter.n1981\ : std_logic;
signal \receive_module.rx_counter.n10\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \receive_module.rx_counter.n9\ : std_logic;
signal \receive_module.rx_counter.n1870\ : std_logic;
signal \receive_module.rx_counter.n8_adj_575\ : std_logic;
signal \receive_module.rx_counter.n1871\ : std_logic;
signal \receive_module.rx_counter.X_3\ : std_logic;
signal \receive_module.rx_counter.n1872\ : std_logic;
signal \receive_module.rx_counter.X_4\ : std_logic;
signal \receive_module.rx_counter.n1873\ : std_logic;
signal \receive_module.rx_counter.X_5\ : std_logic;
signal \receive_module.rx_counter.n1874\ : std_logic;
signal \receive_module.rx_counter.X_6\ : std_logic;
signal \receive_module.rx_counter.n1875\ : std_logic;
signal \receive_module.rx_counter.X_7\ : std_logic;
signal \receive_module.rx_counter.n1876\ : std_logic;
signal \receive_module.rx_counter.n1877\ : std_logic;
signal \receive_module.rx_counter.X_8\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \receive_module.rx_counter.n1878\ : std_logic;
signal \receive_module.rx_counter.X_9\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_4\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \transmit_module.n1823\ : std_logic;
signal \transmit_module.n1824\ : std_logic;
signal \transmit_module.n1825\ : std_logic;
signal \transmit_module.BRAM_ADDR_4\ : std_logic;
signal \transmit_module.n200\ : std_logic;
signal \transmit_module.n1826\ : std_logic;
signal \transmit_module.n1827\ : std_logic;
signal \transmit_module.n1828\ : std_logic;
signal \transmit_module.n1829\ : std_logic;
signal \transmit_module.n1830\ : std_logic;
signal \bfn_5_16_0_\ : std_logic;
signal \transmit_module.n1831\ : std_logic;
signal \transmit_module.n1832\ : std_logic;
signal \transmit_module.n1833\ : std_logic;
signal \transmit_module.n1834\ : std_logic;
signal \transmit_module.n1835\ : std_logic;
signal \transmit_module.n193\ : std_logic;
signal \transmit_module.n196\ : std_logic;
signal \transmit_module.n192\ : std_logic;
signal \transmit_module.n204\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_9\ : std_logic;
signal \transmit_module.n195\ : std_logic;
signal \transmit_module.BRAM_ADDR_9\ : std_logic;
signal \transmit_module.n194\ : std_logic;
signal \transmit_module.n202\ : std_logic;
signal \transmit_module.n2145_cascade_\ : std_logic;
signal n2144 : std_logic;
signal \transmit_module.old_VGA_HS\ : std_logic;
signal \ADV_HSYNC_c\ : std_logic;
signal \transmit_module.n2156_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_0\ : std_logic;
signal \bfn_5_19_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n1844\ : std_logic;
signal \transmit_module.video_signal_controller.n1845\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_3\ : std_logic;
signal \transmit_module.video_signal_controller.n1846\ : std_logic;
signal \transmit_module.video_signal_controller.n1847\ : std_logic;
signal \transmit_module.video_signal_controller.n1848\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_6\ : std_logic;
signal \transmit_module.video_signal_controller.n1849\ : std_logic;
signal \transmit_module.video_signal_controller.n1850\ : std_logic;
signal \transmit_module.video_signal_controller.n1851\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_8\ : std_logic;
signal \bfn_5_20_0_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_9\ : std_logic;
signal \transmit_module.video_signal_controller.n1852\ : std_logic;
signal \transmit_module.video_signal_controller.n1853\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_10\ : std_logic;
signal \transmit_module.video_signal_controller.n528\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_2\ : std_logic;
signal \ADV_G_c_2\ : std_logic;
signal \VGA_Y_4\ : std_logic;
signal \ADV_B_c_4\ : std_logic;
signal \VGA_Y_0\ : std_logic;
signal \ADV_B_c_0\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_4\ : std_logic;
signal \ADV_G_c_4\ : std_logic;
signal \ADV_B_c_7\ : std_logic;
signal \VGA_Y_1\ : std_logic;
signal \ADV_B_c_1\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_7\ : std_logic;
signal \ADV_G_c_7\ : std_logic;
signal \INVADV_G__i3C_net\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_1\ : std_logic;
signal \ADV_G_c_1\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_5\ : std_logic;
signal \ADV_G_c_5\ : std_logic;
signal \VGA_Y_6\ : std_logic;
signal \ADV_B_c_6\ : std_logic;
signal \VGA_Y_7\ : std_logic;
signal \ADV_R_c_7\ : std_logic;
signal \VGA_Y_2\ : std_logic;
signal \ADV_B_c_2\ : std_logic;
signal \INVADV_G__i2C_net\ : std_logic;
signal n1144 : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_99\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_2\ : std_logic;
signal \receive_module.rx_counter.n8\ : std_logic;
signal \receive_module.rx_counter.n7_adj_574\ : std_logic;
signal \receive_module.rx_counter.n2063_cascade_\ : std_logic;
signal \receive_module.rx_counter.n4\ : std_logic;
signal \receive_module.rx_counter.n2007\ : std_logic;
signal \receive_module.rx_counter.n2007_cascade_\ : std_logic;
signal \receive_module.rx_counter.n2069_cascade_\ : std_logic;
signal \receive_module.rx_counter.n2153\ : std_logic;
signal \receive_module.rx_counter.n2071\ : std_logic;
signal n2148 : std_logic;
signal \transmit_module.n199\ : std_logic;
signal \transmit_module.n203\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_6\ : std_logic;
signal \transmit_module.n198\ : std_logic;
signal \transmit_module.BRAM_ADDR_6\ : std_logic;
signal \transmit_module.n201\ : std_logic;
signal \transmit_module.BRAM_ADDR_1\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_1\ : std_logic;
signal \transmit_module.BRAM_ADDR_10\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_10\ : std_logic;
signal \transmit_module.BRAM_ADDR_5\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_5\ : std_logic;
signal \transmit_module.BRAM_ADDR_8\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_8\ : std_logic;
signal \transmit_module.BRAM_ADDR_11\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_11\ : std_logic;
signal \transmit_module.BRAM_ADDR_0\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_0\ : std_logic;
signal \transmit_module.BRAM_ADDR_3\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_3\ : std_logic;
signal \transmit_module.BRAM_ADDR_12\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_12\ : std_logic;
signal \transmit_module.BRAM_ADDR_2\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_2\ : std_logic;
signal \transmit_module.n792\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_33\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_32\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_31\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_30\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_20\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_19\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_18\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_22\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_21\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_17\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_29\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_28\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_27\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_26\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_25\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_24\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_23\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_0\ : std_logic;
signal \TVP_HSYNC_c\ : std_logic;
signal \receive_module.rx_counter.old_HS\ : std_logic;
signal \receive_module.rx_counter.Y_0\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \receive_module.rx_counter.Y_1\ : std_logic;
signal \receive_module.rx_counter.n1836\ : std_logic;
signal \receive_module.rx_counter.Y_2\ : std_logic;
signal \receive_module.rx_counter.n1837\ : std_logic;
signal \receive_module.rx_counter.Y_3\ : std_logic;
signal \receive_module.rx_counter.n1838\ : std_logic;
signal \receive_module.rx_counter.Y_4\ : std_logic;
signal \receive_module.rx_counter.n1839\ : std_logic;
signal \receive_module.rx_counter.Y_5\ : std_logic;
signal \receive_module.rx_counter.n1840\ : std_logic;
signal \receive_module.rx_counter.Y_6\ : std_logic;
signal \receive_module.rx_counter.n1841\ : std_logic;
signal \receive_module.rx_counter.Y_7\ : std_logic;
signal \receive_module.rx_counter.n1842\ : std_logic;
signal \receive_module.rx_counter.n1843\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \receive_module.rx_counter.Y_8\ : std_logic;
signal \receive_module.rx_counter.n752\ : std_logic;
signal \receive_module.n2155\ : std_logic;
signal \transmit_module.n197\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_7\ : std_logic;
signal \transmit_module.BRAM_ADDR_7\ : std_logic;
signal \transmit_module.n2156\ : std_logic;
signal \transmit_module.n191\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_13\ : std_logic;
signal \transmit_module.n1997\ : std_logic;
signal \transmit_module.BRAM_ADDR_13_N_257_13\ : std_logic;
signal \transmit_module.n704\ : std_logic;
signal \DEBUG_c_1\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.n694\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_16\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_8\ : std_logic;
signal \ADV_CLK_c\ : std_logic;
signal \transmit_module.n2158\ : std_logic;
signal \ADV_VSYNC_c\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \receive_module.rx_counter.n1865\ : std_logic;
signal \receive_module.rx_counter.n1866\ : std_logic;
signal \receive_module.rx_counter.n1867\ : std_logic;
signal \receive_module.rx_counter.n1868\ : std_logic;
signal \receive_module.rx_counter.n1869\ : std_logic;
signal \LED_c\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_4\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_2\ : std_logic;
signal \receive_module.rx_counter.n2150\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_5\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_1\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_0\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_3\ : std_logic;
signal \receive_module.rx_counter.n2113_cascade_\ : std_logic;
signal \receive_module.rx_counter.n7\ : std_logic;
signal \receive_module.rx_counter.n11\ : std_logic;
signal \receive_module.rx_counter.n11_cascade_\ : std_logic;
signal \receive_module.rx_counter.n1328\ : std_logic;
signal \TVP_VSYNC_c\ : std_logic;
signal \receive_module.rx_counter.old_VS\ : std_logic;
signal \TVP_CLK_c\ : std_logic;
signal \GB_BUFFER_TVP_CLK_c_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \TVP_CLK_wire\ : std_logic;
signal \ADV_CLK_wire\ : std_logic;
signal \ADV_G_wire\ : std_logic_vector(7 downto 0);
signal \ADV_B_wire\ : std_logic_vector(7 downto 0);
signal \ADV_R_wire\ : std_logic_vector(7 downto 0);
signal \ADV_VSYNC_wire\ : std_logic;
signal \ADV_SYNC_N_wire\ : std_logic;
signal \TVP_HSYNC_wire\ : std_logic;
signal \TVP_VSYNC_wire\ : std_logic;
signal \ADV_BLANK_N_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \ADV_HSYNC_wire\ : std_logic;
signal \pll2.PLL_100_TO_48MHz96_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pll1.PLL_20_TO_100MHz_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \TVP_CLK_wire\ <= TVP_CLK;
    ADV_CLK <= \ADV_CLK_wire\;
    ADV_G <= \ADV_G_wire\;
    ADV_B <= \ADV_B_wire\;
    ADV_R <= \ADV_R_wire\;
    ADV_VSYNC <= \ADV_VSYNC_wire\;
    ADV_SYNC_N <= \ADV_SYNC_N_wire\;
    \TVP_HSYNC_wire\ <= TVP_HSYNC;
    \TVP_VSYNC_wire\ <= TVP_VSYNC;
    ADV_BLANK_N <= \ADV_BLANK_N_wire\;
    LED <= \LED_wire\;
    ADV_HSYNC <= \ADV_HSYNC_wire\;
    \pll2.PLL_100_TO_48MHz96_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pll1.PLL_20_TO_100MHz_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';

    \pll2.PLL_100_TO_48MHz96_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0101",
            DIVQ => "100",
            DIVF => "0101110",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \ADV_CLK_c\,
            REFERENCECLK => \N__4486\,
            RESETB => \N__9807\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll2.PLL_100_TO_48MHz96_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \pll1.PLL_20_TO_100MHz_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0100111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \CLK_100MHz\,
            REFERENCECLK => \N__9823\,
            RESETB => \N__9811\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll1.PLL_20_TO_100MHz_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \TVP_CLK_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__10322\,
            GLOBALBUFFEROUTPUT => \TVP_CLK_c\
        );

    \TVP_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10324\,
            DIN => \N__10323\,
            DOUT => \N__10322\,
            PACKAGEPIN => \TVP_CLK_wire\
        );

    \TVP_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10324\,
            PADOUT => \N__10323\,
            PADIN => \N__10322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10313\,
            DIN => \N__10312\,
            DOUT => \N__10311\,
            PACKAGEPIN => \ADV_CLK_wire\
        );

    \ADV_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10313\,
            PADOUT => \N__10312\,
            PADIN => \N__10311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10304\,
            DIN => \N__10303\,
            DOUT => \N__10302\,
            PACKAGEPIN => DEBUG(3)
        );

    \DEBUG_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10304\,
            PADOUT => \N__10303\,
            PADIN => \N__10302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6241\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10295\,
            DIN => \N__10294\,
            DOUT => \N__10293\,
            PACKAGEPIN => \ADV_G_wire\(5)
        );

    \ADV_G_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10295\,
            PADOUT => \N__10294\,
            PADIN => \N__10293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7129\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10286\,
            DIN => \N__10285\,
            DOUT => \N__10284\,
            PACKAGEPIN => \ADV_B_wire\(3)
        );

    \ADV_B_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10286\,
            PADOUT => \N__10285\,
            PADIN => \N__10284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5671\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10277\,
            DIN => \N__10276\,
            DOUT => \N__10275\,
            PACKAGEPIN => \ADV_R_wire\(4)
        );

    \ADV_R_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10277\,
            PADOUT => \N__10276\,
            PADIN => \N__10275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5611\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10268\,
            DIN => \N__10267\,
            DOUT => \N__10266\,
            PACKAGEPIN => \ADV_B_wire\(0)
        );

    \ADV_B_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10268\,
            PADOUT => \N__10267\,
            PADIN => \N__10266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6568\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10259\,
            DIN => \N__10258\,
            DOUT => \N__10257\,
            PACKAGEPIN => \ADV_G_wire\(2)
        );

    \ADV_G_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10259\,
            PADOUT => \N__10258\,
            PADIN => \N__10257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6688\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10250\,
            DIN => \N__10249\,
            DOUT => \N__10248\,
            PACKAGEPIN => \ADV_VSYNC_wire\
        );

    \ADV_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10250\,
            PADOUT => \N__10249\,
            PADIN => \N__10248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8923\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10241\,
            DIN => \N__10240\,
            DOUT => \N__10239\,
            PACKAGEPIN => \ADV_R_wire\(3)
        );

    \ADV_R_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10241\,
            PADOUT => \N__10240\,
            PADIN => \N__10239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5404\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10232\,
            DIN => \N__10231\,
            DOUT => \N__10230\,
            PACKAGEPIN => \ADV_B_wire\(5)
        );

    \ADV_B_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10232\,
            PADOUT => \N__10231\,
            PADIN => \N__10230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5647\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10223\,
            DIN => \N__10222\,
            DOUT => \N__10221\,
            PACKAGEPIN => DEBUG(7)
        );

    \DEBUG_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10223\,
            PADOUT => \N__10222\,
            PADIN => \N__10221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10214\,
            DIN => \N__10213\,
            DOUT => \N__10212\,
            PACKAGEPIN => \ADV_G_wire\(1)
        );

    \ADV_G_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10214\,
            PADOUT => \N__10213\,
            PADIN => \N__10212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7186\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10205\,
            DIN => \N__10204\,
            DOUT => \N__10203\,
            PACKAGEPIN => \ADV_R_wire\(0)
        );

    \ADV_R_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10205\,
            PADOUT => \N__10204\,
            PADIN => \N__10203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4627\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10196\,
            DIN => \N__10195\,
            DOUT => \N__10194\,
            PACKAGEPIN => DEBUG(2)
        );

    \DEBUG_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10196\,
            PADOUT => \N__10195\,
            PADIN => \N__10194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5242\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10187\,
            DIN => \N__10186\,
            DOUT => \N__10185\,
            PACKAGEPIN => \ADV_G_wire\(4)
        );

    \ADV_G_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10187\,
            PADOUT => \N__10186\,
            PADIN => \N__10185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6526\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10178\,
            DIN => \N__10177\,
            DOUT => \N__10176\,
            PACKAGEPIN => \ADV_R_wire\(5)
        );

    \ADV_R_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10178\,
            PADOUT => \N__10177\,
            PADIN => \N__10176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5419\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10169\,
            DIN => \N__10168\,
            DOUT => \N__10167\,
            PACKAGEPIN => DEBUG(1)
        );

    \DEBUG_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10169\,
            PADOUT => \N__10168\,
            PADIN => \N__10167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10160\,
            DIN => \N__10159\,
            DOUT => \N__10158\,
            PACKAGEPIN => \ADV_B_wire\(1)
        );

    \ADV_B_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10160\,
            PADOUT => \N__10159\,
            PADIN => \N__10158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6448\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_SYNC_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10151\,
            DIN => \N__10150\,
            DOUT => \N__10149\,
            PACKAGEPIN => \ADV_SYNC_N_wire\
        );

    \ADV_SYNC_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10151\,
            PADOUT => \N__10150\,
            PADIN => \N__10149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10142\,
            DIN => \N__10141\,
            DOUT => \N__10140\,
            PACKAGEPIN => \ADV_B_wire\(6)
        );

    \ADV_B_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10142\,
            PADOUT => \N__10141\,
            PADIN => \N__10140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7060\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10133\,
            DIN => \N__10132\,
            DOUT => \N__10131\,
            PACKAGEPIN => \ADV_G_wire\(0)
        );

    \ADV_G_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10133\,
            PADOUT => \N__10132\,
            PADIN => \N__10131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5629\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10124\,
            DIN => \N__10123\,
            DOUT => \N__10122\,
            PACKAGEPIN => \ADV_R_wire\(1)
        );

    \ADV_R_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10124\,
            PADOUT => \N__10123\,
            PADIN => \N__10122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5059\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10115\,
            DIN => \N__10114\,
            DOUT => \N__10113\,
            PACKAGEPIN => DEBUG(5)
        );

    \DEBUG_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10115\,
            PADOUT => \N__10114\,
            PADIN => \N__10113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5932\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10106\,
            DIN => \N__10105\,
            DOUT => \N__10104\,
            PACKAGEPIN => \TVP_HSYNC_wire\
        );

    \TVP_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10106\,
            PADOUT => \N__10105\,
            PADIN => \N__10104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_HSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10097\,
            DIN => \N__10096\,
            DOUT => \N__10095\,
            PACKAGEPIN => \ADV_G_wire\(7)
        );

    \ADV_G_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10097\,
            PADOUT => \N__10096\,
            PADIN => \N__10095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10088\,
            DIN => \N__10087\,
            DOUT => \N__10086\,
            PACKAGEPIN => \ADV_R_wire\(6)
        );

    \ADV_R_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10088\,
            PADOUT => \N__10087\,
            PADIN => \N__10086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4612\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10079\,
            DIN => \N__10078\,
            DOUT => \N__10077\,
            PACKAGEPIN => \TVP_VSYNC_wire\
        );

    \TVP_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10079\,
            PADOUT => \N__10078\,
            PADIN => \N__10077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_BLANK_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10070\,
            DIN => \N__10069\,
            DOUT => \N__10068\,
            PACKAGEPIN => \ADV_BLANK_N_wire\
        );

    \ADV_BLANK_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10070\,
            PADOUT => \N__10069\,
            PADIN => \N__10068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9806\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__10061\,
            DIN => \N__10060\,
            DOUT => \N__10059\,
            PACKAGEPIN => DEBUG(0)
        );

    \DEBUG_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10061\,
            PADOUT => \N__10060\,
            PADIN => \N__10059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10052\,
            DIN => \N__10051\,
            DOUT => \N__10050\,
            PACKAGEPIN => \ADV_B_wire\(2)
        );

    \ADV_B_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10052\,
            PADOUT => \N__10051\,
            PADIN => \N__10050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6928\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10043\,
            DIN => \N__10042\,
            DOUT => \N__10041\,
            PACKAGEPIN => \ADV_B_wire\(7)
        );

    \ADV_B_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10043\,
            PADOUT => \N__10042\,
            PADIN => \N__10041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6514\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10034\,
            DIN => \N__10033\,
            DOUT => \N__10032\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10034\,
            PADOUT => \N__10033\,
            PADIN => \N__10032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9754\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10025\,
            DIN => \N__10024\,
            DOUT => \N__10023\,
            PACKAGEPIN => \ADV_G_wire\(3)
        );

    \ADV_G_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10025\,
            PADOUT => \N__10024\,
            PADIN => \N__10023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5722\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10016\,
            DIN => \N__10015\,
            DOUT => \N__10014\,
            PACKAGEPIN => \ADV_HSYNC_wire\
        );

    \ADV_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10016\,
            PADOUT => \N__10015\,
            PADIN => \N__10014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6196\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10007\,
            DIN => \N__10006\,
            DOUT => \N__10005\,
            PACKAGEPIN => \ADV_R_wire\(2)
        );

    \ADV_R_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__10007\,
            PADOUT => \N__10006\,
            PADIN => \N__10005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4639\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9998\,
            DIN => \N__9997\,
            DOUT => \N__9996\,
            PACKAGEPIN => \ADV_B_wire\(4)
        );

    \ADV_B_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9998\,
            PADOUT => \N__9997\,
            PADIN => \N__9996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6628\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__9989\,
            DIN => \N__9988\,
            DOUT => \N__9987\,
            PACKAGEPIN => DEBUG(4)
        );

    \DEBUG_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9989\,
            PADOUT => \N__9988\,
            PADIN => \N__9987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5899\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9980\,
            DIN => \N__9979\,
            DOUT => \N__9978\,
            PACKAGEPIN => \ADV_G_wire\(6)
        );

    \ADV_G_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9980\,
            PADOUT => \N__9979\,
            PADIN => \N__9978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5080\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9971\,
            DIN => \N__9970\,
            DOUT => \N__9969\,
            PACKAGEPIN => \ADV_R_wire\(7)
        );

    \ADV_R_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__9971\,
            PADOUT => \N__9970\,
            PADIN => \N__9969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__9952\,
            I => \receive_module.rx_counter.n11_cascade_\
        );

    \I__2211\ : SRMux
    port map (
            O => \N__9949\,
            I => \N__9946\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9946\,
            I => \N__9943\
        );

    \I__2209\ : Odrv12
    port map (
            O => \N__9943\,
            I => \receive_module.rx_counter.n1328\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9936\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9933\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9936\,
            I => \N__9925\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9933\,
            I => \N__9925\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9919\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9931\,
            I => \N__9919\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9930\,
            I => \N__9916\
        );

    \I__2201\ : Span4Mux_v
    port map (
            O => \N__9925\,
            I => \N__9913\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9910\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9919\,
            I => \N__9907\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9916\,
            I => \N__9904\
        );

    \I__2197\ : Sp12to4
    port map (
            O => \N__9913\,
            I => \N__9899\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9910\,
            I => \N__9899\
        );

    \I__2195\ : Span4Mux_v
    port map (
            O => \N__9907\,
            I => \N__9896\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__9904\,
            I => \N__9893\
        );

    \I__2193\ : Span12Mux_h
    port map (
            O => \N__9899\,
            I => \N__9890\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__9896\,
            I => \N__9885\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__9893\,
            I => \N__9885\
        );

    \I__2190\ : Odrv12
    port map (
            O => \N__9890\,
            I => \TVP_VSYNC_c\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__9885\,
            I => \TVP_VSYNC_c\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9874\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9879\,
            I => \N__9874\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9874\,
            I => \receive_module.rx_counter.old_VS\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9868\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9868\,
            I => \N__9854\
        );

    \I__2183\ : ClkMux
    port map (
            O => \N__9867\,
            I => \N__9829\
        );

    \I__2182\ : ClkMux
    port map (
            O => \N__9866\,
            I => \N__9829\
        );

    \I__2181\ : ClkMux
    port map (
            O => \N__9865\,
            I => \N__9829\
        );

    \I__2180\ : ClkMux
    port map (
            O => \N__9864\,
            I => \N__9829\
        );

    \I__2179\ : ClkMux
    port map (
            O => \N__9863\,
            I => \N__9829\
        );

    \I__2178\ : ClkMux
    port map (
            O => \N__9862\,
            I => \N__9829\
        );

    \I__2177\ : ClkMux
    port map (
            O => \N__9861\,
            I => \N__9829\
        );

    \I__2176\ : ClkMux
    port map (
            O => \N__9860\,
            I => \N__9829\
        );

    \I__2175\ : ClkMux
    port map (
            O => \N__9859\,
            I => \N__9829\
        );

    \I__2174\ : ClkMux
    port map (
            O => \N__9858\,
            I => \N__9829\
        );

    \I__2173\ : ClkMux
    port map (
            O => \N__9857\,
            I => \N__9829\
        );

    \I__2172\ : Glb2LocalMux
    port map (
            O => \N__9854\,
            I => \N__9829\
        );

    \I__2171\ : GlobalMux
    port map (
            O => \N__9829\,
            I => \N__9826\
        );

    \I__2170\ : gio2CtrlBuf
    port map (
            O => \N__9826\,
            I => \TVP_CLK_c\
        );

    \I__2169\ : IoInMux
    port map (
            O => \N__9823\,
            I => \N__9820\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9820\,
            I => \N__9817\
        );

    \I__2167\ : Span4Mux_s0_v
    port map (
            O => \N__9817\,
            I => \N__9814\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__9814\,
            I => \GB_BUFFER_TVP_CLK_c_THRU_CO\
        );

    \I__2165\ : IoInMux
    port map (
            O => \N__9811\,
            I => \N__9808\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9808\,
            I => \N__9803\
        );

    \I__2163\ : IoInMux
    port map (
            O => \N__9807\,
            I => \N__9800\
        );

    \I__2162\ : IoInMux
    port map (
            O => \N__9806\,
            I => \N__9797\
        );

    \I__2161\ : IoSpan4Mux
    port map (
            O => \N__9803\,
            I => \N__9794\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9800\,
            I => \N__9789\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9789\
        );

    \I__2158\ : Span4Mux_s2_v
    port map (
            O => \N__9794\,
            I => \N__9786\
        );

    \I__2157\ : Span4Mux_s1_v
    port map (
            O => \N__9789\,
            I => \N__9783\
        );

    \I__2156\ : Sp12to4
    port map (
            O => \N__9786\,
            I => \N__9780\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__9783\,
            I => \N__9777\
        );

    \I__2154\ : Span12Mux_v
    port map (
            O => \N__9780\,
            I => \N__9774\
        );

    \I__2153\ : Span4Mux_v
    port map (
            O => \N__9777\,
            I => \N__9771\
        );

    \I__2152\ : Odrv12
    port map (
            O => \N__9774\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__9771\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9766\,
            I => \receive_module.rx_counter.n1866\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9763\,
            I => \receive_module.rx_counter.n1867\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9760\,
            I => \receive_module.rx_counter.n1868\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9757\,
            I => \receive_module.rx_counter.n1869\
        );

    \I__2146\ : IoInMux
    port map (
            O => \N__9754\,
            I => \N__9751\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9748\
        );

    \I__2144\ : Span12Mux_s1_v
    port map (
            O => \N__9748\,
            I => \N__9745\
        );

    \I__2143\ : Span12Mux_h
    port map (
            O => \N__9745\,
            I => \N__9741\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9744\,
            I => \N__9738\
        );

    \I__2141\ : Odrv12
    port map (
            O => \N__9741\,
            I => \LED_c\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9738\,
            I => \LED_c\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9729\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9726\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9729\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9726\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__2135\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9717\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9714\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9717\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9714\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__2131\ : CEMux
    port map (
            O => \N__9709\,
            I => \N__9705\
        );

    \I__2130\ : CEMux
    port map (
            O => \N__9708\,
            I => \N__9702\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9705\,
            I => \receive_module.rx_counter.n2150\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9702\,
            I => \receive_module.rx_counter.n2150\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9693\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9690\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9693\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9690\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9685\,
            I => \N__9681\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9684\,
            I => \N__9678\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9681\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9678\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9669\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9666\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9669\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9666\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__2115\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9657\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9654\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9657\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9654\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__9649\,
            I => \receive_module.rx_counter.n2113_cascade_\
        );

    \I__2110\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9643\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9643\,
            I => \receive_module.rx_counter.n7\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9637\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9637\,
            I => \receive_module.rx_counter.n11\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9631\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9631\,
            I => \transmit_module.Y_DELTA_PATTERN_14\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9625\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9625\,
            I => \transmit_module.Y_DELTA_PATTERN_13\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9619\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9619\,
            I => \transmit_module.Y_DELTA_PATTERN_12\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9613\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9613\,
            I => \transmit_module.Y_DELTA_PATTERN_11\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9607\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9607\,
            I => \transmit_module.Y_DELTA_PATTERN_10\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9601\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9601\,
            I => \transmit_module.Y_DELTA_PATTERN_7\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9598\,
            I => \N__9595\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9595\,
            I => \transmit_module.Y_DELTA_PATTERN_9\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9589\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9589\,
            I => \transmit_module.Y_DELTA_PATTERN_8\
        );

    \I__2090\ : ClkMux
    port map (
            O => \N__9586\,
            I => \N__9581\
        );

    \I__2089\ : ClkMux
    port map (
            O => \N__9585\,
            I => \N__9578\
        );

    \I__2088\ : ClkMux
    port map (
            O => \N__9584\,
            I => \N__9572\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__9581\,
            I => \N__9560\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9578\,
            I => \N__9560\
        );

    \I__2085\ : ClkMux
    port map (
            O => \N__9577\,
            I => \N__9557\
        );

    \I__2084\ : ClkMux
    port map (
            O => \N__9576\,
            I => \N__9554\
        );

    \I__2083\ : ClkMux
    port map (
            O => \N__9575\,
            I => \N__9551\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9545\
        );

    \I__2081\ : ClkMux
    port map (
            O => \N__9571\,
            I => \N__9542\
        );

    \I__2080\ : ClkMux
    port map (
            O => \N__9570\,
            I => \N__9536\
        );

    \I__2079\ : ClkMux
    port map (
            O => \N__9569\,
            I => \N__9533\
        );

    \I__2078\ : ClkMux
    port map (
            O => \N__9568\,
            I => \N__9528\
        );

    \I__2077\ : ClkMux
    port map (
            O => \N__9567\,
            I => \N__9525\
        );

    \I__2076\ : ClkMux
    port map (
            O => \N__9566\,
            I => \N__9522\
        );

    \I__2075\ : ClkMux
    port map (
            O => \N__9565\,
            I => \N__9516\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__9560\,
            I => \N__9509\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9557\,
            I => \N__9509\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__9554\,
            I => \N__9509\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9551\,
            I => \N__9506\
        );

    \I__2070\ : ClkMux
    port map (
            O => \N__9550\,
            I => \N__9503\
        );

    \I__2069\ : ClkMux
    port map (
            O => \N__9549\,
            I => \N__9500\
        );

    \I__2068\ : ClkMux
    port map (
            O => \N__9548\,
            I => \N__9497\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__9545\,
            I => \N__9490\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9542\,
            I => \N__9490\
        );

    \I__2065\ : ClkMux
    port map (
            O => \N__9541\,
            I => \N__9487\
        );

    \I__2064\ : ClkMux
    port map (
            O => \N__9540\,
            I => \N__9484\
        );

    \I__2063\ : ClkMux
    port map (
            O => \N__9539\,
            I => \N__9481\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9536\,
            I => \N__9478\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9533\,
            I => \N__9475\
        );

    \I__2060\ : ClkMux
    port map (
            O => \N__9532\,
            I => \N__9472\
        );

    \I__2059\ : ClkMux
    port map (
            O => \N__9531\,
            I => \N__9468\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9528\,
            I => \N__9463\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__9525\,
            I => \N__9463\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9522\,
            I => \N__9457\
        );

    \I__2055\ : ClkMux
    port map (
            O => \N__9521\,
            I => \N__9454\
        );

    \I__2054\ : ClkMux
    port map (
            O => \N__9520\,
            I => \N__9451\
        );

    \I__2053\ : ClkMux
    port map (
            O => \N__9519\,
            I => \N__9443\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9516\,
            I => \N__9439\
        );

    \I__2051\ : Span4Mux_v
    port map (
            O => \N__9509\,
            I => \N__9436\
        );

    \I__2050\ : Span4Mux_h
    port map (
            O => \N__9506\,
            I => \N__9427\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9503\,
            I => \N__9427\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9427\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9497\,
            I => \N__9427\
        );

    \I__2046\ : ClkMux
    port map (
            O => \N__9496\,
            I => \N__9424\
        );

    \I__2045\ : ClkMux
    port map (
            O => \N__9495\,
            I => \N__9419\
        );

    \I__2044\ : Span4Mux_h
    port map (
            O => \N__9490\,
            I => \N__9414\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9487\,
            I => \N__9414\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9484\,
            I => \N__9409\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9481\,
            I => \N__9409\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__9478\,
            I => \N__9402\
        );

    \I__2039\ : Span4Mux_h
    port map (
            O => \N__9475\,
            I => \N__9402\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9472\,
            I => \N__9402\
        );

    \I__2037\ : ClkMux
    port map (
            O => \N__9471\,
            I => \N__9399\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9468\,
            I => \N__9395\
        );

    \I__2035\ : Span4Mux_v
    port map (
            O => \N__9463\,
            I => \N__9392\
        );

    \I__2034\ : ClkMux
    port map (
            O => \N__9462\,
            I => \N__9389\
        );

    \I__2033\ : ClkMux
    port map (
            O => \N__9461\,
            I => \N__9386\
        );

    \I__2032\ : ClkMux
    port map (
            O => \N__9460\,
            I => \N__9380\
        );

    \I__2031\ : Span4Mux_v
    port map (
            O => \N__9457\,
            I => \N__9373\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9454\,
            I => \N__9373\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9451\,
            I => \N__9373\
        );

    \I__2028\ : ClkMux
    port map (
            O => \N__9450\,
            I => \N__9370\
        );

    \I__2027\ : ClkMux
    port map (
            O => \N__9449\,
            I => \N__9367\
        );

    \I__2026\ : ClkMux
    port map (
            O => \N__9448\,
            I => \N__9364\
        );

    \I__2025\ : ClkMux
    port map (
            O => \N__9447\,
            I => \N__9361\
        );

    \I__2024\ : ClkMux
    port map (
            O => \N__9446\,
            I => \N__9357\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9443\,
            I => \N__9351\
        );

    \I__2022\ : ClkMux
    port map (
            O => \N__9442\,
            I => \N__9348\
        );

    \I__2021\ : Span4Mux_h
    port map (
            O => \N__9439\,
            I => \N__9339\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__9436\,
            I => \N__9339\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__9427\,
            I => \N__9339\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9424\,
            I => \N__9339\
        );

    \I__2017\ : ClkMux
    port map (
            O => \N__9423\,
            I => \N__9336\
        );

    \I__2016\ : ClkMux
    port map (
            O => \N__9422\,
            I => \N__9333\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9419\,
            I => \N__9329\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__9414\,
            I => \N__9320\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__9409\,
            I => \N__9320\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__9402\,
            I => \N__9320\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9399\,
            I => \N__9320\
        );

    \I__2010\ : ClkMux
    port map (
            O => \N__9398\,
            I => \N__9317\
        );

    \I__2009\ : Span4Mux_v
    port map (
            O => \N__9395\,
            I => \N__9308\
        );

    \I__2008\ : Span4Mux_h
    port map (
            O => \N__9392\,
            I => \N__9308\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__9389\,
            I => \N__9308\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9386\,
            I => \N__9308\
        );

    \I__2005\ : ClkMux
    port map (
            O => \N__9385\,
            I => \N__9305\
        );

    \I__2004\ : ClkMux
    port map (
            O => \N__9384\,
            I => \N__9302\
        );

    \I__2003\ : ClkMux
    port map (
            O => \N__9383\,
            I => \N__9299\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9380\,
            I => \N__9296\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__9373\,
            I => \N__9289\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9370\,
            I => \N__9289\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__9367\,
            I => \N__9289\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9364\,
            I => \N__9284\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9361\,
            I => \N__9284\
        );

    \I__1996\ : ClkMux
    port map (
            O => \N__9360\,
            I => \N__9281\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__9357\,
            I => \N__9277\
        );

    \I__1994\ : ClkMux
    port map (
            O => \N__9356\,
            I => \N__9274\
        );

    \I__1993\ : ClkMux
    port map (
            O => \N__9355\,
            I => \N__9271\
        );

    \I__1992\ : ClkMux
    port map (
            O => \N__9354\,
            I => \N__9268\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__9351\,
            I => \N__9264\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9348\,
            I => \N__9255\
        );

    \I__1989\ : Span4Mux_h
    port map (
            O => \N__9339\,
            I => \N__9255\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9336\,
            I => \N__9255\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__9333\,
            I => \N__9255\
        );

    \I__1986\ : ClkMux
    port map (
            O => \N__9332\,
            I => \N__9252\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__9329\,
            I => \N__9249\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__9320\,
            I => \N__9244\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__9317\,
            I => \N__9244\
        );

    \I__1982\ : Span4Mux_v
    port map (
            O => \N__9308\,
            I => \N__9235\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9305\,
            I => \N__9235\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9302\,
            I => \N__9235\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9299\,
            I => \N__9235\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__9296\,
            I => \N__9226\
        );

    \I__1977\ : Span4Mux_h
    port map (
            O => \N__9289\,
            I => \N__9226\
        );

    \I__1976\ : Span4Mux_h
    port map (
            O => \N__9284\,
            I => \N__9226\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__9281\,
            I => \N__9226\
        );

    \I__1974\ : ClkMux
    port map (
            O => \N__9280\,
            I => \N__9223\
        );

    \I__1973\ : Span4Mux_v
    port map (
            O => \N__9277\,
            I => \N__9216\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__9274\,
            I => \N__9216\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9271\,
            I => \N__9211\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__9268\,
            I => \N__9211\
        );

    \I__1969\ : ClkMux
    port map (
            O => \N__9267\,
            I => \N__9208\
        );

    \I__1968\ : Span4Mux_h
    port map (
            O => \N__9264\,
            I => \N__9201\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__9255\,
            I => \N__9201\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9201\
        );

    \I__1965\ : Span4Mux_h
    port map (
            O => \N__9249\,
            I => \N__9190\
        );

    \I__1964\ : Span4Mux_v
    port map (
            O => \N__9244\,
            I => \N__9190\
        );

    \I__1963\ : Span4Mux_v
    port map (
            O => \N__9235\,
            I => \N__9190\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__9226\,
            I => \N__9190\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9223\,
            I => \N__9190\
        );

    \I__1960\ : IoInMux
    port map (
            O => \N__9222\,
            I => \N__9187\
        );

    \I__1959\ : ClkMux
    port map (
            O => \N__9221\,
            I => \N__9184\
        );

    \I__1958\ : Span4Mux_v
    port map (
            O => \N__9216\,
            I => \N__9177\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__9211\,
            I => \N__9177\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__9208\,
            I => \N__9177\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__9201\,
            I => \N__9174\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__9190\,
            I => \N__9171\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__9187\,
            I => \N__9168\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__9184\,
            I => \N__9165\
        );

    \I__1951\ : Sp12to4
    port map (
            O => \N__9177\,
            I => \N__9162\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__9174\,
            I => \N__9159\
        );

    \I__1949\ : Span4Mux_v
    port map (
            O => \N__9171\,
            I => \N__9156\
        );

    \I__1948\ : IoSpan4Mux
    port map (
            O => \N__9168\,
            I => \N__9153\
        );

    \I__1947\ : Span12Mux_h
    port map (
            O => \N__9165\,
            I => \N__9150\
        );

    \I__1946\ : Span12Mux_v
    port map (
            O => \N__9162\,
            I => \N__9147\
        );

    \I__1945\ : Sp12to4
    port map (
            O => \N__9159\,
            I => \N__9142\
        );

    \I__1944\ : Sp12to4
    port map (
            O => \N__9156\,
            I => \N__9142\
        );

    \I__1943\ : IoSpan4Mux
    port map (
            O => \N__9153\,
            I => \N__9139\
        );

    \I__1942\ : Span12Mux_v
    port map (
            O => \N__9150\,
            I => \N__9134\
        );

    \I__1941\ : Span12Mux_h
    port map (
            O => \N__9147\,
            I => \N__9134\
        );

    \I__1940\ : Span12Mux_h
    port map (
            O => \N__9142\,
            I => \N__9131\
        );

    \I__1939\ : IoSpan4Mux
    port map (
            O => \N__9139\,
            I => \N__9128\
        );

    \I__1938\ : Odrv12
    port map (
            O => \N__9134\,
            I => \ADV_CLK_c\
        );

    \I__1937\ : Odrv12
    port map (
            O => \N__9131\,
            I => \ADV_CLK_c\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__9128\,
            I => \ADV_CLK_c\
        );

    \I__1935\ : CEMux
    port map (
            O => \N__9121\,
            I => \N__9118\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__9118\,
            I => \N__9111\
        );

    \I__1933\ : CEMux
    port map (
            O => \N__9117\,
            I => \N__9106\
        );

    \I__1932\ : CEMux
    port map (
            O => \N__9116\,
            I => \N__9103\
        );

    \I__1931\ : CEMux
    port map (
            O => \N__9115\,
            I => \N__9100\
        );

    \I__1930\ : CEMux
    port map (
            O => \N__9114\,
            I => \N__9096\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__9111\,
            I => \N__9093\
        );

    \I__1928\ : CEMux
    port map (
            O => \N__9110\,
            I => \N__9090\
        );

    \I__1927\ : CEMux
    port map (
            O => \N__9109\,
            I => \N__9087\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__9106\,
            I => \N__9077\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9103\,
            I => \N__9077\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9100\,
            I => \N__9077\
        );

    \I__1923\ : CEMux
    port map (
            O => \N__9099\,
            I => \N__9074\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9096\,
            I => \N__9071\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__9093\,
            I => \N__9063\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__9090\,
            I => \N__9063\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9063\
        );

    \I__1918\ : SRMux
    port map (
            O => \N__9086\,
            I => \N__9060\
        );

    \I__1917\ : SRMux
    port map (
            O => \N__9085\,
            I => \N__9057\
        );

    \I__1916\ : CEMux
    port map (
            O => \N__9084\,
            I => \N__9054\
        );

    \I__1915\ : Span4Mux_v
    port map (
            O => \N__9077\,
            I => \N__9049\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__9074\,
            I => \N__9049\
        );

    \I__1913\ : Span4Mux_h
    port map (
            O => \N__9071\,
            I => \N__9045\
        );

    \I__1912\ : CEMux
    port map (
            O => \N__9070\,
            I => \N__9042\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__9063\,
            I => \N__9037\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9037\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9034\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__9054\,
            I => \N__9031\
        );

    \I__1907\ : Span4Mux_v
    port map (
            O => \N__9049\,
            I => \N__9028\
        );

    \I__1906\ : SRMux
    port map (
            O => \N__9048\,
            I => \N__9025\
        );

    \I__1905\ : Sp12to4
    port map (
            O => \N__9045\,
            I => \N__9020\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9042\,
            I => \N__9020\
        );

    \I__1903\ : Span4Mux_h
    port map (
            O => \N__9037\,
            I => \N__9017\
        );

    \I__1902\ : Span4Mux_h
    port map (
            O => \N__9034\,
            I => \N__9014\
        );

    \I__1901\ : Span4Mux_h
    port map (
            O => \N__9031\,
            I => \N__9007\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__9028\,
            I => \N__9007\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__9025\,
            I => \N__9007\
        );

    \I__1898\ : Odrv12
    port map (
            O => \N__9020\,
            I => \transmit_module.n2158\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__9017\,
            I => \transmit_module.n2158\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__9014\,
            I => \transmit_module.n2158\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__9007\,
            I => \transmit_module.n2158\
        );

    \I__1894\ : SRMux
    port map (
            O => \N__8998\,
            I => \N__8986\
        );

    \I__1893\ : SRMux
    port map (
            O => \N__8997\,
            I => \N__8983\
        );

    \I__1892\ : SRMux
    port map (
            O => \N__8996\,
            I => \N__8969\
        );

    \I__1891\ : SRMux
    port map (
            O => \N__8995\,
            I => \N__8965\
        );

    \I__1890\ : SRMux
    port map (
            O => \N__8994\,
            I => \N__8961\
        );

    \I__1889\ : SRMux
    port map (
            O => \N__8993\,
            I => \N__8957\
        );

    \I__1888\ : SRMux
    port map (
            O => \N__8992\,
            I => \N__8954\
        );

    \I__1887\ : SRMux
    port map (
            O => \N__8991\,
            I => \N__8951\
        );

    \I__1886\ : SRMux
    port map (
            O => \N__8990\,
            I => \N__8947\
        );

    \I__1885\ : SRMux
    port map (
            O => \N__8989\,
            I => \N__8944\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8986\,
            I => \N__8940\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8983\,
            I => \N__8937\
        );

    \I__1882\ : SRMux
    port map (
            O => \N__8982\,
            I => \N__8934\
        );

    \I__1881\ : SRMux
    port map (
            O => \N__8981\,
            I => \N__8930\
        );

    \I__1880\ : SRMux
    port map (
            O => \N__8980\,
            I => \N__8927\
        );

    \I__1879\ : SRMux
    port map (
            O => \N__8979\,
            I => \N__8920\
        );

    \I__1878\ : SRMux
    port map (
            O => \N__8978\,
            I => \N__8917\
        );

    \I__1877\ : SRMux
    port map (
            O => \N__8977\,
            I => \N__8913\
        );

    \I__1876\ : SRMux
    port map (
            O => \N__8976\,
            I => \N__8910\
        );

    \I__1875\ : SRMux
    port map (
            O => \N__8975\,
            I => \N__8905\
        );

    \I__1874\ : SRMux
    port map (
            O => \N__8974\,
            I => \N__8902\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__8973\,
            I => \N__8899\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__8972\,
            I => \N__8896\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8969\,
            I => \N__8890\
        );

    \I__1870\ : SRMux
    port map (
            O => \N__8968\,
            I => \N__8887\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8965\,
            I => \N__8884\
        );

    \I__1868\ : SRMux
    port map (
            O => \N__8964\,
            I => \N__8881\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8961\,
            I => \N__8878\
        );

    \I__1866\ : SRMux
    port map (
            O => \N__8960\,
            I => \N__8875\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8957\,
            I => \N__8872\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8954\,
            I => \N__8869\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8951\,
            I => \N__8866\
        );

    \I__1862\ : SRMux
    port map (
            O => \N__8950\,
            I => \N__8863\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8947\,
            I => \N__8860\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8944\,
            I => \N__8857\
        );

    \I__1859\ : SRMux
    port map (
            O => \N__8943\,
            I => \N__8854\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__8940\,
            I => \N__8847\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__8937\,
            I => \N__8847\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8934\,
            I => \N__8847\
        );

    \I__1855\ : SRMux
    port map (
            O => \N__8933\,
            I => \N__8844\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8930\,
            I => \N__8837\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8927\,
            I => \N__8837\
        );

    \I__1852\ : SRMux
    port map (
            O => \N__8926\,
            I => \N__8834\
        );

    \I__1851\ : SRMux
    port map (
            O => \N__8925\,
            I => \N__8831\
        );

    \I__1850\ : SRMux
    port map (
            O => \N__8924\,
            I => \N__8828\
        );

    \I__1849\ : IoInMux
    port map (
            O => \N__8923\,
            I => \N__8824\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8920\,
            I => \N__8821\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8917\,
            I => \N__8818\
        );

    \I__1846\ : SRMux
    port map (
            O => \N__8916\,
            I => \N__8815\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8913\,
            I => \N__8810\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8810\
        );

    \I__1843\ : SRMux
    port map (
            O => \N__8909\,
            I => \N__8807\
        );

    \I__1842\ : SRMux
    port map (
            O => \N__8908\,
            I => \N__8804\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8905\,
            I => \N__8801\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8902\,
            I => \N__8798\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8793\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8793\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8786\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8786\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8786\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__8890\,
            I => \N__8781\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8887\,
            I => \N__8781\
        );

    \I__1832\ : Span4Mux_h
    port map (
            O => \N__8884\,
            I => \N__8778\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8881\,
            I => \N__8771\
        );

    \I__1830\ : Span4Mux_h
    port map (
            O => \N__8878\,
            I => \N__8771\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8875\,
            I => \N__8771\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__8872\,
            I => \N__8762\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__8869\,
            I => \N__8762\
        );

    \I__1826\ : Span4Mux_h
    port map (
            O => \N__8866\,
            I => \N__8762\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8863\,
            I => \N__8762\
        );

    \I__1824\ : Span4Mux_v
    port map (
            O => \N__8860\,
            I => \N__8755\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__8857\,
            I => \N__8755\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8854\,
            I => \N__8755\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__8847\,
            I => \N__8750\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8844\,
            I => \N__8750\
        );

    \I__1819\ : SRMux
    port map (
            O => \N__8843\,
            I => \N__8747\
        );

    \I__1818\ : SRMux
    port map (
            O => \N__8842\,
            I => \N__8744\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__8837\,
            I => \N__8737\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8737\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8831\,
            I => \N__8737\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8734\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__8827\,
            I => \N__8731\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8824\,
            I => \N__8728\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__8821\,
            I => \N__8721\
        );

    \I__1810\ : Span4Mux_v
    port map (
            O => \N__8818\,
            I => \N__8721\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8815\,
            I => \N__8721\
        );

    \I__1808\ : Span4Mux_h
    port map (
            O => \N__8810\,
            I => \N__8716\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8807\,
            I => \N__8716\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8804\,
            I => \N__8713\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__8801\,
            I => \N__8704\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__8798\,
            I => \N__8704\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8793\,
            I => \N__8704\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8786\,
            I => \N__8704\
        );

    \I__1801\ : Span4Mux_v
    port map (
            O => \N__8781\,
            I => \N__8697\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__8778\,
            I => \N__8697\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__8771\,
            I => \N__8697\
        );

    \I__1798\ : Span4Mux_h
    port map (
            O => \N__8762\,
            I => \N__8690\
        );

    \I__1797\ : Span4Mux_h
    port map (
            O => \N__8755\,
            I => \N__8690\
        );

    \I__1796\ : Span4Mux_s2_h
    port map (
            O => \N__8750\,
            I => \N__8690\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8687\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8684\
        );

    \I__1793\ : Span4Mux_v
    port map (
            O => \N__8737\,
            I => \N__8679\
        );

    \I__1792\ : Span4Mux_s3_h
    port map (
            O => \N__8734\,
            I => \N__8679\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8676\
        );

    \I__1790\ : Span4Mux_s2_h
    port map (
            O => \N__8728\,
            I => \N__8665\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__8721\,
            I => \N__8665\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__8716\,
            I => \N__8665\
        );

    \I__1787\ : Span4Mux_s2_h
    port map (
            O => \N__8713\,
            I => \N__8665\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__8704\,
            I => \N__8665\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__8697\,
            I => \ADV_VSYNC_c\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__8690\,
            I => \ADV_VSYNC_c\
        );

    \I__1783\ : Odrv12
    port map (
            O => \N__8687\,
            I => \ADV_VSYNC_c\
        );

    \I__1782\ : Odrv12
    port map (
            O => \N__8684\,
            I => \ADV_VSYNC_c\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__8679\,
            I => \ADV_VSYNC_c\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8676\,
            I => \ADV_VSYNC_c\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__8665\,
            I => \ADV_VSYNC_c\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8650\,
            I => \bfn_9_7_0_\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8647\,
            I => \receive_module.rx_counter.n1865\
        );

    \I__1776\ : SRMux
    port map (
            O => \N__8644\,
            I => \N__8641\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8641\,
            I => \N__8637\
        );

    \I__1774\ : SRMux
    port map (
            O => \N__8640\,
            I => \N__8632\
        );

    \I__1773\ : Span4Mux_v
    port map (
            O => \N__8637\,
            I => \N__8629\
        );

    \I__1772\ : SRMux
    port map (
            O => \N__8636\,
            I => \N__8626\
        );

    \I__1771\ : SRMux
    port map (
            O => \N__8635\,
            I => \N__8623\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8632\,
            I => \N__8620\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__8629\,
            I => \N__8615\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8626\,
            I => \N__8615\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8623\,
            I => \N__8612\
        );

    \I__1766\ : Span4Mux_h
    port map (
            O => \N__8620\,
            I => \N__8609\
        );

    \I__1765\ : Sp12to4
    port map (
            O => \N__8615\,
            I => \N__8606\
        );

    \I__1764\ : Span4Mux_h
    port map (
            O => \N__8612\,
            I => \N__8603\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__8609\,
            I => \receive_module.n2155\
        );

    \I__1762\ : Odrv12
    port map (
            O => \N__8606\,
            I => \receive_module.n2155\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__8603\,
            I => \receive_module.n2155\
        );

    \I__1760\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8593\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8593\,
            I => \N__8590\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__8590\,
            I => \N__8587\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__8587\,
            I => \transmit_module.n197\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__8584\,
            I => \N__8581\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8578\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8578\,
            I => \transmit_module.ADDR_Y_COMPONENT_7\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8572\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8572\,
            I => \N__8568\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8565\
        );

    \I__1750\ : Span4Mux_h
    port map (
            O => \N__8568\,
            I => \N__8562\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8565\,
            I => \transmit_module.BRAM_ADDR_7\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__8562\,
            I => \transmit_module.BRAM_ADDR_7\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8551\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__8556\,
            I => \N__8544\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__8555\,
            I => \N__8541\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__8554\,
            I => \N__8538\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8551\,
            I => \N__8534\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8531\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8528\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__8548\,
            I => \N__8521\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8516\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8507\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8507\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8507\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8507\
        );

    \I__1734\ : Span4Mux_h
    port map (
            O => \N__8534\,
            I => \N__8502\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8531\,
            I => \N__8502\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8528\,
            I => \N__8499\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8484\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8526\,
            I => \N__8484\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8484\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8484\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8484\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8484\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8484\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8516\,
            I => \N__8481\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8478\
        );

    \I__1722\ : Span4Mux_v
    port map (
            O => \N__8502\,
            I => \N__8473\
        );

    \I__1721\ : Span4Mux_v
    port map (
            O => \N__8499\,
            I => \N__8473\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8484\,
            I => \transmit_module.n2156\
        );

    \I__1719\ : Odrv12
    port map (
            O => \N__8481\,
            I => \transmit_module.n2156\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__8478\,
            I => \transmit_module.n2156\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__8473\,
            I => \transmit_module.n2156\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8461\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8461\,
            I => \N__8458\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__8458\,
            I => \transmit_module.n191\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__8455\,
            I => \N__8452\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8449\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8449\,
            I => \transmit_module.ADDR_Y_COMPONENT_13\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8446\,
            I => \N__8432\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8432\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8432\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8432\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8442\,
            I => \N__8428\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8418\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8415\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8412\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8428\,
            I => \N__8403\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8388\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8388\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8388\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8388\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8388\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8388\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8388\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8418\,
            I => \N__8385\
        );

    \I__1693\ : Span4Mux_h
    port map (
            O => \N__8415\,
            I => \N__8381\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8412\,
            I => \N__8378\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8371\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8410\,
            I => \N__8371\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8371\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8366\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8366\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8363\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__8403\,
            I => \N__8356\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__8388\,
            I => \N__8356\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__8385\,
            I => \N__8356\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8353\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__8381\,
            I => \N__8350\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__8378\,
            I => \N__8345\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8345\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8366\,
            I => \N__8336\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8363\,
            I => \N__8336\
        );

    \I__1676\ : Span4Mux_h
    port map (
            O => \N__8356\,
            I => \N__8336\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8353\,
            I => \N__8336\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__8350\,
            I => \transmit_module.n1997\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__8345\,
            I => \transmit_module.n1997\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__8336\,
            I => \transmit_module.n1997\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8326\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8323\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__8323\,
            I => \transmit_module.BRAM_ADDR_13_N_257_13\
        );

    \I__1668\ : CEMux
    port map (
            O => \N__8320\,
            I => \N__8317\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8317\,
            I => \N__8312\
        );

    \I__1666\ : CEMux
    port map (
            O => \N__8316\,
            I => \N__8309\
        );

    \I__1665\ : CEMux
    port map (
            O => \N__8315\,
            I => \N__8306\
        );

    \I__1664\ : Span4Mux_h
    port map (
            O => \N__8312\,
            I => \N__8299\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8309\,
            I => \N__8299\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__8306\,
            I => \N__8296\
        );

    \I__1661\ : CEMux
    port map (
            O => \N__8305\,
            I => \N__8293\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8290\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__8299\,
            I => \N__8287\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__8296\,
            I => \N__8284\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__8293\,
            I => \N__8281\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__8290\,
            I => \N__8278\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__8287\,
            I => \transmit_module.n704\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__8284\,
            I => \transmit_module.n704\
        );

    \I__1653\ : Odrv12
    port map (
            O => \N__8281\,
            I => \transmit_module.n704\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__8278\,
            I => \transmit_module.n704\
        );

    \I__1651\ : IoInMux
    port map (
            O => \N__8269\,
            I => \N__8266\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8266\,
            I => \N__8261\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8258\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8255\
        );

    \I__1647\ : Span12Mux_s6_h
    port map (
            O => \N__8261\,
            I => \N__8252\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8246\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8255\,
            I => \N__8246\
        );

    \I__1644\ : Span12Mux_v
    port map (
            O => \N__8252\,
            I => \N__8243\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8240\
        );

    \I__1642\ : Span4Mux_h
    port map (
            O => \N__8246\,
            I => \N__8237\
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__8243\,
            I => \DEBUG_c_1\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__8240\,
            I => \DEBUG_c_1\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__8237\,
            I => \DEBUG_c_1\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8227\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8227\,
            I => \transmit_module.X_DELTA_PATTERN_10\
        );

    \I__1636\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8221\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8221\,
            I => \transmit_module.X_DELTA_PATTERN_11\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__8215\,
            I => \transmit_module.X_DELTA_PATTERN_13\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__8209\,
            I => \transmit_module.X_DELTA_PATTERN_12\
        );

    \I__1630\ : CEMux
    port map (
            O => \N__8206\,
            I => \N__8202\
        );

    \I__1629\ : CEMux
    port map (
            O => \N__8205\,
            I => \N__8199\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8196\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8193\
        );

    \I__1626\ : Span4Mux_v
    port map (
            O => \N__8196\,
            I => \N__8187\
        );

    \I__1625\ : Span4Mux_h
    port map (
            O => \N__8193\,
            I => \N__8187\
        );

    \I__1624\ : CEMux
    port map (
            O => \N__8192\,
            I => \N__8184\
        );

    \I__1623\ : Sp12to4
    port map (
            O => \N__8187\,
            I => \N__8179\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__8184\,
            I => \N__8179\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__8179\,
            I => \transmit_module.n694\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8176\,
            I => \N__8173\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8173\,
            I => \transmit_module.Y_DELTA_PATTERN_16\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8170\,
            I => \N__8167\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8167\,
            I => \transmit_module.Y_DELTA_PATTERN_15\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8159\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8154\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8154\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8159\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8154\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8149\,
            I => \receive_module.rx_counter.n1836\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__8146\,
            I => \N__8140\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8145\,
            I => \N__8137\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8134\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8129\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8129\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8137\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__8134\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__8129\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8122\,
            I => \receive_module.rx_counter.n1837\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__8119\,
            I => \N__8115\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8110\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8107\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8102\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8102\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__8110\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8107\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8102\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__1593\ : InMux
    port map (
            O => \N__8095\,
            I => \receive_module.rx_counter.n1838\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8086\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8083\
        );

    \I__1590\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8078\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8078\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__8086\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__8083\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__8078\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__1585\ : InMux
    port map (
            O => \N__8071\,
            I => \receive_module.rx_counter.n1839\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8068\,
            I => \N__8063\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8067\,
            I => \N__8058\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8058\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__8063\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__8058\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1579\ : InMux
    port map (
            O => \N__8053\,
            I => \receive_module.rx_counter.n1840\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8045\
        );

    \I__1577\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8042\
        );

    \I__1576\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8039\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8045\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__8042\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__8039\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1572\ : InMux
    port map (
            O => \N__8032\,
            I => \receive_module.rx_counter.n1841\
        );

    \I__1571\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8026\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__8026\,
            I => \N__8022\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8017\
        );

    \I__1568\ : Span4Mux_h
    port map (
            O => \N__8022\,
            I => \N__8014\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8021\,
            I => \N__8009\
        );

    \I__1566\ : InMux
    port map (
            O => \N__8020\,
            I => \N__8009\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__8017\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__8014\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__8009\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__1562\ : InMux
    port map (
            O => \N__8002\,
            I => \receive_module.rx_counter.n1842\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7999\,
            I => \bfn_7_7_0_\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7993\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7993\,
            I => \N__7989\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7984\
        );

    \I__1557\ : Span4Mux_h
    port map (
            O => \N__7989\,
            I => \N__7981\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7978\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7975\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__7984\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__7981\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7978\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7975\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__1550\ : CEMux
    port map (
            O => \N__7966\,
            I => \N__7962\
        );

    \I__1549\ : CEMux
    port map (
            O => \N__7965\,
            I => \N__7959\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7962\,
            I => \N__7956\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7959\,
            I => \N__7953\
        );

    \I__1546\ : Span4Mux_h
    port map (
            O => \N__7956\,
            I => \N__7950\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__7953\,
            I => \receive_module.rx_counter.n752\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__7950\,
            I => \receive_module.rx_counter.n752\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7942\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7942\,
            I => \transmit_module.Y_DELTA_PATTERN_28\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7936\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7936\,
            I => \transmit_module.Y_DELTA_PATTERN_27\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7933\,
            I => \N__7930\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7930\,
            I => \transmit_module.Y_DELTA_PATTERN_26\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7927\,
            I => \N__7924\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7924\,
            I => \transmit_module.Y_DELTA_PATTERN_6\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7921\,
            I => \N__7918\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7918\,
            I => \transmit_module.Y_DELTA_PATTERN_25\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7912\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7912\,
            I => \transmit_module.Y_DELTA_PATTERN_24\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7906\,
            I => \N__7903\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__7903\,
            I => \transmit_module.Y_DELTA_PATTERN_23\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7897\,
            I => \transmit_module.Y_DELTA_PATTERN_1\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7890\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7887\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7890\,
            I => \N__7883\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7887\,
            I => \N__7880\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7877\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__7883\,
            I => \N__7872\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__7880\,
            I => \N__7872\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7877\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__7872\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7867\,
            I => \N__7864\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7864\,
            I => \N__7859\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7863\,
            I => \N__7854\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7854\
        );

    \I__1513\ : Span4Mux_v
    port map (
            O => \N__7859\,
            I => \N__7849\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7854\,
            I => \N__7849\
        );

    \I__1511\ : Sp12to4
    port map (
            O => \N__7849\,
            I => \N__7846\
        );

    \I__1510\ : Span12Mux_h
    port map (
            O => \N__7846\,
            I => \N__7843\
        );

    \I__1509\ : Odrv12
    port map (
            O => \N__7843\,
            I => \TVP_HSYNC_c\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7837\,
            I => \receive_module.rx_counter.old_HS\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7829\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7824\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7824\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7829\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7824\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7819\,
            I => \bfn_7_6_0_\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7813\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7813\,
            I => \transmit_module.Y_DELTA_PATTERN_20\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7807\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7807\,
            I => \transmit_module.Y_DELTA_PATTERN_19\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7801\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7801\,
            I => \transmit_module.Y_DELTA_PATTERN_18\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7795\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7795\,
            I => \transmit_module.Y_DELTA_PATTERN_22\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7792\,
            I => \N__7789\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7789\,
            I => \transmit_module.Y_DELTA_PATTERN_21\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7783\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7783\,
            I => \transmit_module.Y_DELTA_PATTERN_17\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7780\,
            I => \N__7777\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7777\,
            I => \N__7774\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__7774\,
            I => \transmit_module.Y_DELTA_PATTERN_29\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7768\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7768\,
            I => \transmit_module.X_DELTA_PATTERN_7\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7765\,
            I => \N__7762\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7762\,
            I => \transmit_module.X_DELTA_PATTERN_9\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7756\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7756\,
            I => \transmit_module.X_DELTA_PATTERN_8\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7750\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7750\,
            I => \transmit_module.X_DELTA_PATTERN_15\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7744\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7744\,
            I => \transmit_module.X_DELTA_PATTERN_6\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7738\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7738\,
            I => \transmit_module.X_DELTA_PATTERN_5\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7732\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7732\,
            I => \transmit_module.X_DELTA_PATTERN_14\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7726\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7726\,
            I => \N__7723\
        );

    \I__1469\ : Span4Mux_h
    port map (
            O => \N__7723\,
            I => \N__7720\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__7720\,
            I => \N__7717\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__7717\,
            I => \transmit_module.Y_DELTA_PATTERN_33\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7711\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7711\,
            I => \transmit_module.Y_DELTA_PATTERN_32\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7705\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7705\,
            I => \transmit_module.Y_DELTA_PATTERN_31\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7699\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7699\,
            I => \transmit_module.Y_DELTA_PATTERN_30\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7692\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7689\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7692\,
            I => \transmit_module.BRAM_ADDR_12\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7689\,
            I => \transmit_module.BRAM_ADDR_12\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__7684\,
            I => \N__7681\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7678\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7678\,
            I => \transmit_module.ADDR_Y_COMPONENT_12\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7675\,
            I => \N__7671\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7674\,
            I => \N__7668\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7671\,
            I => \N__7665\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7668\,
            I => \transmit_module.BRAM_ADDR_2\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__7665\,
            I => \transmit_module.BRAM_ADDR_2\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__7660\,
            I => \N__7657\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7654\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7654\,
            I => \transmit_module.ADDR_Y_COMPONENT_2\
        );

    \I__1445\ : CEMux
    port map (
            O => \N__7651\,
            I => \N__7646\
        );

    \I__1444\ : CEMux
    port map (
            O => \N__7650\,
            I => \N__7642\
        );

    \I__1443\ : CEMux
    port map (
            O => \N__7649\,
            I => \N__7638\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7646\,
            I => \N__7635\
        );

    \I__1441\ : CEMux
    port map (
            O => \N__7645\,
            I => \N__7632\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7642\,
            I => \N__7629\
        );

    \I__1439\ : CEMux
    port map (
            O => \N__7641\,
            I => \N__7626\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7638\,
            I => \N__7623\
        );

    \I__1437\ : Span4Mux_h
    port map (
            O => \N__7635\,
            I => \N__7618\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7632\,
            I => \N__7618\
        );

    \I__1435\ : Span4Mux_h
    port map (
            O => \N__7629\,
            I => \N__7613\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7626\,
            I => \N__7613\
        );

    \I__1433\ : Span4Mux_v
    port map (
            O => \N__7623\,
            I => \N__7610\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__7618\,
            I => \N__7605\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__7613\,
            I => \N__7605\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__7610\,
            I => \transmit_module.n792\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__7605\,
            I => \transmit_module.n792\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7597\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7597\,
            I => \transmit_module.X_DELTA_PATTERN_2\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7591\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7591\,
            I => \transmit_module.X_DELTA_PATTERN_4\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7585\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7585\,
            I => \transmit_module.X_DELTA_PATTERN_3\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7579\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7579\,
            I => \transmit_module.X_DELTA_PATTERN_1\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__7576\,
            I => \N__7573\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7573\,
            I => \N__7570\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7570\,
            I => \N__7566\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7563\
        );

    \I__1416\ : Span4Mux_h
    port map (
            O => \N__7566\,
            I => \N__7560\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7563\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__7560\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7555\,
            I => \N__7551\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7554\,
            I => \N__7548\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__7551\,
            I => \transmit_module.BRAM_ADDR_1\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__7548\,
            I => \transmit_module.BRAM_ADDR_1\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7537\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7537\,
            I => \transmit_module.ADDR_Y_COMPONENT_1\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7530\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7527\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7530\,
            I => \transmit_module.BRAM_ADDR_10\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7527\,
            I => \transmit_module.BRAM_ADDR_10\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7519\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7519\,
            I => \transmit_module.ADDR_Y_COMPONENT_10\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7512\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7509\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7512\,
            I => \transmit_module.BRAM_ADDR_5\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7509\,
            I => \transmit_module.BRAM_ADDR_5\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7501\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7501\,
            I => \N__7498\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__7498\,
            I => \transmit_module.ADDR_Y_COMPONENT_5\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7495\,
            I => \N__7491\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7494\,
            I => \N__7488\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7491\,
            I => \transmit_module.BRAM_ADDR_8\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7488\,
            I => \transmit_module.BRAM_ADDR_8\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7483\,
            I => \N__7480\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7480\,
            I => \N__7477\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7477\,
            I => \transmit_module.ADDR_Y_COMPONENT_8\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7470\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7473\,
            I => \N__7467\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__7470\,
            I => \transmit_module.BRAM_ADDR_11\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7467\,
            I => \transmit_module.BRAM_ADDR_11\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__7462\,
            I => \N__7459\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7459\,
            I => \N__7456\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7456\,
            I => \transmit_module.ADDR_Y_COMPONENT_11\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7453\,
            I => \N__7449\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7452\,
            I => \N__7446\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7449\,
            I => \N__7443\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7446\,
            I => \transmit_module.BRAM_ADDR_0\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__7443\,
            I => \transmit_module.BRAM_ADDR_0\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7435\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7435\,
            I => \transmit_module.ADDR_Y_COMPONENT_0\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7429\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7429\,
            I => \N__7425\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7428\,
            I => \N__7422\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__7425\,
            I => \transmit_module.BRAM_ADDR_3\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7422\,
            I => \transmit_module.BRAM_ADDR_3\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7414\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7414\,
            I => \N__7411\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__7411\,
            I => \transmit_module.ADDR_Y_COMPONENT_3\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__7408\,
            I => \receive_module.rx_counter.n2007_cascade_\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__7405\,
            I => \receive_module.rx_counter.n2069_cascade_\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7396\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7396\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7396\,
            I => \receive_module.rx_counter.n2153\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7390\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7390\,
            I => \receive_module.rx_counter.n2071\
        );

    \I__1357\ : SRMux
    port map (
            O => \N__7387\,
            I => \N__7383\
        );

    \I__1356\ : SRMux
    port map (
            O => \N__7386\,
            I => \N__7380\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7383\,
            I => \N__7377\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7380\,
            I => \N__7374\
        );

    \I__1353\ : Span4Mux_v
    port map (
            O => \N__7377\,
            I => \N__7371\
        );

    \I__1352\ : Span4Mux_v
    port map (
            O => \N__7374\,
            I => \N__7368\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__7371\,
            I => n2148
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__7368\,
            I => n2148
        );

    \I__1349\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7360\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7360\,
            I => \transmit_module.n199\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7354\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7354\,
            I => \transmit_module.n203\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7348\,
            I => \N__7345\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__7345\,
            I => \transmit_module.ADDR_Y_COMPONENT_6\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7339\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__7339\,
            I => \transmit_module.n198\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7332\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7329\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7332\,
            I => \transmit_module.BRAM_ADDR_6\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7329\,
            I => \transmit_module.BRAM_ADDR_6\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7321\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7321\,
            I => \transmit_module.n201\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7315\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7315\,
            I => \transmit_module.Y_DELTA_PATTERN_5\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7312\,
            I => \N__7309\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7309\,
            I => \transmit_module.Y_DELTA_PATTERN_4\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7303\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7303\,
            I => \transmit_module.Y_DELTA_PATTERN_3\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7300\,
            I => \N__7297\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__7297\,
            I => \transmit_module.Y_DELTA_PATTERN_2\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__7294\,
            I => \N__7291\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7288\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7288\,
            I => \N__7285\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__7285\,
            I => \receive_module.rx_counter.n8\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7279\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__7279\,
            I => \receive_module.rx_counter.n7_adj_574\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__7276\,
            I => \receive_module.rx_counter.n2063_cascade_\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7270\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7270\,
            I => \receive_module.rx_counter.n4\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7264\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7264\,
            I => \receive_module.rx_counter.n2007\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7255\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7248\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7248\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7245\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7255\,
            I => \N__7242\
        );

    \I__1310\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7237\
        );

    \I__1309\ : InMux
    port map (
            O => \N__7253\,
            I => \N__7237\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7248\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__7245\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__7242\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7237\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1304\ : IoInMux
    port map (
            O => \N__7228\,
            I => \N__7225\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7225\,
            I => \N__7222\
        );

    \I__1302\ : IoSpan4Mux
    port map (
            O => \N__7222\,
            I => \N__7219\
        );

    \I__1301\ : Span4Mux_s3_v
    port map (
            O => \N__7219\,
            I => \N__7216\
        );

    \I__1300\ : Span4Mux_v
    port map (
            O => \N__7216\,
            I => \N__7213\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__7213\,
            I => \N__7210\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__7210\,
            I => \ADV_G_c_7\
        );

    \I__1297\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7203\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7199\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7203\,
            I => \N__7196\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7193\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7199\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__7196\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__7193\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__1290\ : IoInMux
    port map (
            O => \N__7186\,
            I => \N__7183\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__7183\,
            I => \N__7180\
        );

    \I__1288\ : Span4Mux_s2_v
    port map (
            O => \N__7180\,
            I => \N__7177\
        );

    \I__1287\ : Span4Mux_v
    port map (
            O => \N__7177\,
            I => \N__7174\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__7174\,
            I => \N__7171\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__7171\,
            I => \ADV_G_c_1\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__7168\,
            I => \N__7163\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7159\
        );

    \I__1282\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7152\
        );

    \I__1281\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7152\
        );

    \I__1280\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7149\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__7159\,
            I => \N__7146\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7158\,
            I => \N__7141\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7141\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7152\,
            I => \N__7138\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__7149\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__7146\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__7141\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__7138\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1271\ : IoInMux
    port map (
            O => \N__7129\,
            I => \N__7126\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__7126\,
            I => \N__7123\
        );

    \I__1269\ : Span4Mux_s3_v
    port map (
            O => \N__7123\,
            I => \N__7120\
        );

    \I__1268\ : Span4Mux_h
    port map (
            O => \N__7120\,
            I => \N__7117\
        );

    \I__1267\ : Span4Mux_v
    port map (
            O => \N__7117\,
            I => \N__7114\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__7114\,
            I => \ADV_G_c_5\
        );

    \I__1265\ : InMux
    port map (
            O => \N__7111\,
            I => \N__7107\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__7110\,
            I => \N__7102\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7107\,
            I => \N__7099\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7092\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7105\,
            I => \N__7089\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7086\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__7099\,
            I => \N__7083\
        );

    \I__1258\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7078\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7078\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7096\,
            I => \N__7073\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7095\,
            I => \N__7073\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__7092\,
            I => \VGA_Y_6\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7089\,
            I => \VGA_Y_6\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__7086\,
            I => \VGA_Y_6\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__7083\,
            I => \VGA_Y_6\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__7078\,
            I => \VGA_Y_6\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__7073\,
            I => \VGA_Y_6\
        );

    \I__1248\ : IoInMux
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__7057\,
            I => \N__7054\
        );

    \I__1246\ : Span4Mux_s2_v
    port map (
            O => \N__7054\,
            I => \N__7051\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__7048\,
            I => \N__7045\
        );

    \I__1243\ : Sp12to4
    port map (
            O => \N__7045\,
            I => \N__7042\
        );

    \I__1242\ : Span12Mux_h
    port map (
            O => \N__7042\,
            I => \N__7039\
        );

    \I__1241\ : Odrv12
    port map (
            O => \N__7039\,
            I => \ADV_B_c_6\
        );

    \I__1240\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7032\
        );

    \I__1239\ : InMux
    port map (
            O => \N__7035\,
            I => \N__7028\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__7032\,
            I => \N__7025\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7019\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__7028\,
            I => \N__7016\
        );

    \I__1235\ : Span4Mux_h
    port map (
            O => \N__7025\,
            I => \N__7013\
        );

    \I__1234\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7010\
        );

    \I__1233\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7005\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7005\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__7019\,
            I => \VGA_Y_7\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__7016\,
            I => \VGA_Y_7\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__7013\,
            I => \VGA_Y_7\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__7010\,
            I => \VGA_Y_7\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__7005\,
            I => \VGA_Y_7\
        );

    \I__1226\ : IoInMux
    port map (
            O => \N__6994\,
            I => \N__6991\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6991\,
            I => \N__6988\
        );

    \I__1224\ : Span4Mux_s3_h
    port map (
            O => \N__6988\,
            I => \N__6985\
        );

    \I__1223\ : Span4Mux_v
    port map (
            O => \N__6985\,
            I => \N__6982\
        );

    \I__1222\ : Span4Mux_v
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1221\ : Odrv4
    port map (
            O => \N__6979\,
            I => \ADV_R_c_7\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6973\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6973\,
            I => \N__6968\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__6972\,
            I => \N__6961\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6958\
        );

    \I__1216\ : Span4Mux_h
    port map (
            O => \N__6968\,
            I => \N__6955\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6952\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6949\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6946\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6964\,
            I => \N__6941\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6941\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6958\,
            I => \VGA_Y_2\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__6955\,
            I => \VGA_Y_2\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6952\,
            I => \VGA_Y_2\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6949\,
            I => \VGA_Y_2\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6946\,
            I => \VGA_Y_2\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6941\,
            I => \VGA_Y_2\
        );

    \I__1204\ : IoInMux
    port map (
            O => \N__6928\,
            I => \N__6925\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6925\,
            I => \N__6922\
        );

    \I__1202\ : IoSpan4Mux
    port map (
            O => \N__6922\,
            I => \N__6919\
        );

    \I__1201\ : Span4Mux_s3_v
    port map (
            O => \N__6919\,
            I => \N__6916\
        );

    \I__1200\ : Sp12to4
    port map (
            O => \N__6916\,
            I => \N__6913\
        );

    \I__1199\ : Span12Mux_h
    port map (
            O => \N__6913\,
            I => \N__6910\
        );

    \I__1198\ : Odrv12
    port map (
            O => \N__6910\,
            I => \ADV_B_c_2\
        );

    \I__1197\ : SRMux
    port map (
            O => \N__6907\,
            I => \N__6902\
        );

    \I__1196\ : SRMux
    port map (
            O => \N__6906\,
            I => \N__6899\
        );

    \I__1195\ : SRMux
    port map (
            O => \N__6905\,
            I => \N__6896\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6902\,
            I => \N__6893\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6899\,
            I => \N__6890\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6896\,
            I => \N__6886\
        );

    \I__1191\ : Span4Mux_h
    port map (
            O => \N__6893\,
            I => \N__6883\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__6890\,
            I => \N__6878\
        );

    \I__1189\ : SRMux
    port map (
            O => \N__6889\,
            I => \N__6875\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__6886\,
            I => \N__6872\
        );

    \I__1187\ : Span4Mux_s0_h
    port map (
            O => \N__6883\,
            I => \N__6869\
        );

    \I__1186\ : SRMux
    port map (
            O => \N__6882\,
            I => \N__6866\
        );

    \I__1185\ : SRMux
    port map (
            O => \N__6881\,
            I => \N__6863\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__6878\,
            I => n1144
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6875\,
            I => n1144
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__6872\,
            I => n1144
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__6869\,
            I => n1144
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6866\,
            I => n1144
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6863\,
            I => n1144
        );

    \I__1178\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6847\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6847\,
            I => \N__6844\
        );

    \I__1176\ : Span4Mux_h
    port map (
            O => \N__6844\,
            I => \N__6841\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__6841\,
            I => \transmit_module.Y_DELTA_PATTERN_99\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6838\,
            I => \bfn_5_20_0_\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6832\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6832\,
            I => \N__6824\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6821\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6830\,
            I => \N__6814\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6814\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6814\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6827\,
            I => \N__6811\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__6824\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6821\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6814\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6811\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6802\,
            I => \transmit_module.video_signal_controller.n1852\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6799\,
            I => \transmit_module.video_signal_controller.n1853\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6796\,
            I => \N__6792\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6785\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6792\,
            I => \N__6782\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6775\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6775\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6775\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6772\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6785\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6782\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6775\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6772\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1149\ : CEMux
    port map (
            O => \N__6763\,
            I => \N__6759\
        );

    \I__1148\ : CEMux
    port map (
            O => \N__6762\,
            I => \N__6755\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6759\,
            I => \N__6752\
        );

    \I__1146\ : SRMux
    port map (
            O => \N__6758\,
            I => \N__6749\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6755\,
            I => \N__6745\
        );

    \I__1144\ : Span4Mux_v
    port map (
            O => \N__6752\,
            I => \N__6740\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6749\,
            I => \N__6740\
        );

    \I__1142\ : SRMux
    port map (
            O => \N__6748\,
            I => \N__6737\
        );

    \I__1141\ : Span4Mux_v
    port map (
            O => \N__6745\,
            I => \N__6731\
        );

    \I__1140\ : Span4Mux_h
    port map (
            O => \N__6740\,
            I => \N__6728\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6737\,
            I => \N__6725\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6718\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6718\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6718\
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__6731\,
            I => \transmit_module.video_signal_controller.n528\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__6728\,
            I => \transmit_module.video_signal_controller.n528\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__6725\,
            I => \transmit_module.video_signal_controller.n528\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6718\,
            I => \transmit_module.video_signal_controller.n528\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6705\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6708\,
            I => \N__6701\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6705\,
            I => \N__6698\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6704\,
            I => \N__6695\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6701\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__6698\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6695\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__1124\ : IoInMux
    port map (
            O => \N__6688\,
            I => \N__6685\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6685\,
            I => \N__6682\
        );

    \I__1122\ : Span4Mux_s3_v
    port map (
            O => \N__6682\,
            I => \N__6679\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__6676\,
            I => \N__6673\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__6673\,
            I => \ADV_G_c_2\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6670\,
            I => \N__6666\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6658\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6666\,
            I => \N__6655\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6665\,
            I => \N__6652\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6664\,
            I => \N__6647\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6663\,
            I => \N__6647\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6644\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6641\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6658\,
            I => \VGA_Y_4\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__6655\,
            I => \VGA_Y_4\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6652\,
            I => \VGA_Y_4\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6647\,
            I => \VGA_Y_4\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6644\,
            I => \VGA_Y_4\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6641\,
            I => \VGA_Y_4\
        );

    \I__1104\ : IoInMux
    port map (
            O => \N__6628\,
            I => \N__6625\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1102\ : IoSpan4Mux
    port map (
            O => \N__6622\,
            I => \N__6619\
        );

    \I__1101\ : Span4Mux_s2_v
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1100\ : Span4Mux_h
    port map (
            O => \N__6616\,
            I => \N__6613\
        );

    \I__1099\ : Sp12to4
    port map (
            O => \N__6613\,
            I => \N__6610\
        );

    \I__1098\ : Span12Mux_h
    port map (
            O => \N__6610\,
            I => \N__6607\
        );

    \I__1097\ : Odrv12
    port map (
            O => \N__6607\,
            I => \ADV_B_c_4\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6599\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__6603\,
            I => \N__6594\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6602\,
            I => \N__6591\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6599\,
            I => \N__6588\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6585\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6597\,
            I => \N__6582\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6579\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6591\,
            I => \VGA_Y_0\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__6588\,
            I => \VGA_Y_0\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6585\,
            I => \VGA_Y_0\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6582\,
            I => \VGA_Y_0\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6579\,
            I => \VGA_Y_0\
        );

    \I__1084\ : IoInMux
    port map (
            O => \N__6568\,
            I => \N__6565\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6565\,
            I => \N__6562\
        );

    \I__1082\ : Span12Mux_s11_v
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__6559\,
            I => \ADV_B_c_0\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6552\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6546\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6552\,
            I => \N__6543\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6538\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6538\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6535\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6546\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__6543\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6538\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6535\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1070\ : IoInMux
    port map (
            O => \N__6526\,
            I => \N__6523\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__1068\ : Span12Mux_s11_v
    port map (
            O => \N__6520\,
            I => \N__6517\
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__6517\,
            I => \ADV_G_c_4\
        );

    \I__1066\ : IoInMux
    port map (
            O => \N__6514\,
            I => \N__6511\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__6511\,
            I => \N__6508\
        );

    \I__1064\ : IoSpan4Mux
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__1063\ : Span4Mux_s0_v
    port map (
            O => \N__6505\,
            I => \N__6502\
        );

    \I__1062\ : Sp12to4
    port map (
            O => \N__6502\,
            I => \N__6499\
        );

    \I__1061\ : Span12Mux_s11_v
    port map (
            O => \N__6499\,
            I => \N__6496\
        );

    \I__1060\ : Span12Mux_h
    port map (
            O => \N__6496\,
            I => \N__6493\
        );

    \I__1059\ : Odrv12
    port map (
            O => \N__6493\,
            I => \ADV_B_c_7\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6486\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6482\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6486\,
            I => \N__6475\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6472\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6482\,
            I => \N__6469\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6464\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6464\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6459\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6459\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__6475\,
            I => \VGA_Y_1\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6472\,
            I => \VGA_Y_1\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__6469\,
            I => \VGA_Y_1\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6464\,
            I => \VGA_Y_1\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6459\,
            I => \VGA_Y_1\
        );

    \I__1044\ : IoInMux
    port map (
            O => \N__6448\,
            I => \N__6445\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6445\,
            I => \N__6442\
        );

    \I__1042\ : Span12Mux_s11_v
    port map (
            O => \N__6442\,
            I => \N__6439\
        );

    \I__1041\ : Span12Mux_h
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__1040\ : Odrv12
    port map (
            O => \N__6436\,
            I => \ADV_B_c_1\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6428\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6425\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6431\,
            I => \N__6422\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6428\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6425\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6422\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6415\,
            I => \bfn_5_19_0_\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6412\,
            I => \transmit_module.video_signal_controller.n1844\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6409\,
            I => \transmit_module.video_signal_controller.n1845\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6403\,
            I => \N__6398\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6394\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6391\
        );

    \I__1026\ : Span4Mux_v
    port map (
            O => \N__6398\,
            I => \N__6388\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6385\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6394\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6391\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__6388\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6385\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6376\,
            I => \transmit_module.video_signal_controller.n1846\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6373\,
            I => \transmit_module.video_signal_controller.n1847\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6370\,
            I => \transmit_module.video_signal_controller.n1848\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6363\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6358\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6363\,
            I => \N__6355\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6348\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6348\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6358\,
            I => \N__6343\
        );

    \I__1011\ : Span4Mux_v
    port map (
            O => \N__6355\,
            I => \N__6343\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6354\,
            I => \N__6338\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6338\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6348\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__6343\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6338\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6331\,
            I => \transmit_module.video_signal_controller.n1849\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6328\,
            I => \transmit_module.video_signal_controller.n1850\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6319\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6316\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6323\,
            I => \N__6313\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6310\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__6319\,
            I => \N__6305\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6305\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6313\,
            I => \N__6302\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6310\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__6305\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__6302\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__993\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__991\ : Odrv12
    port map (
            O => \N__6289\,
            I => \transmit_module.n204\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__6286\,
            I => \N__6283\
        );

    \I__989\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6280\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6280\,
            I => \transmit_module.ADDR_Y_COMPONENT_9\
        );

    \I__987\ : InMux
    port map (
            O => \N__6277\,
            I => \N__6274\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__6274\,
            I => \transmit_module.n195\
        );

    \I__985\ : InMux
    port map (
            O => \N__6271\,
            I => \N__6265\
        );

    \I__984\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6265\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6265\,
            I => \transmit_module.BRAM_ADDR_9\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__6262\,
            I => \N__6259\
        );

    \I__981\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6256\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6256\,
            I => \transmit_module.n194\
        );

    \I__979\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6250\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6250\,
            I => \N__6247\
        );

    \I__977\ : Odrv12
    port map (
            O => \N__6247\,
            I => \transmit_module.n202\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__6244\,
            I => \transmit_module.n2145_cascade_\
        );

    \I__975\ : IoInMux
    port map (
            O => \N__6241\,
            I => \N__6238\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__6238\,
            I => \N__6235\
        );

    \I__973\ : Span4Mux_s3_h
    port map (
            O => \N__6235\,
            I => \N__6232\
        );

    \I__972\ : Span4Mux_v
    port map (
            O => \N__6232\,
            I => \N__6228\
        );

    \I__971\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6225\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__6228\,
            I => n2144
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6225\,
            I => n2144
        );

    \I__968\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6211\
        );

    \I__967\ : InMux
    port map (
            O => \N__6219\,
            I => \N__6211\
        );

    \I__966\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6206\
        );

    \I__965\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6206\
        );

    \I__964\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6203\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6211\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6206\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__6203\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__960\ : IoInMux
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6193\,
            I => \N__6189\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__6192\,
            I => \N__6182\
        );

    \I__957\ : Span4Mux_s3_h
    port map (
            O => \N__6189\,
            I => \N__6178\
        );

    \I__956\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6175\
        );

    \I__955\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6170\
        );

    \I__954\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6170\
        );

    \I__953\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6163\
        );

    \I__952\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6163\
        );

    \I__951\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6163\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__6178\,
            I => \ADV_HSYNC_c\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6175\,
            I => \ADV_HSYNC_c\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__6170\,
            I => \ADV_HSYNC_c\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__6163\,
            I => \ADV_HSYNC_c\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__6154\,
            I => \transmit_module.n2156_cascade_\
        );

    \I__945\ : InMux
    port map (
            O => \N__6151\,
            I => \bfn_5_16_0_\
        );

    \I__944\ : InMux
    port map (
            O => \N__6148\,
            I => \transmit_module.n1831\
        );

    \I__943\ : InMux
    port map (
            O => \N__6145\,
            I => \transmit_module.n1832\
        );

    \I__942\ : InMux
    port map (
            O => \N__6142\,
            I => \transmit_module.n1833\
        );

    \I__941\ : InMux
    port map (
            O => \N__6139\,
            I => \transmit_module.n1834\
        );

    \I__940\ : InMux
    port map (
            O => \N__6136\,
            I => \transmit_module.n1835\
        );

    \I__939\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6130\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__6130\,
            I => \transmit_module.n193\
        );

    \I__937\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6124\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6124\,
            I => \transmit_module.n196\
        );

    \I__935\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6118\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__6118\,
            I => \transmit_module.n192\
        );

    \I__933\ : InMux
    port map (
            O => \N__6115\,
            I => \transmit_module.n1823\
        );

    \I__932\ : InMux
    port map (
            O => \N__6112\,
            I => \transmit_module.n1824\
        );

    \I__931\ : InMux
    port map (
            O => \N__6109\,
            I => \transmit_module.n1825\
        );

    \I__930\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6102\
        );

    \I__929\ : InMux
    port map (
            O => \N__6105\,
            I => \N__6099\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6102\,
            I => \transmit_module.BRAM_ADDR_4\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__6099\,
            I => \transmit_module.BRAM_ADDR_4\
        );

    \I__926\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6091\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__6091\,
            I => \transmit_module.n200\
        );

    \I__924\ : InMux
    port map (
            O => \N__6088\,
            I => \transmit_module.n1826\
        );

    \I__923\ : InMux
    port map (
            O => \N__6085\,
            I => \transmit_module.n1827\
        );

    \I__922\ : InMux
    port map (
            O => \N__6082\,
            I => \transmit_module.n1828\
        );

    \I__921\ : InMux
    port map (
            O => \N__6079\,
            I => \transmit_module.n1829\
        );

    \I__920\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6073\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__6073\,
            I => \receive_module.rx_counter.n8_adj_575\
        );

    \I__918\ : InMux
    port map (
            O => \N__6070\,
            I => \receive_module.rx_counter.n1871\
        );

    \I__917\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6063\
        );

    \I__916\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6060\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__6063\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__6060\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__913\ : InMux
    port map (
            O => \N__6055\,
            I => \receive_module.rx_counter.n1872\
        );

    \I__912\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6048\
        );

    \I__911\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6045\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__6048\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__6045\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__908\ : InMux
    port map (
            O => \N__6040\,
            I => \receive_module.rx_counter.n1873\
        );

    \I__907\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6033\
        );

    \I__906\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6030\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6033\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__6030\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__903\ : InMux
    port map (
            O => \N__6025\,
            I => \receive_module.rx_counter.n1874\
        );

    \I__902\ : InMux
    port map (
            O => \N__6022\,
            I => \N__6015\
        );

    \I__901\ : InMux
    port map (
            O => \N__6021\,
            I => \N__6015\
        );

    \I__900\ : InMux
    port map (
            O => \N__6020\,
            I => \N__6012\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6015\,
            I => \N__6009\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__6012\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__6009\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__896\ : InMux
    port map (
            O => \N__6004\,
            I => \receive_module.rx_counter.n1875\
        );

    \I__895\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5994\
        );

    \I__894\ : InMux
    port map (
            O => \N__6000\,
            I => \N__5994\
        );

    \I__893\ : InMux
    port map (
            O => \N__5999\,
            I => \N__5991\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5994\,
            I => \N__5988\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5991\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__5988\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__889\ : InMux
    port map (
            O => \N__5983\,
            I => \receive_module.rx_counter.n1876\
        );

    \I__888\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5977\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5977\,
            I => \N__5973\
        );

    \I__886\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5970\
        );

    \I__885\ : Span4Mux_h
    port map (
            O => \N__5973\,
            I => \N__5967\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5970\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__5967\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__882\ : InMux
    port map (
            O => \N__5962\,
            I => \bfn_5_12_0_\
        );

    \I__881\ : InMux
    port map (
            O => \N__5959\,
            I => \receive_module.rx_counter.n1878\
        );

    \I__880\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5952\
        );

    \I__879\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5949\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5952\,
            I => \N__5946\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5949\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__5946\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__5941\,
            I => \N__5938\
        );

    \I__874\ : InMux
    port map (
            O => \N__5938\,
            I => \N__5935\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5935\,
            I => \transmit_module.ADDR_Y_COMPONENT_4\
        );

    \I__872\ : IoInMux
    port map (
            O => \N__5932\,
            I => \N__5929\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5929\,
            I => \N__5925\
        );

    \I__870\ : InMux
    port map (
            O => \N__5928\,
            I => \N__5922\
        );

    \I__869\ : IoSpan4Mux
    port map (
            O => \N__5925\,
            I => \N__5919\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5922\,
            I => \N__5916\
        );

    \I__867\ : Span4Mux_s3_h
    port map (
            O => \N__5919\,
            I => \N__5911\
        );

    \I__866\ : Span4Mux_v
    port map (
            O => \N__5916\,
            I => \N__5911\
        );

    \I__865\ : Span4Mux_v
    port map (
            O => \N__5911\,
            I => \N__5908\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__5908\,
            I => \N__5905\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__5905\,
            I => \DEBUG_c_5\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__5902\,
            I => \receive_module.rx_counter.n28_cascade_\
        );

    \I__861\ : IoInMux
    port map (
            O => \N__5899\,
            I => \N__5896\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__859\ : Span4Mux_s2_h
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__5890\,
            I => \N__5887\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__5884\,
            I => \DEBUG_c_4\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__5881\,
            I => \DEBUG_c_4_cascade_\
        );

    \I__854\ : CEMux
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5875\,
            I => \N__5871\
        );

    \I__852\ : CEMux
    port map (
            O => \N__5874\,
            I => \N__5868\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__5871\,
            I => \N__5865\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5868\,
            I => \N__5862\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__5865\,
            I => \receive_module.n788\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__5862\,
            I => \receive_module.n788\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__5857\,
            I => \N__5854\
        );

    \I__846\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5851\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5851\,
            I => \receive_module.rx_counter.n2083\
        );

    \I__844\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5845\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5845\,
            I => \receive_module.rx_counter.n2033\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__5842\,
            I => \N__5839\
        );

    \I__841\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5833\
        );

    \I__840\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5833\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5833\,
            I => \receive_module.rx_counter.n1981\
        );

    \I__838\ : InMux
    port map (
            O => \N__5830\,
            I => \N__5827\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5827\,
            I => \receive_module.rx_counter.n10\
        );

    \I__836\ : InMux
    port map (
            O => \N__5824\,
            I => \bfn_5_11_0_\
        );

    \I__835\ : InMux
    port map (
            O => \N__5821\,
            I => \N__5818\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5818\,
            I => \receive_module.rx_counter.n9\
        );

    \I__833\ : InMux
    port map (
            O => \N__5815\,
            I => \receive_module.rx_counter.n1870\
        );

    \I__832\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5806\
        );

    \I__831\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5806\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5803\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__5803\,
            I => \transmit_module.video_signal_controller.n679\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__5800\,
            I => \transmit_module.video_signal_controller.n679_cascade_\
        );

    \I__827\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5794\,
            I => \transmit_module.video_signal_controller.n2151\
        );

    \I__825\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5788\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5788\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_552\
        );

    \I__823\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5775\
        );

    \I__822\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5770\
        );

    \I__821\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5770\
        );

    \I__820\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5763\
        );

    \I__819\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5763\
        );

    \I__818\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5763\
        );

    \I__817\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5758\
        );

    \I__816\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5758\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5775\,
            I => \VGA_Y_5\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5770\,
            I => \VGA_Y_5\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5763\,
            I => \VGA_Y_5\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5758\,
            I => \VGA_Y_5\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__5749\,
            I => \transmit_module.video_signal_controller.n2149_cascade_\
        );

    \I__810\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5743\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5743\,
            I => \transmit_module.video_signal_controller.n2152\
        );

    \I__808\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5737\,
            I => \transmit_module.video_signal_controller.n2006\
        );

    \I__806\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5731\,
            I => \transmit_module.video_signal_controller.n8\
        );

    \I__804\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5725\,
            I => \transmit_module.video_signal_controller.n2140\
        );

    \I__802\ : IoInMux
    port map (
            O => \N__5722\,
            I => \N__5719\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5719\,
            I => \N__5716\
        );

    \I__800\ : Span12Mux_s9_v
    port map (
            O => \N__5716\,
            I => \N__5713\
        );

    \I__799\ : Odrv12
    port map (
            O => \N__5713\,
            I => \ADV_G_c_3\
        );

    \I__798\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5706\
        );

    \I__797\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5698\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5706\,
            I => \N__5695\
        );

    \I__795\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5692\
        );

    \I__794\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5687\
        );

    \I__793\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5687\
        );

    \I__792\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5682\
        );

    \I__791\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5682\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5698\,
            I => \VGA_Y_3\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__5695\,
            I => \VGA_Y_3\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5692\,
            I => \VGA_Y_3\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5687\,
            I => \VGA_Y_3\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5682\,
            I => \VGA_Y_3\
        );

    \I__785\ : IoInMux
    port map (
            O => \N__5671\,
            I => \N__5668\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__783\ : Span4Mux_s1_v
    port map (
            O => \N__5665\,
            I => \N__5662\
        );

    \I__782\ : Span4Mux_v
    port map (
            O => \N__5662\,
            I => \N__5659\
        );

    \I__781\ : Span4Mux_v
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__780\ : Sp12to4
    port map (
            O => \N__5656\,
            I => \N__5653\
        );

    \I__779\ : Span12Mux_h
    port map (
            O => \N__5653\,
            I => \N__5650\
        );

    \I__778\ : Odrv12
    port map (
            O => \N__5650\,
            I => \ADV_B_c_3\
        );

    \I__777\ : IoInMux
    port map (
            O => \N__5647\,
            I => \N__5644\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5644\,
            I => \N__5641\
        );

    \I__775\ : Span12Mux_s0_v
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__774\ : Span12Mux_v
    port map (
            O => \N__5638\,
            I => \N__5635\
        );

    \I__773\ : Span12Mux_h
    port map (
            O => \N__5635\,
            I => \N__5632\
        );

    \I__772\ : Odrv12
    port map (
            O => \N__5632\,
            I => \ADV_B_c_5\
        );

    \I__771\ : IoInMux
    port map (
            O => \N__5629\,
            I => \N__5626\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5626\,
            I => \N__5623\
        );

    \I__769\ : IoSpan4Mux
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__768\ : Sp12to4
    port map (
            O => \N__5620\,
            I => \N__5617\
        );

    \I__767\ : Span12Mux_v
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__766\ : Odrv12
    port map (
            O => \N__5614\,
            I => \ADV_G_c_0\
        );

    \I__765\ : IoInMux
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5608\,
            I => \N__5605\
        );

    \I__763\ : Span4Mux_s3_h
    port map (
            O => \N__5605\,
            I => \N__5602\
        );

    \I__762\ : Span4Mux_v
    port map (
            O => \N__5602\,
            I => \N__5599\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__5599\,
            I => \ADV_R_c_4\
        );

    \I__760\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5593\,
            I => \transmit_module.video_signal_controller.n2076\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__5590\,
            I => \transmit_module.video_signal_controller.n2011_cascade_\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__5587\,
            I => \transmit_module.n1997_cascade_\
        );

    \I__756\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5580\
        );

    \I__755\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5577\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5580\,
            I => \N__5574\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5577\,
            I => \transmit_module.video_signal_controller.n18\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__5574\,
            I => \transmit_module.video_signal_controller.n18\
        );

    \I__751\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5559\
        );

    \I__750\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5559\
        );

    \I__749\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5559\
        );

    \I__748\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5554\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5559\,
            I => \N__5551\
        );

    \I__746\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5548\
        );

    \I__745\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5545\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5554\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__5551\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5548\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5545\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__5536\,
            I => \N__5533\
        );

    \I__739\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5528\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__5532\,
            I => \N__5524\
        );

    \I__737\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5521\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5528\,
            I => \N__5518\
        );

    \I__735\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5513\
        );

    \I__734\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5513\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5521\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__732\ : Odrv4
    port map (
            O => \N__5518\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5513\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__730\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5500\
        );

    \I__729\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5497\
        );

    \I__728\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5494\
        );

    \I__727\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5491\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5500\,
            I => \N__5488\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5497\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5494\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5491\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__5488\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__721\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5473\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__5478\,
            I => \N__5470\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__5477\,
            I => \N__5467\
        );

    \I__718\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5464\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5461\
        );

    \I__716\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5458\
        );

    \I__715\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5455\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5464\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__713\ : Odrv4
    port map (
            O => \N__5461\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5458\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5455\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__710\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5443\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5443\,
            I => \transmit_module.video_signal_controller.n12\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__5440\,
            I => \transmit_module.video_signal_controller.n2146_cascade_\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__5437\,
            I => \transmit_module.video_signal_controller.n1769_cascade_\
        );

    \I__706\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5431\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5431\,
            I => \transmit_module.n2147\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__5428\,
            I => \transmit_module.video_signal_controller.n18_cascade_\
        );

    \I__703\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5422\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5422\,
            I => \transmit_module.video_signal_controller.n8_adj_572\
        );

    \I__701\ : IoInMux
    port map (
            O => \N__5419\,
            I => \N__5416\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5416\,
            I => \N__5413\
        );

    \I__699\ : IoSpan4Mux
    port map (
            O => \N__5413\,
            I => \N__5410\
        );

    \I__698\ : Span4Mux_s3_h
    port map (
            O => \N__5410\,
            I => \N__5407\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__5407\,
            I => \ADV_R_c_5\
        );

    \I__696\ : IoInMux
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5401\,
            I => \N__5398\
        );

    \I__694\ : Span4Mux_s3_h
    port map (
            O => \N__5398\,
            I => \N__5395\
        );

    \I__693\ : Odrv4
    port map (
            O => \N__5395\,
            I => \ADV_R_c_3\
        );

    \I__692\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5389\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5389\,
            I => \transmit_module.Y_DELTA_PATTERN_49\
        );

    \I__690\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5383\,
            I => \transmit_module.Y_DELTA_PATTERN_43\
        );

    \I__688\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__686\ : Odrv4
    port map (
            O => \N__5374\,
            I => \transmit_module.Y_DELTA_PATTERN_42\
        );

    \I__685\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5368\,
            I => \transmit_module.Y_DELTA_PATTERN_52\
        );

    \I__683\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5362\,
            I => \transmit_module.Y_DELTA_PATTERN_51\
        );

    \I__681\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5356\,
            I => \transmit_module.Y_DELTA_PATTERN_50\
        );

    \I__679\ : CEMux
    port map (
            O => \N__5353\,
            I => \N__5346\
        );

    \I__678\ : CEMux
    port map (
            O => \N__5352\,
            I => \N__5343\
        );

    \I__677\ : CEMux
    port map (
            O => \N__5351\,
            I => \N__5338\
        );

    \I__676\ : CEMux
    port map (
            O => \N__5350\,
            I => \N__5335\
        );

    \I__675\ : CEMux
    port map (
            O => \N__5349\,
            I => \N__5331\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5346\,
            I => \N__5328\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5343\,
            I => \N__5325\
        );

    \I__672\ : CEMux
    port map (
            O => \N__5342\,
            I => \N__5322\
        );

    \I__671\ : CEMux
    port map (
            O => \N__5341\,
            I => \N__5319\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__5338\,
            I => \N__5316\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5335\,
            I => \N__5313\
        );

    \I__668\ : CEMux
    port map (
            O => \N__5334\,
            I => \N__5310\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5331\,
            I => \N__5305\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__5328\,
            I => \N__5296\
        );

    \I__665\ : Span4Mux_h
    port map (
            O => \N__5325\,
            I => \N__5296\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5322\,
            I => \N__5296\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5319\,
            I => \N__5296\
        );

    \I__662\ : Span4Mux_v
    port map (
            O => \N__5316\,
            I => \N__5292\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__5313\,
            I => \N__5289\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5286\
        );

    \I__659\ : CEMux
    port map (
            O => \N__5309\,
            I => \N__5283\
        );

    \I__658\ : CEMux
    port map (
            O => \N__5308\,
            I => \N__5280\
        );

    \I__657\ : Span12Mux_h
    port map (
            O => \N__5305\,
            I => \N__5275\
        );

    \I__656\ : Sp12to4
    port map (
            O => \N__5296\,
            I => \N__5275\
        );

    \I__655\ : CEMux
    port map (
            O => \N__5295\,
            I => \N__5272\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__5292\,
            I => \transmit_module.n2159\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__5289\,
            I => \transmit_module.n2159\
        );

    \I__652\ : Odrv12
    port map (
            O => \N__5286\,
            I => \transmit_module.n2159\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__5283\,
            I => \transmit_module.n2159\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5280\,
            I => \transmit_module.n2159\
        );

    \I__649\ : Odrv12
    port map (
            O => \N__5275\,
            I => \transmit_module.n2159\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__5272\,
            I => \transmit_module.n2159\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__5257\,
            I => \transmit_module.video_signal_controller.n2079_cascade_\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__5254\,
            I => \transmit_module.video_signal_controller.n2117_cascade_\
        );

    \I__645\ : InMux
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5248\,
            I => \transmit_module.video_signal_controller.n2154\
        );

    \I__643\ : InMux
    port map (
            O => \N__5245\,
            I => \receive_module.n1822\
        );

    \I__642\ : IoInMux
    port map (
            O => \N__5242\,
            I => \N__5239\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__5239\,
            I => \N__5236\
        );

    \I__640\ : Span4Mux_s3_h
    port map (
            O => \N__5236\,
            I => \N__5232\
        );

    \I__639\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5229\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__5232\,
            I => \DEBUG_c_2\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__5229\,
            I => \DEBUG_c_2\
        );

    \I__636\ : InMux
    port map (
            O => \N__5224\,
            I => \N__5221\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__5221\,
            I => \transmit_module.Y_DELTA_PATTERN_34\
        );

    \I__634\ : InMux
    port map (
            O => \N__5218\,
            I => \N__5215\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5215\,
            I => \transmit_module.Y_DELTA_PATTERN_68\
        );

    \I__632\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5209\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5209\,
            I => \transmit_module.Y_DELTA_PATTERN_67\
        );

    \I__630\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5203\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__5203\,
            I => \transmit_module.Y_DELTA_PATTERN_66\
        );

    \I__628\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5197\,
            I => \transmit_module.Y_DELTA_PATTERN_53\
        );

    \I__626\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5191\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__5191\,
            I => \transmit_module.Y_DELTA_PATTERN_55\
        );

    \I__624\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5185\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5185\,
            I => \transmit_module.Y_DELTA_PATTERN_54\
        );

    \I__622\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5179\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__5179\,
            I => \transmit_module.Y_DELTA_PATTERN_44\
        );

    \I__620\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5173\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5173\,
            I => \receive_module.BRAM_ADDR_5\
        );

    \I__618\ : InMux
    port map (
            O => \N__5170\,
            I => \receive_module.n1814\
        );

    \I__617\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__5164\,
            I => \receive_module.BRAM_ADDR_6\
        );

    \I__615\ : InMux
    port map (
            O => \N__5161\,
            I => \receive_module.n1815\
        );

    \I__614\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5155\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5155\,
            I => \receive_module.BRAM_ADDR_7\
        );

    \I__612\ : InMux
    port map (
            O => \N__5152\,
            I => \receive_module.n1816\
        );

    \I__611\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5146\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__5146\,
            I => \receive_module.BRAM_ADDR_8\
        );

    \I__609\ : InMux
    port map (
            O => \N__5143\,
            I => \bfn_4_8_0_\
        );

    \I__608\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5137\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5137\,
            I => \receive_module.BRAM_ADDR_9\
        );

    \I__606\ : InMux
    port map (
            O => \N__5134\,
            I => \receive_module.n1818\
        );

    \I__605\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5128\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__5128\,
            I => \receive_module.BRAM_ADDR_10\
        );

    \I__603\ : InMux
    port map (
            O => \N__5125\,
            I => \receive_module.n1819\
        );

    \I__602\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__5119\,
            I => \receive_module.BRAM_ADDR_11\
        );

    \I__600\ : InMux
    port map (
            O => \N__5116\,
            I => \receive_module.n1820\
        );

    \I__599\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5110\,
            I => \receive_module.BRAM_ADDR_12\
        );

    \I__597\ : InMux
    port map (
            O => \N__5107\,
            I => \receive_module.n1821\
        );

    \I__596\ : InMux
    port map (
            O => \N__5104\,
            I => \transmit_module.video_signal_controller.n1863\
        );

    \I__595\ : InMux
    port map (
            O => \N__5101\,
            I => \transmit_module.video_signal_controller.n1864\
        );

    \I__594\ : SRMux
    port map (
            O => \N__5098\,
            I => \N__5094\
        );

    \I__593\ : SRMux
    port map (
            O => \N__5097\,
            I => \N__5091\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__5094\,
            I => \N__5088\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__5091\,
            I => \N__5085\
        );

    \I__590\ : Odrv4
    port map (
            O => \N__5088\,
            I => \transmit_module.video_signal_controller.n1582\
        );

    \I__589\ : Odrv12
    port map (
            O => \N__5085\,
            I => \transmit_module.video_signal_controller.n1582\
        );

    \I__588\ : IoInMux
    port map (
            O => \N__5080\,
            I => \N__5077\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__586\ : IoSpan4Mux
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__585\ : Span4Mux_s2_v
    port map (
            O => \N__5071\,
            I => \N__5068\
        );

    \I__584\ : Span4Mux_h
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__583\ : Span4Mux_v
    port map (
            O => \N__5065\,
            I => \N__5062\
        );

    \I__582\ : Odrv4
    port map (
            O => \N__5062\,
            I => \ADV_G_c_6\
        );

    \I__581\ : IoInMux
    port map (
            O => \N__5059\,
            I => \N__5056\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__5056\,
            I => \N__5053\
        );

    \I__579\ : Span4Mux_s1_h
    port map (
            O => \N__5053\,
            I => \N__5050\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__577\ : Odrv4
    port map (
            O => \N__5047\,
            I => \ADV_R_c_1\
        );

    \I__576\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__5041\,
            I => \receive_module.BRAM_ADDR_0\
        );

    \I__574\ : InMux
    port map (
            O => \N__5038\,
            I => \bfn_4_7_0_\
        );

    \I__573\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5032\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__5032\,
            I => \receive_module.BRAM_ADDR_1\
        );

    \I__571\ : InMux
    port map (
            O => \N__5029\,
            I => \receive_module.n1810\
        );

    \I__570\ : InMux
    port map (
            O => \N__5026\,
            I => \N__5023\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__5023\,
            I => \receive_module.BRAM_ADDR_2\
        );

    \I__568\ : InMux
    port map (
            O => \N__5020\,
            I => \receive_module.n1811\
        );

    \I__567\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5014\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__5014\,
            I => \receive_module.BRAM_ADDR_3\
        );

    \I__565\ : InMux
    port map (
            O => \N__5011\,
            I => \receive_module.n1812\
        );

    \I__564\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__5005\,
            I => \receive_module.BRAM_ADDR_4\
        );

    \I__562\ : InMux
    port map (
            O => \N__5002\,
            I => \receive_module.n1813\
        );

    \I__561\ : InMux
    port map (
            O => \N__4999\,
            I => \transmit_module.video_signal_controller.n1854\
        );

    \I__560\ : InMux
    port map (
            O => \N__4996\,
            I => \transmit_module.video_signal_controller.n1855\
        );

    \I__559\ : InMux
    port map (
            O => \N__4993\,
            I => \transmit_module.video_signal_controller.n1856\
        );

    \I__558\ : InMux
    port map (
            O => \N__4990\,
            I => \transmit_module.video_signal_controller.n1857\
        );

    \I__557\ : InMux
    port map (
            O => \N__4987\,
            I => \transmit_module.video_signal_controller.n1858\
        );

    \I__556\ : InMux
    port map (
            O => \N__4984\,
            I => \transmit_module.video_signal_controller.n1859\
        );

    \I__555\ : InMux
    port map (
            O => \N__4981\,
            I => \transmit_module.video_signal_controller.n1860\
        );

    \I__554\ : InMux
    port map (
            O => \N__4978\,
            I => \bfn_3_22_0_\
        );

    \I__553\ : InMux
    port map (
            O => \N__4975\,
            I => \transmit_module.video_signal_controller.n1862\
        );

    \I__552\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4966\
        );

    \I__551\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4966\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4966\,
            I => \transmit_module.video_signal_controller.n1983\
        );

    \I__549\ : CascadeMux
    port map (
            O => \N__4963\,
            I => \transmit_module.video_signal_controller.n2004_cascade_\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__4960\,
            I => \N__4957\
        );

    \I__547\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4954\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4954\,
            I => \transmit_module.video_signal_controller.n9\
        );

    \I__545\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4948\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4948\,
            I => \transmit_module.video_signal_controller.n11\
        );

    \I__543\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4942\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4942\,
            I => \transmit_module.video_signal_controller.n2121\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__4939\,
            I => \transmit_module.video_signal_controller.n7_cascade_\
        );

    \I__540\ : InMux
    port map (
            O => \N__4936\,
            I => \bfn_3_21_0_\
        );

    \I__539\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4930\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4930\,
            I => \transmit_module.Y_DELTA_PATTERN_47\
        );

    \I__537\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4924\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4924\,
            I => \transmit_module.Y_DELTA_PATTERN_46\
        );

    \I__535\ : CEMux
    port map (
            O => \N__4921\,
            I => \N__4918\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4918\,
            I => \N__4914\
        );

    \I__533\ : CEMux
    port map (
            O => \N__4917\,
            I => \N__4911\
        );

    \I__532\ : Span4Mux_v
    port map (
            O => \N__4914\,
            I => \N__4906\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4906\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__4906\,
            I => \N__4903\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__4903\,
            I => \transmit_module.n868\
        );

    \I__528\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4897\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4897\,
            I => \transmit_module.video_signal_controller.SYNC_BUFF1\
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__4894\,
            I => \N__4891\
        );

    \I__525\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4885\
        );

    \I__524\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4885\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4885\,
            I => \N__4882\
        );

    \I__522\ : Span4Mux_v
    port map (
            O => \N__4882\,
            I => \N__4879\
        );

    \I__521\ : Odrv4
    port map (
            O => \N__4879\,
            I => \DEBUG_c_7\
        );

    \I__520\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4867\
        );

    \I__519\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4867\
        );

    \I__518\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4867\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4867\,
            I => \N__4864\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__4864\,
            I => \transmit_module.video_signal_controller.SYNC_BUFF2\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4861\,
            I => \transmit_module.video_signal_controller.n2067_cascade_\
        );

    \I__514\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4855\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4855\,
            I => \transmit_module.video_signal_controller.n4\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__4852\,
            I => \N__4849\
        );

    \I__511\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4845\
        );

    \I__510\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4842\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4845\,
            I => \N__4839\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4842\,
            I => \transmit_module.video_signal_controller.SYNC_EN_SMOOTH\
        );

    \I__507\ : Odrv4
    port map (
            O => \N__4839\,
            I => \transmit_module.video_signal_controller.SYNC_EN_SMOOTH\
        );

    \I__506\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4831\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4831\,
            I => \N__4828\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__4828\,
            I => \transmit_module.Y_DELTA_PATTERN_74\
        );

    \I__503\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4822\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4822\,
            I => \transmit_module.Y_DELTA_PATTERN_73\
        );

    \I__501\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4816\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4816\,
            I => \transmit_module.Y_DELTA_PATTERN_72\
        );

    \I__499\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4810\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4810\,
            I => \transmit_module.Y_DELTA_PATTERN_71\
        );

    \I__497\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4804\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4804\,
            I => \transmit_module.Y_DELTA_PATTERN_45\
        );

    \I__495\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4798\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__493\ : Odrv4
    port map (
            O => \N__4795\,
            I => \transmit_module.Y_DELTA_PATTERN_58\
        );

    \I__492\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4789\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4789\,
            I => \transmit_module.Y_DELTA_PATTERN_57\
        );

    \I__490\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4783\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4783\,
            I => \transmit_module.Y_DELTA_PATTERN_48\
        );

    \I__488\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4777\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4777\,
            I => \transmit_module.Y_DELTA_PATTERN_56\
        );

    \I__486\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4771\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4771\,
            I => \transmit_module.Y_DELTA_PATTERN_76\
        );

    \I__484\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4765\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4765\,
            I => \transmit_module.Y_DELTA_PATTERN_75\
        );

    \I__482\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4759\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4759\,
            I => \transmit_module.Y_DELTA_PATTERN_78\
        );

    \I__480\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4753\,
            I => \transmit_module.Y_DELTA_PATTERN_77\
        );

    \I__478\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4747\,
            I => \transmit_module.Y_DELTA_PATTERN_37\
        );

    \I__476\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4741\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__4741\,
            I => \transmit_module.Y_DELTA_PATTERN_69\
        );

    \I__474\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4735\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4735\,
            I => \transmit_module.Y_DELTA_PATTERN_70\
        );

    \I__472\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4729\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4729\,
            I => \transmit_module.Y_DELTA_PATTERN_36\
        );

    \I__470\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4723\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4723\,
            I => \transmit_module.Y_DELTA_PATTERN_35\
        );

    \I__468\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4717\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4717\,
            I => \transmit_module.Y_DELTA_PATTERN_61\
        );

    \I__466\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4711\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4711\,
            I => \transmit_module.Y_DELTA_PATTERN_65\
        );

    \I__464\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4705\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4705\,
            I => \transmit_module.Y_DELTA_PATTERN_62\
        );

    \I__462\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4699\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4699\,
            I => \transmit_module.Y_DELTA_PATTERN_64\
        );

    \I__460\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4693\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4693\,
            I => \transmit_module.Y_DELTA_PATTERN_63\
        );

    \I__458\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4687\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4687\,
            I => \N__4684\
        );

    \I__456\ : Odrv4
    port map (
            O => \N__4684\,
            I => \transmit_module.Y_DELTA_PATTERN_60\
        );

    \I__455\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4678\,
            I => \transmit_module.Y_DELTA_PATTERN_59\
        );

    \I__453\ : InMux
    port map (
            O => \N__4675\,
            I => \N__4672\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4672\,
            I => \transmit_module.Y_DELTA_PATTERN_97\
        );

    \I__451\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4666\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4666\,
            I => \transmit_module.Y_DELTA_PATTERN_98\
        );

    \I__449\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4660\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4660\,
            I => \transmit_module.Y_DELTA_PATTERN_93\
        );

    \I__447\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4654\,
            I => \transmit_module.Y_DELTA_PATTERN_96\
        );

    \I__445\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4648\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4648\,
            I => \transmit_module.Y_DELTA_PATTERN_95\
        );

    \I__443\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4642\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4642\,
            I => \transmit_module.Y_DELTA_PATTERN_94\
        );

    \I__441\ : IoInMux
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4636\,
            I => \N__4633\
        );

    \I__439\ : Span4Mux_s1_h
    port map (
            O => \N__4633\,
            I => \N__4630\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__4630\,
            I => \ADV_R_c_2\
        );

    \I__437\ : IoInMux
    port map (
            O => \N__4627\,
            I => \N__4624\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4621\
        );

    \I__435\ : IoSpan4Mux
    port map (
            O => \N__4621\,
            I => \N__4618\
        );

    \I__434\ : Span4Mux_s1_h
    port map (
            O => \N__4618\,
            I => \N__4615\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__4615\,
            I => \ADV_R_c_0\
        );

    \I__432\ : IoInMux
    port map (
            O => \N__4612\,
            I => \N__4609\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4609\,
            I => \N__4606\
        );

    \I__430\ : IoSpan4Mux
    port map (
            O => \N__4606\,
            I => \N__4603\
        );

    \I__429\ : Span4Mux_s1_h
    port map (
            O => \N__4603\,
            I => \N__4600\
        );

    \I__428\ : Span4Mux_v
    port map (
            O => \N__4600\,
            I => \N__4597\
        );

    \I__427\ : Odrv4
    port map (
            O => \N__4597\,
            I => \ADV_R_c_6\
        );

    \I__426\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4591\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__4591\,
            I => \transmit_module.Y_DELTA_PATTERN_86\
        );

    \I__424\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4585\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4585\,
            I => \transmit_module.Y_DELTA_PATTERN_90\
        );

    \I__422\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4579\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4579\,
            I => \transmit_module.Y_DELTA_PATTERN_89\
        );

    \I__420\ : InMux
    port map (
            O => \N__4576\,
            I => \N__4573\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4573\,
            I => \transmit_module.Y_DELTA_PATTERN_85\
        );

    \I__418\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4567\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4567\,
            I => \transmit_module.Y_DELTA_PATTERN_88\
        );

    \I__416\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__4561\,
            I => \transmit_module.Y_DELTA_PATTERN_87\
        );

    \I__414\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4555\,
            I => \transmit_module.Y_DELTA_PATTERN_84\
        );

    \I__412\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4549\,
            I => \transmit_module.Y_DELTA_PATTERN_83\
        );

    \I__410\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4543\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4543\,
            I => \transmit_module.Y_DELTA_PATTERN_92\
        );

    \I__408\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__4537\,
            I => \transmit_module.Y_DELTA_PATTERN_91\
        );

    \I__406\ : InMux
    port map (
            O => \N__4534\,
            I => \N__4531\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4531\,
            I => \transmit_module.Y_DELTA_PATTERN_79\
        );

    \I__404\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4525\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4525\,
            I => \transmit_module.Y_DELTA_PATTERN_40\
        );

    \I__402\ : InMux
    port map (
            O => \N__4522\,
            I => \N__4519\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4519\,
            I => \transmit_module.Y_DELTA_PATTERN_39\
        );

    \I__400\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__4513\,
            I => \transmit_module.Y_DELTA_PATTERN_41\
        );

    \I__398\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__4507\,
            I => \transmit_module.Y_DELTA_PATTERN_82\
        );

    \I__396\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4501\,
            I => \transmit_module.Y_DELTA_PATTERN_81\
        );

    \I__394\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__4495\,
            I => \transmit_module.Y_DELTA_PATTERN_80\
        );

    \I__392\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__4489\,
            I => \transmit_module.Y_DELTA_PATTERN_38\
        );

    \I__390\ : IoInMux
    port map (
            O => \N__4486\,
            I => \N__4483\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__388\ : IoSpan4Mux
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__387\ : Span4Mux_s1_v
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__386\ : Sp12to4
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__385\ : Span12Mux_s9_v
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__384\ : Span12Mux_v
    port map (
            O => \N__4468\,
            I => \N__4465\
        );

    \I__383\ : Odrv12
    port map (
            O => \N__4465\,
            I => \CLK_100MHz\
        );

    \INVADV_G__i2C\ : INV
    port map (
            O => \INVADV_G__i2C_net\,
            I => \N__9422\
        );

    \INVADV_G__i3C\ : INV
    port map (
            O => \INVADV_G__i3C_net\,
            I => \N__9519\
        );

    \INVADV_G__i4C\ : INV
    port map (
            O => \INVADV_G__i4C_net\,
            I => \N__9448\
        );

    \INVADV_R__i6C\ : INV
    port map (
            O => \INVADV_R__i6C_net\,
            I => \N__9442\
        );

    \INVADV_G__i7C\ : INV
    port map (
            O => \INVADV_G__i7C_net\,
            I => \N__9450\
        );

    \INVADV_R__i3C\ : INV
    port map (
            O => \INVADV_R__i3C_net\,
            I => \N__9521\
        );

    \IN_MUX_bfv_3_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_21_0_\
        );

    \IN_MUX_bfv_3_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n1861\,
            carryinitout => \bfn_3_22_0_\
        );

    \IN_MUX_bfv_5_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_19_0_\
        );

    \IN_MUX_bfv_5_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n1851\,
            carryinitout => \bfn_5_20_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_5_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.n1830\,
            carryinitout => \bfn_5_16_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n1843\,
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n1877\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_4_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.n1817\,
            carryinitout => \bfn_4_8_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i37_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4492\,
            lcout => \transmit_module.Y_DELTA_PATTERN_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9575\,
            ce => \N__5350\,
            sr => \N__8997\
        );

    \transmit_module.Y_DELTA_PATTERN_i38_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4522\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9575\,
            ce => \N__5350\,
            sr => \N__8997\
        );

    \transmit_module.Y_DELTA_PATTERN_i79_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4498\,
            lcout => \transmit_module.Y_DELTA_PATTERN_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9568\,
            ce => \N__5342\,
            sr => \N__8974\
        );

    \transmit_module.Y_DELTA_PATTERN_i78_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4534\,
            lcout => \transmit_module.Y_DELTA_PATTERN_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9568\,
            ce => \N__5342\,
            sr => \N__8974\
        );

    \transmit_module.Y_DELTA_PATTERN_i40_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4516\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9568\,
            ce => \N__5342\,
            sr => \N__8974\
        );

    \transmit_module.Y_DELTA_PATTERN_i39_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4528\,
            lcout => \transmit_module.Y_DELTA_PATTERN_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9568\,
            ce => \N__5342\,
            sr => \N__8974\
        );

    \transmit_module.Y_DELTA_PATTERN_i41_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5380\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9566\,
            ce => \N__5308\,
            sr => \N__8933\
        );

    \transmit_module.Y_DELTA_PATTERN_i81_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4510\,
            lcout => \transmit_module.Y_DELTA_PATTERN_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9566\,
            ce => \N__5308\,
            sr => \N__8933\
        );

    \transmit_module.Y_DELTA_PATTERN_i82_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4552\,
            lcout => \transmit_module.Y_DELTA_PATTERN_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9566\,
            ce => \N__5308\,
            sr => \N__8933\
        );

    \transmit_module.Y_DELTA_PATTERN_i80_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4504\,
            lcout => \transmit_module.Y_DELTA_PATTERN_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9566\,
            ce => \N__5308\,
            sr => \N__8933\
        );

    \transmit_module.Y_DELTA_PATTERN_i88_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4582\,
            lcout => \transmit_module.Y_DELTA_PATTERN_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => \N__4917\,
            sr => \N__8908\
        );

    \transmit_module.Y_DELTA_PATTERN_i85_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4594\,
            lcout => \transmit_module.Y_DELTA_PATTERN_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => \N__4917\,
            sr => \N__8908\
        );

    \transmit_module.Y_DELTA_PATTERN_i90_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4540\,
            lcout => \transmit_module.Y_DELTA_PATTERN_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => \N__4917\,
            sr => \N__8908\
        );

    \transmit_module.Y_DELTA_PATTERN_i86_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4564\,
            lcout => \transmit_module.Y_DELTA_PATTERN_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => \N__4917\,
            sr => \N__8908\
        );

    \transmit_module.Y_DELTA_PATTERN_i89_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4588\,
            lcout => \transmit_module.Y_DELTA_PATTERN_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => \N__4917\,
            sr => \N__8908\
        );

    \transmit_module.Y_DELTA_PATTERN_i84_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4576\,
            lcout => \transmit_module.Y_DELTA_PATTERN_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => \N__4917\,
            sr => \N__8908\
        );

    \transmit_module.Y_DELTA_PATTERN_i87_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4570\,
            lcout => \transmit_module.Y_DELTA_PATTERN_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => \N__4917\,
            sr => \N__8908\
        );

    \transmit_module.Y_DELTA_PATTERN_i83_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4558\,
            lcout => \transmit_module.Y_DELTA_PATTERN_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => \N__4917\,
            sr => \N__8908\
        );

    \transmit_module.Y_DELTA_PATTERN_i96_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4675\,
            lcout => \transmit_module.Y_DELTA_PATTERN_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => \N__4921\,
            sr => \N__8924\
        );

    \transmit_module.Y_DELTA_PATTERN_i92_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4663\,
            lcout => \transmit_module.Y_DELTA_PATTERN_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => \N__4921\,
            sr => \N__8924\
        );

    \transmit_module.Y_DELTA_PATTERN_i91_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4546\,
            lcout => \transmit_module.Y_DELTA_PATTERN_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => \N__4921\,
            sr => \N__8924\
        );

    \transmit_module.Y_DELTA_PATTERN_i97_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4669\,
            lcout => \transmit_module.Y_DELTA_PATTERN_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => \N__4921\,
            sr => \N__8924\
        );

    \transmit_module.Y_DELTA_PATTERN_i98_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6850\,
            lcout => \transmit_module.Y_DELTA_PATTERN_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => \N__4921\,
            sr => \N__8924\
        );

    \transmit_module.Y_DELTA_PATTERN_i93_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4645\,
            lcout => \transmit_module.Y_DELTA_PATTERN_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => \N__4921\,
            sr => \N__8924\
        );

    \transmit_module.Y_DELTA_PATTERN_i95_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4657\,
            lcout => \transmit_module.Y_DELTA_PATTERN_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => \N__4921\,
            sr => \N__8924\
        );

    \transmit_module.Y_DELTA_PATTERN_i94_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4651\,
            lcout => \transmit_module.Y_DELTA_PATTERN_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => \N__4921\,
            sr => \N__8924\
        );

    \ADV_R__i3_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6966\,
            lcout => \ADV_R_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i3C_net\,
            ce => 'H',
            sr => \N__6907\
        );

    \ADV_R__i1_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6597\,
            lcout => \ADV_R_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i3C_net\,
            ce => 'H',
            sr => \N__6907\
        );

    \ADV_R__i7_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7105\,
            lcout => \ADV_R_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i3C_net\,
            ce => 'H',
            sr => \N__6907\
        );

    \transmit_module.Y_DELTA_PATTERN_i60_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4720\,
            lcout => \transmit_module.Y_DELTA_PATTERN_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9446\,
            ce => \N__5353\,
            sr => \N__8981\
        );

    \transmit_module.Y_DELTA_PATTERN_i74_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4768\,
            lcout => \transmit_module.Y_DELTA_PATTERN_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9584\,
            ce => \N__5352\,
            sr => \N__8989\
        );

    \transmit_module.Y_DELTA_PATTERN_i61_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4708\,
            lcout => \transmit_module.Y_DELTA_PATTERN_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9584\,
            ce => \N__5352\,
            sr => \N__8989\
        );

    \transmit_module.Y_DELTA_PATTERN_i64_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4714\,
            lcout => \transmit_module.Y_DELTA_PATTERN_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9584\,
            ce => \N__5352\,
            sr => \N__8989\
        );

    \transmit_module.Y_DELTA_PATTERN_i65_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5206\,
            lcout => \transmit_module.Y_DELTA_PATTERN_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9584\,
            ce => \N__5352\,
            sr => \N__8989\
        );

    \transmit_module.Y_DELTA_PATTERN_i62_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4696\,
            lcout => \transmit_module.Y_DELTA_PATTERN_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9584\,
            ce => \N__5352\,
            sr => \N__8989\
        );

    \transmit_module.Y_DELTA_PATTERN_i63_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4702\,
            lcout => \transmit_module.Y_DELTA_PATTERN_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9584\,
            ce => \N__5352\,
            sr => \N__8989\
        );

    \transmit_module.Y_DELTA_PATTERN_i58_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4681\,
            lcout => \transmit_module.Y_DELTA_PATTERN_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => \N__5334\,
            sr => \N__8909\
        );

    \transmit_module.Y_DELTA_PATTERN_i34_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4726\,
            lcout => \transmit_module.Y_DELTA_PATTERN_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => \N__5334\,
            sr => \N__8909\
        );

    \transmit_module.Y_DELTA_PATTERN_i59_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4690\,
            lcout => \transmit_module.Y_DELTA_PATTERN_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => \N__5334\,
            sr => \N__8909\
        );

    \transmit_module.Y_DELTA_PATTERN_i76_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4756\,
            lcout => \transmit_module.Y_DELTA_PATTERN_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => \N__5334\,
            sr => \N__8909\
        );

    \transmit_module.Y_DELTA_PATTERN_i68_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4744\,
            lcout => \transmit_module.Y_DELTA_PATTERN_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => \N__5334\,
            sr => \N__8909\
        );

    \transmit_module.Y_DELTA_PATTERN_i75_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4774\,
            lcout => \transmit_module.Y_DELTA_PATTERN_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => \N__5334\,
            sr => \N__8909\
        );

    \transmit_module.Y_DELTA_PATTERN_i77_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4762\,
            lcout => \transmit_module.Y_DELTA_PATTERN_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => \N__5334\,
            sr => \N__8909\
        );

    \transmit_module.Y_DELTA_PATTERN_i36_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4750\,
            lcout => \transmit_module.Y_DELTA_PATTERN_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => \N__5334\,
            sr => \N__8909\
        );

    \transmit_module.Y_DELTA_PATTERN_i69_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4738\,
            lcout => \transmit_module.Y_DELTA_PATTERN_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9355\,
            ce => \N__5341\,
            sr => \N__8925\
        );

    \transmit_module.Y_DELTA_PATTERN_i70_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4813\,
            lcout => \transmit_module.Y_DELTA_PATTERN_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9355\,
            ce => \N__5341\,
            sr => \N__8925\
        );

    \transmit_module.Y_DELTA_PATTERN_i72_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4825\,
            lcout => \transmit_module.Y_DELTA_PATTERN_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9355\,
            ce => \N__5341\,
            sr => \N__8925\
        );

    \transmit_module.Y_DELTA_PATTERN_i35_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4732\,
            lcout => \transmit_module.Y_DELTA_PATTERN_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9355\,
            ce => \N__5341\,
            sr => \N__8925\
        );

    \transmit_module.Y_DELTA_PATTERN_i73_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4834\,
            lcout => \transmit_module.Y_DELTA_PATTERN_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9355\,
            ce => \N__5341\,
            sr => \N__8925\
        );

    \transmit_module.Y_DELTA_PATTERN_i71_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4819\,
            lcout => \transmit_module.Y_DELTA_PATTERN_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9355\,
            ce => \N__5341\,
            sr => \N__8925\
        );

    \transmit_module.Y_DELTA_PATTERN_i45_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4927\,
            lcout => \transmit_module.Y_DELTA_PATTERN_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9356\,
            ce => \N__5295\,
            sr => \N__8842\
        );

    \transmit_module.Y_DELTA_PATTERN_i44_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4807\,
            lcout => \transmit_module.Y_DELTA_PATTERN_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9356\,
            ce => \N__5295\,
            sr => \N__8842\
        );

    \transmit_module.Y_DELTA_PATTERN_i48_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5392\,
            lcout => \transmit_module.Y_DELTA_PATTERN_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9356\,
            ce => \N__5295\,
            sr => \N__8842\
        );

    \transmit_module.Y_DELTA_PATTERN_i56_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4792\,
            lcout => \transmit_module.Y_DELTA_PATTERN_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9356\,
            ce => \N__5295\,
            sr => \N__8842\
        );

    \transmit_module.Y_DELTA_PATTERN_i57_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4801\,
            lcout => \transmit_module.Y_DELTA_PATTERN_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9356\,
            ce => \N__5295\,
            sr => \N__8842\
        );

    \transmit_module.Y_DELTA_PATTERN_i47_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4786\,
            lcout => \transmit_module.Y_DELTA_PATTERN_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9356\,
            ce => \N__5295\,
            sr => \N__8842\
        );

    \transmit_module.Y_DELTA_PATTERN_i55_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4780\,
            lcout => \transmit_module.Y_DELTA_PATTERN_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9356\,
            ce => \N__5295\,
            sr => \N__8842\
        );

    \transmit_module.Y_DELTA_PATTERN_i46_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4933\,
            lcout => \transmit_module.Y_DELTA_PATTERN_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9356\,
            ce => \N__5295\,
            sr => \N__8842\
        );

    \transmit_module.video_signal_controller.i280_2_lut_3_lut_4_lut_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__8407\,
            in1 => \N__6219\,
            in2 => \N__8972\,
            in3 => \N__6187\,
            lcout => \transmit_module.n868\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i280_2_lut_3_lut_4_lut_rep_23_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__8408\,
            in1 => \N__6220\,
            in2 => \N__8973\,
            in3 => \N__6186\,
            lcout => \transmit_module.n2159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.SYNC_BUFF1_57_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5928\,
            lcout => \transmit_module.video_signal_controller.SYNC_BUFF1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9354\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.SYNC_BUFF2_58_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4900\,
            lcout => \transmit_module.video_signal_controller.SYNC_BUFF2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9354\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i2_4_lut_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__8549\,
            in1 => \N__5434\,
            in2 => \N__8827\,
            in3 => \N__8406\,
            lcout => \transmit_module.n694\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__6735\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4890\,
            lcout => \transmit_module.video_signal_controller.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_16_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__4875\,
            in1 => \N__6736\,
            in2 => \N__4852\,
            in3 => \N__4972\,
            lcout => \transmit_module.video_signal_controller.n1582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i3_4_lut_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4874\,
            in1 => \N__6734\,
            in2 => \N__4894\,
            in3 => \N__4971\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2067_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.SYNC_EN_SMOOTH_64_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110010"
        )
    port map (
            in0 => \N__4848\,
            in1 => \N__4876\,
            in2 => \N__4861\,
            in3 => \N__4858\,
            lcout => \transmit_module.video_signal_controller.SYNC_EN_SMOOTH\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i6_4_lut_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4951\,
            in1 => \N__6480\,
            in2 => \N__4960\,
            in3 => \N__6663\,
            lcout => \transmit_module.video_signal_controller.n1983\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1958_2_lut_4_lut_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5782\,
            in1 => \N__6971\,
            in2 => \N__7110\,
            in3 => \N__5569\,
            lcout => \transmit_module.video_signal_controller.n2121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_4_lut_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__7097\,
            in1 => \N__5780\,
            in2 => \N__5536\,
            in3 => \N__7024\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2004_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_adj_12_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__5479\,
            in1 => \N__5506\,
            in2 => \N__4963\,
            in3 => \N__5567\,
            lcout => \transmit_module.video_signal_controller.n2076\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_adj_15_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5568\,
            in1 => \N__6965\,
            in2 => \_gnd_net_\,
            in3 => \N__5703\,
            lcout => \transmit_module.video_signal_controller.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i4_4_lut_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5781\,
            in1 => \N__5811\,
            in2 => \N__6603\,
            in3 => \N__7098\,
            lcout => \transmit_module.video_signal_controller.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_3_lut_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__6602\,
            in1 => \N__6481\,
            in2 => \_gnd_net_\,
            in3 => \N__6664\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VS_61_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5704\,
            in1 => \N__4945\,
            in2 => \N__4939\,
            in3 => \N__5812\,
            lcout => \ADV_VSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i0_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6598\,
            in2 => \_gnd_net_\,
            in3 => \N__4936\,
            lcout => \VGA_Y_0\,
            ltout => OPEN,
            carryin => \bfn_3_21_0_\,
            carryout => \transmit_module.video_signal_controller.n1854\,
            clk => \N__9520\,
            ce => \N__6762\,
            sr => \N__5097\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i1_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6485\,
            in2 => \_gnd_net_\,
            in3 => \N__4999\,
            lcout => \VGA_Y_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1854\,
            carryout => \transmit_module.video_signal_controller.n1855\,
            clk => \N__9520\,
            ce => \N__6762\,
            sr => \N__5097\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i2_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6967\,
            in2 => \_gnd_net_\,
            in3 => \N__4996\,
            lcout => \VGA_Y_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1855\,
            carryout => \transmit_module.video_signal_controller.n1856\,
            clk => \N__9520\,
            ce => \N__6762\,
            sr => \N__5097\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i3_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5709\,
            in2 => \_gnd_net_\,
            in3 => \N__4993\,
            lcout => \VGA_Y_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1856\,
            carryout => \transmit_module.video_signal_controller.n1857\,
            clk => \N__9520\,
            ce => \N__6762\,
            sr => \N__5097\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i4_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6669\,
            in2 => \_gnd_net_\,
            in3 => \N__4990\,
            lcout => \VGA_Y_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1857\,
            carryout => \transmit_module.video_signal_controller.n1858\,
            clk => \N__9520\,
            ce => \N__6762\,
            sr => \N__5097\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i5_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5785\,
            in2 => \_gnd_net_\,
            in3 => \N__4987\,
            lcout => \VGA_Y_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1858\,
            carryout => \transmit_module.video_signal_controller.n1859\,
            clk => \N__9520\,
            ce => \N__6762\,
            sr => \N__5097\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i6_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7106\,
            in2 => \_gnd_net_\,
            in3 => \N__4984\,
            lcout => \VGA_Y_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1859\,
            carryout => \transmit_module.video_signal_controller.n1860\,
            clk => \N__9520\,
            ce => \N__6762\,
            sr => \N__5097\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i7_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7031\,
            in2 => \_gnd_net_\,
            in3 => \N__4981\,
            lcout => \VGA_Y_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1860\,
            carryout => \transmit_module.video_signal_controller.n1861\,
            clk => \N__9520\,
            ce => \N__6762\,
            sr => \N__5097\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i8_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5531\,
            in2 => \_gnd_net_\,
            in3 => \N__4978\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_8\,
            ltout => OPEN,
            carryin => \bfn_3_22_0_\,
            carryout => \transmit_module.video_signal_controller.n1862\,
            clk => \N__9495\,
            ce => \N__6763\,
            sr => \N__5098\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i9_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5566\,
            in2 => \_gnd_net_\,
            in3 => \N__4975\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1862\,
            carryout => \transmit_module.video_signal_controller.n1863\,
            clk => \N__9495\,
            ce => \N__6763\,
            sr => \N__5098\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i10_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5476\,
            in2 => \_gnd_net_\,
            in3 => \N__5104\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1863\,
            carryout => \transmit_module.video_signal_controller.n1864\,
            clk => \N__9495\,
            ce => \N__6763\,
            sr => \N__5098\
        );

    \transmit_module.video_signal_controller.VGA_Y_274__i11_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5505\,
            in2 => \_gnd_net_\,
            in3 => \N__5101\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9495\,
            ce => \N__6763\,
            sr => \N__5098\
        );

    \ADV_G__i7_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6367\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ADV_G_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i7C_net\,
            ce => 'H',
            sr => \N__6906\
        );

    \ADV_R__i2_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6489\,
            lcout => \ADV_R_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i7C_net\,
            ce => 'H',
            sr => \N__6906\
        );

    \receive_module.BRAM_ADDR__i0_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5044\,
            in2 => \_gnd_net_\,
            in3 => \N__5038\,
            lcout => \receive_module.BRAM_ADDR_0\,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => \receive_module.n1810\,
            clk => \N__9863\,
            ce => \N__5878\,
            sr => \N__8636\
        );

    \receive_module.BRAM_ADDR__i1_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5035\,
            in2 => \_gnd_net_\,
            in3 => \N__5029\,
            lcout => \receive_module.BRAM_ADDR_1\,
            ltout => OPEN,
            carryin => \receive_module.n1810\,
            carryout => \receive_module.n1811\,
            clk => \N__9863\,
            ce => \N__5878\,
            sr => \N__8636\
        );

    \receive_module.BRAM_ADDR__i2_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5026\,
            in2 => \_gnd_net_\,
            in3 => \N__5020\,
            lcout => \receive_module.BRAM_ADDR_2\,
            ltout => OPEN,
            carryin => \receive_module.n1811\,
            carryout => \receive_module.n1812\,
            clk => \N__9863\,
            ce => \N__5878\,
            sr => \N__8636\
        );

    \receive_module.BRAM_ADDR__i3_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5017\,
            in2 => \_gnd_net_\,
            in3 => \N__5011\,
            lcout => \receive_module.BRAM_ADDR_3\,
            ltout => OPEN,
            carryin => \receive_module.n1812\,
            carryout => \receive_module.n1813\,
            clk => \N__9863\,
            ce => \N__5878\,
            sr => \N__8636\
        );

    \receive_module.BRAM_ADDR__i4_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5008\,
            in2 => \_gnd_net_\,
            in3 => \N__5002\,
            lcout => \receive_module.BRAM_ADDR_4\,
            ltout => OPEN,
            carryin => \receive_module.n1813\,
            carryout => \receive_module.n1814\,
            clk => \N__9863\,
            ce => \N__5878\,
            sr => \N__8636\
        );

    \receive_module.BRAM_ADDR__i5_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5176\,
            in2 => \_gnd_net_\,
            in3 => \N__5170\,
            lcout => \receive_module.BRAM_ADDR_5\,
            ltout => OPEN,
            carryin => \receive_module.n1814\,
            carryout => \receive_module.n1815\,
            clk => \N__9863\,
            ce => \N__5878\,
            sr => \N__8636\
        );

    \receive_module.BRAM_ADDR__i6_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5167\,
            in2 => \_gnd_net_\,
            in3 => \N__5161\,
            lcout => \receive_module.BRAM_ADDR_6\,
            ltout => OPEN,
            carryin => \receive_module.n1815\,
            carryout => \receive_module.n1816\,
            clk => \N__9863\,
            ce => \N__5878\,
            sr => \N__8636\
        );

    \receive_module.BRAM_ADDR__i7_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5158\,
            in2 => \_gnd_net_\,
            in3 => \N__5152\,
            lcout => \receive_module.BRAM_ADDR_7\,
            ltout => OPEN,
            carryin => \receive_module.n1816\,
            carryout => \receive_module.n1817\,
            clk => \N__9863\,
            ce => \N__5878\,
            sr => \N__8636\
        );

    \receive_module.BRAM_ADDR__i8_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5149\,
            in2 => \_gnd_net_\,
            in3 => \N__5143\,
            lcout => \receive_module.BRAM_ADDR_8\,
            ltout => OPEN,
            carryin => \bfn_4_8_0_\,
            carryout => \receive_module.n1818\,
            clk => \N__9865\,
            ce => \N__5874\,
            sr => \N__8644\
        );

    \receive_module.BRAM_ADDR__i9_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5140\,
            in2 => \_gnd_net_\,
            in3 => \N__5134\,
            lcout => \receive_module.BRAM_ADDR_9\,
            ltout => OPEN,
            carryin => \receive_module.n1818\,
            carryout => \receive_module.n1819\,
            clk => \N__9865\,
            ce => \N__5874\,
            sr => \N__8644\
        );

    \receive_module.BRAM_ADDR__i10_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5131\,
            in2 => \_gnd_net_\,
            in3 => \N__5125\,
            lcout => \receive_module.BRAM_ADDR_10\,
            ltout => OPEN,
            carryin => \receive_module.n1819\,
            carryout => \receive_module.n1820\,
            clk => \N__9865\,
            ce => \N__5874\,
            sr => \N__8644\
        );

    \receive_module.BRAM_ADDR__i11_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5122\,
            in2 => \_gnd_net_\,
            in3 => \N__5116\,
            lcout => \receive_module.BRAM_ADDR_11\,
            ltout => OPEN,
            carryin => \receive_module.n1820\,
            carryout => \receive_module.n1821\,
            clk => \N__9865\,
            ce => \N__5874\,
            sr => \N__8644\
        );

    \receive_module.BRAM_ADDR__i12_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5113\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => \receive_module.BRAM_ADDR_12\,
            ltout => OPEN,
            carryin => \receive_module.n1821\,
            carryout => \receive_module.n1822\,
            clk => \N__9865\,
            ce => \N__5874\,
            sr => \N__8644\
        );

    \receive_module.BRAM_ADDR__i13_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5235\,
            in2 => \_gnd_net_\,
            in3 => \N__5245\,
            lcout => \DEBUG_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9865\,
            ce => \N__5874\,
            sr => \N__8644\
        );

    \transmit_module.ADDR_Y_COMPONENT__i4_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6106\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9586\,
            ce => \N__7651\,
            sr => \N__8976\
        );

    \transmit_module.Y_DELTA_PATTERN_i33_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5224\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9221\,
            ce => \N__5351\,
            sr => \N__8980\
        );

    \transmit_module.Y_DELTA_PATTERN_i67_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5218\,
            lcout => \transmit_module.Y_DELTA_PATTERN_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9221\,
            ce => \N__5351\,
            sr => \N__8980\
        );

    \transmit_module.Y_DELTA_PATTERN_i66_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5212\,
            lcout => \transmit_module.Y_DELTA_PATTERN_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9221\,
            ce => \N__5351\,
            sr => \N__8980\
        );

    \transmit_module.Y_DELTA_PATTERN_i53_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5188\,
            lcout => \transmit_module.Y_DELTA_PATTERN_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9550\,
            ce => \N__5349\,
            sr => \N__8926\
        );

    \transmit_module.Y_DELTA_PATTERN_i52_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5200\,
            lcout => \transmit_module.Y_DELTA_PATTERN_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9550\,
            ce => \N__5349\,
            sr => \N__8926\
        );

    \transmit_module.Y_DELTA_PATTERN_i54_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5194\,
            lcout => \transmit_module.Y_DELTA_PATTERN_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9550\,
            ce => \N__5349\,
            sr => \N__8926\
        );

    \transmit_module.Y_DELTA_PATTERN_i43_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5182\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9577\,
            ce => \N__5309\,
            sr => \N__8943\
        );

    \transmit_module.Y_DELTA_PATTERN_i49_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5359\,
            lcout => \transmit_module.Y_DELTA_PATTERN_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9577\,
            ce => \N__5309\,
            sr => \N__8943\
        );

    \transmit_module.Y_DELTA_PATTERN_i42_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5386\,
            lcout => \transmit_module.Y_DELTA_PATTERN_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9577\,
            ce => \N__5309\,
            sr => \N__8943\
        );

    \transmit_module.Y_DELTA_PATTERN_i51_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5371\,
            lcout => \transmit_module.Y_DELTA_PATTERN_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9577\,
            ce => \N__5309\,
            sr => \N__8943\
        );

    \transmit_module.Y_DELTA_PATTERN_i50_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5365\,
            lcout => \transmit_module.Y_DELTA_PATTERN_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9577\,
            ce => \N__5309\,
            sr => \N__8943\
        );

    \transmit_module.video_signal_controller.i2_3_lut_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6550\,
            in1 => \N__7157\,
            in2 => \_gnd_net_\,
            in3 => \N__6362\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2079_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1954_4_lut_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__7260\,
            in1 => \N__6796\,
            in2 => \N__5257\,
            in3 => \N__6835\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_HS_60_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__5446\,
            in1 => \N__5251\,
            in2 => \N__5254\,
            in3 => \N__6325\,
            lcout => \ADV_HSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i433_2_lut_rep_18_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7259\,
            in2 => \_gnd_net_\,
            in3 => \N__6361\,
            lcout => \transmit_module.video_signal_controller.n2154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.old_VGA_HS_34_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6188\,
            lcout => \transmit_module.old_VGA_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i319_3_lut_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7158\,
            in1 => \N__6551\,
            in2 => \_gnd_net_\,
            in3 => \N__6402\,
            lcout => \transmit_module.video_signal_controller.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_10_3_lut_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7166\,
            in1 => \N__7254\,
            in2 => \_gnd_net_\,
            in3 => \N__6354\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1677_4_lut_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6431\,
            in1 => \N__6549\,
            in2 => \N__5440\,
            in3 => \N__5425\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n1769_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1690_4_lut_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__6829\,
            in1 => \N__6324\,
            in2 => \N__5437\,
            in3 => \N__6790\,
            lcout => \transmit_module.video_signal_controller.n528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_3_lut_rep_11_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__6789\,
            in1 => \N__6828\,
            in2 => \_gnd_net_\,
            in3 => \N__5583\,
            lcout => \transmit_module.n2147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i357_2_lut_3_lut_4_lut_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__6323\,
            in1 => \N__7253\,
            in2 => \N__7168\,
            in3 => \N__6353\,
            lcout => \transmit_module.video_signal_controller.n18\,
            ltout => \transmit_module.video_signal_controller.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_8_4_lut_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011000000000"
        )
    port map (
            in0 => \N__6791\,
            in1 => \N__6830\,
            in2 => \N__5428\,
            in3 => \N__8384\,
            lcout => n2144,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i3_3_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6704\,
            in1 => \N__6397\,
            in2 => \_gnd_net_\,
            in3 => \N__7202\,
            lcout => \transmit_module.video_signal_controller.n8_adj_572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADV_R__i6_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5783\,
            lcout => \ADV_R_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i6C_net\,
            ce => 'H',
            sr => \N__6881\
        );

    \ADV_R__i4_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5705\,
            lcout => \ADV_R_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i6C_net\,
            ce => 'H',
            sr => \N__6881\
        );

    \ADV_B__i6_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5784\,
            lcout => \ADV_B_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i6C_net\,
            ce => 'H',
            sr => \N__6881\
        );

    \ADV_G__i1_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6432\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ADV_G_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i6C_net\,
            ce => 'H',
            sr => \N__6881\
        );

    \ADV_R__i5_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6665\,
            lcout => \ADV_R_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i6C_net\,
            ce => 'H',
            sr => \N__6881\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_13_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__5504\,
            in1 => \N__5558\,
            in2 => \N__5478\,
            in3 => \N__5740\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2011_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_10_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100000000"
        )
    port map (
            in0 => \N__5596\,
            in1 => \N__6662\,
            in2 => \N__5590\,
            in3 => \N__5791\,
            lcout => \transmit_module.n1997\,
            ltout => \transmit_module.n1997_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1055_1_lut_2_lut_4_lut_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110011111"
        )
    port map (
            in0 => \N__6827\,
            in1 => \N__6788\,
            in2 => \N__5587\,
            in3 => \N__5584\,
            lcout => n1144,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_16_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5532\,
            in3 => \N__7022\,
            lcout => \transmit_module.video_signal_controller.n2152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_rep_15_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5779\,
            in1 => \N__5557\,
            in2 => \_gnd_net_\,
            in3 => \N__7095\,
            lcout => \transmit_module.video_signal_controller.n2151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_3_lut_4_lut_adj_14_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5527\,
            in1 => \N__5503\,
            in2 => \N__5477\,
            in3 => \N__7023\,
            lcout => \transmit_module.video_signal_controller.n679\,
            ltout => \transmit_module.video_signal_controller.n679_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6661\,
            in1 => \N__5734\,
            in2 => \N__5800\,
            in3 => \N__5797\,
            lcout => \transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_13_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5778\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_11_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__6479\,
            in1 => \N__5728\,
            in2 => \N__5749\,
            in3 => \N__5746\,
            lcout => \transmit_module.video_signal_controller.n2006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i335_3_lut_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__5702\,
            in1 => \N__6478\,
            in2 => \_gnd_net_\,
            in3 => \N__6964\,
            lcout => \transmit_module.video_signal_controller.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_rep_4_2_lut_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6972\,
            in3 => \N__5701\,
            lcout => \transmit_module.video_signal_controller.n2140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADV_G__i4_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6406\,
            lcout => \ADV_G_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i4C_net\,
            ce => 'H',
            sr => \N__6905\
        );

    \ADV_B__i4_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5710\,
            lcout => \ADV_B_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i4C_net\,
            ce => 'H',
            sr => \N__6905\
        );

    \receive_module.rx_counter.i26_1_lut_rep_19_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9939\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.n2155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.SYNC_45_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7267\,
            in1 => \N__7282\,
            in2 => \N__7294\,
            in3 => \N__7996\,
            lcout => \DEBUG_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i35_4_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010111001"
        )
    port map (
            in0 => \N__5956\,
            in1 => \N__5980\,
            in2 => \N__5857\,
            in3 => \N__5848\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1973_4_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__8029\,
            in1 => \N__7273\,
            in2 => \N__5902\,
            in3 => \N__7393\,
            lcout => \DEBUG_c_4\,
            ltout => \DEBUG_c_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i1969_2_lut_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5881\,
            in3 => \N__9940\,
            lcout => \receive_module.n788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_adj_19_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6000\,
            in1 => \N__6021\,
            in2 => \_gnd_net_\,
            in3 => \N__5838\,
            lcout => \receive_module.rx_counter.n2083\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1871_3_lut_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__6022\,
            in1 => \_gnd_net_\,
            in2 => \N__5842\,
            in3 => \N__6001\,
            lcout => \receive_module.rx_counter.n2033\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__6051\,
            in2 => \_gnd_net_\,
            in3 => \N__6066\,
            lcout => \receive_module.rx_counter.n1981\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.X_272__i0_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5830\,
            in2 => \_gnd_net_\,
            in3 => \N__5824\,
            lcout => \receive_module.rx_counter.n10\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \receive_module.rx_counter.n1870\,
            clk => \N__9866\,
            ce => 'H',
            sr => \N__7386\
        );

    \receive_module.rx_counter.X_272__i1_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5821\,
            in2 => \_gnd_net_\,
            in3 => \N__5815\,
            lcout => \receive_module.rx_counter.n9\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1870\,
            carryout => \receive_module.rx_counter.n1871\,
            clk => \N__9866\,
            ce => 'H',
            sr => \N__7386\
        );

    \receive_module.rx_counter.X_272__i2_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6076\,
            in2 => \_gnd_net_\,
            in3 => \N__6070\,
            lcout => \receive_module.rx_counter.n8_adj_575\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1871\,
            carryout => \receive_module.rx_counter.n1872\,
            clk => \N__9866\,
            ce => 'H',
            sr => \N__7386\
        );

    \receive_module.rx_counter.X_272__i3_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6067\,
            in2 => \_gnd_net_\,
            in3 => \N__6055\,
            lcout => \receive_module.rx_counter.X_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1872\,
            carryout => \receive_module.rx_counter.n1873\,
            clk => \N__9866\,
            ce => 'H',
            sr => \N__7386\
        );

    \receive_module.rx_counter.X_272__i4_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6052\,
            in2 => \_gnd_net_\,
            in3 => \N__6040\,
            lcout => \receive_module.rx_counter.X_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1873\,
            carryout => \receive_module.rx_counter.n1874\,
            clk => \N__9866\,
            ce => 'H',
            sr => \N__7386\
        );

    \receive_module.rx_counter.X_272__i5_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6037\,
            in2 => \_gnd_net_\,
            in3 => \N__6025\,
            lcout => \receive_module.rx_counter.X_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1874\,
            carryout => \receive_module.rx_counter.n1875\,
            clk => \N__9866\,
            ce => 'H',
            sr => \N__7386\
        );

    \receive_module.rx_counter.X_272__i6_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6020\,
            in2 => \_gnd_net_\,
            in3 => \N__6004\,
            lcout => \receive_module.rx_counter.X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1875\,
            carryout => \receive_module.rx_counter.n1876\,
            clk => \N__9866\,
            ce => 'H',
            sr => \N__7386\
        );

    \receive_module.rx_counter.X_272__i7_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5999\,
            in2 => \_gnd_net_\,
            in3 => \N__5983\,
            lcout => \receive_module.rx_counter.X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1876\,
            carryout => \receive_module.rx_counter.n1877\,
            clk => \N__9866\,
            ce => 'H',
            sr => \N__7386\
        );

    \receive_module.rx_counter.X_272__i8_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5976\,
            in2 => \_gnd_net_\,
            in3 => \N__5962\,
            lcout => \receive_module.rx_counter.X_8\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \receive_module.rx_counter.n1878\,
            clk => \N__9867\,
            ce => 'H',
            sr => \N__7387\
        );

    \receive_module.rx_counter.X_272__i9_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5955\,
            in2 => \_gnd_net_\,
            in3 => \N__5959\,
            lcout => \receive_module.rx_counter.X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9867\,
            ce => 'H',
            sr => \N__7387\
        );

    \transmit_module.BRAM_ADDR__i4_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__6094\,
            in1 => \N__8547\,
            in2 => \N__5941\,
            in3 => \N__8431\,
            lcout => \transmit_module.BRAM_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9585\,
            ce => \N__8315\,
            sr => \N__8996\
        );

    \transmit_module.add_13_2_lut_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7453\,
            in2 => \N__7576\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n204\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \transmit_module.n1823\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_3_lut_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7554\,
            in2 => \_gnd_net_\,
            in3 => \N__6115\,
            lcout => \transmit_module.n203\,
            ltout => OPEN,
            carryin => \transmit_module.n1823\,
            carryout => \transmit_module.n1824\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_4_lut_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7675\,
            in2 => \_gnd_net_\,
            in3 => \N__6112\,
            lcout => \transmit_module.n202\,
            ltout => OPEN,
            carryin => \transmit_module.n1824\,
            carryout => \transmit_module.n1825\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_5_lut_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7428\,
            in2 => \_gnd_net_\,
            in3 => \N__6109\,
            lcout => \transmit_module.n201\,
            ltout => OPEN,
            carryin => \transmit_module.n1825\,
            carryout => \transmit_module.n1826\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_6_lut_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6105\,
            in2 => \_gnd_net_\,
            in3 => \N__6088\,
            lcout => \transmit_module.n200\,
            ltout => OPEN,
            carryin => \transmit_module.n1826\,
            carryout => \transmit_module.n1827\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_7_lut_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7515\,
            in2 => \_gnd_net_\,
            in3 => \N__6085\,
            lcout => \transmit_module.n199\,
            ltout => OPEN,
            carryin => \transmit_module.n1827\,
            carryout => \transmit_module.n1828\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_8_lut_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7335\,
            in2 => \_gnd_net_\,
            in3 => \N__6082\,
            lcout => \transmit_module.n198\,
            ltout => OPEN,
            carryin => \transmit_module.n1828\,
            carryout => \transmit_module.n1829\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_9_lut_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8575\,
            in2 => \_gnd_net_\,
            in3 => \N__6079\,
            lcout => \transmit_module.n197\,
            ltout => OPEN,
            carryin => \transmit_module.n1829\,
            carryout => \transmit_module.n1830\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_10_lut_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7494\,
            in2 => \_gnd_net_\,
            in3 => \N__6151\,
            lcout => \transmit_module.n196\,
            ltout => OPEN,
            carryin => \bfn_5_16_0_\,
            carryout => \transmit_module.n1831\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_11_lut_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6270\,
            in2 => \_gnd_net_\,
            in3 => \N__6148\,
            lcout => \transmit_module.n195\,
            ltout => OPEN,
            carryin => \transmit_module.n1831\,
            carryout => \transmit_module.n1832\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_12_lut_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7533\,
            in2 => \_gnd_net_\,
            in3 => \N__6145\,
            lcout => \transmit_module.n194\,
            ltout => OPEN,
            carryin => \transmit_module.n1832\,
            carryout => \transmit_module.n1833\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_13_lut_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7473\,
            in2 => \_gnd_net_\,
            in3 => \N__6142\,
            lcout => \transmit_module.n193\,
            ltout => OPEN,
            carryin => \transmit_module.n1833\,
            carryout => \transmit_module.n1834\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_14_lut_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7695\,
            in2 => \_gnd_net_\,
            in3 => \N__6139\,
            lcout => \transmit_module.n192\,
            ltout => OPEN,
            carryin => \transmit_module.n1834\,
            carryout => \transmit_module.n1835\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_15_lut_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8264\,
            in2 => \_gnd_net_\,
            in3 => \N__6136\,
            lcout => \transmit_module.n191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i9_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9549\,
            ce => \N__7641\,
            sr => \N__8995\
        );

    \transmit_module.BRAM_ADDR__i11_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__8520\,
            in1 => \N__6133\,
            in2 => \N__7462\,
            in3 => \N__8423\,
            lcout => \transmit_module.BRAM_ADDR_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9576\,
            ce => \N__8305\,
            sr => \N__8982\
        );

    \transmit_module.BRAM_ADDR__i8_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__8426\,
            in1 => \N__6127\,
            in2 => \N__7483\,
            in3 => \N__8527\,
            lcout => \transmit_module.BRAM_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9576\,
            ce => \N__8305\,
            sr => \N__8982\
        );

    \transmit_module.BRAM_ADDR__i12_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__8424\,
            in1 => \N__8524\,
            in2 => \N__7684\,
            in3 => \N__6121\,
            lcout => \transmit_module.BRAM_ADDR_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9576\,
            ce => \N__8305\,
            sr => \N__8982\
        );

    \transmit_module.BRAM_ADDR__i0_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__6295\,
            in1 => \N__7438\,
            in2 => \N__8548\,
            in3 => \N__8421\,
            lcout => \transmit_module.BRAM_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9576\,
            ce => \N__8305\,
            sr => \N__8982\
        );

    \transmit_module.BRAM_ADDR__i9_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__8427\,
            in1 => \N__8525\,
            in2 => \N__6286\,
            in3 => \N__6277\,
            lcout => \transmit_module.BRAM_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9576\,
            ce => \N__8305\,
            sr => \N__8982\
        );

    \transmit_module.BRAM_ADDR__i10_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__8519\,
            in1 => \N__7522\,
            in2 => \N__6262\,
            in3 => \N__8422\,
            lcout => \transmit_module.BRAM_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9576\,
            ce => \N__8305\,
            sr => \N__8982\
        );

    \transmit_module.BRAM_ADDR__i2_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__8425\,
            in1 => \N__6253\,
            in2 => \N__7660\,
            in3 => \N__8526\,
            lcout => \transmit_module.BRAM_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9576\,
            ce => \N__8305\,
            sr => \N__8982\
        );

    \transmit_module.video_signal_controller.i280_2_lut_3_lut_4_lut_rep_22_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__8410\,
            in1 => \N__6218\,
            in2 => \N__6192\,
            in3 => \N__8894\,
            lcout => \transmit_module.n2158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_9_3_lut_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6217\,
            in1 => \N__6185\,
            in2 => \_gnd_net_\,
            in3 => \N__8409\,
            lcout => OPEN,
            ltout => \transmit_module.n2145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1633_4_lut_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011100"
        )
    port map (
            in0 => \N__7893\,
            in1 => \N__8893\,
            in2 => \N__6244\,
            in3 => \N__6231\,
            lcout => \transmit_module.n704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_20_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6216\,
            in2 => \_gnd_net_\,
            in3 => \N__6181\,
            lcout => \transmit_module.n2156\,
            ltout => \transmit_module.n2156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__8411\,
            in1 => \N__7894\,
            in2 => \N__6154\,
            in3 => \N__8895\,
            lcout => \transmit_module.n792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i1_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6433\,
            in2 => \_gnd_net_\,
            in3 => \N__6415\,
            lcout => \transmit_module.video_signal_controller.VGA_X_0\,
            ltout => OPEN,
            carryin => \bfn_5_19_0_\,
            carryout => \transmit_module.video_signal_controller.n1844\,
            clk => \N__9539\,
            ce => 'H',
            sr => \N__6748\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i2_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7206\,
            in2 => \_gnd_net_\,
            in3 => \N__6412\,
            lcout => \transmit_module.video_signal_controller.VGA_X_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1844\,
            carryout => \transmit_module.video_signal_controller.n1845\,
            clk => \N__9539\,
            ce => 'H',
            sr => \N__6748\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i3_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6708\,
            in2 => \_gnd_net_\,
            in3 => \N__6409\,
            lcout => \transmit_module.video_signal_controller.VGA_X_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1845\,
            carryout => \transmit_module.video_signal_controller.n1846\,
            clk => \N__9539\,
            ce => 'H',
            sr => \N__6748\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i4_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6401\,
            in2 => \_gnd_net_\,
            in3 => \N__6376\,
            lcout => \transmit_module.video_signal_controller.VGA_X_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1846\,
            carryout => \transmit_module.video_signal_controller.n1847\,
            clk => \N__9539\,
            ce => 'H',
            sr => \N__6748\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i5_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6555\,
            in2 => \_gnd_net_\,
            in3 => \N__6373\,
            lcout => \transmit_module.video_signal_controller.VGA_X_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1847\,
            carryout => \transmit_module.video_signal_controller.n1848\,
            clk => \N__9539\,
            ce => 'H',
            sr => \N__6748\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i6_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7162\,
            in2 => \_gnd_net_\,
            in3 => \N__6370\,
            lcout => \transmit_module.video_signal_controller.VGA_X_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1848\,
            carryout => \transmit_module.video_signal_controller.n1849\,
            clk => \N__9539\,
            ce => 'H',
            sr => \N__6748\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i7_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6366\,
            in2 => \_gnd_net_\,
            in3 => \N__6331\,
            lcout => \transmit_module.video_signal_controller.VGA_X_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1849\,
            carryout => \transmit_module.video_signal_controller.n1850\,
            clk => \N__9539\,
            ce => 'H',
            sr => \N__6748\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i8_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7258\,
            in2 => \_gnd_net_\,
            in3 => \N__6328\,
            lcout => \transmit_module.video_signal_controller.VGA_X_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1850\,
            carryout => \transmit_module.video_signal_controller.n1851\,
            clk => \N__9539\,
            ce => 'H',
            sr => \N__6748\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i9_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6322\,
            in2 => \_gnd_net_\,
            in3 => \N__6838\,
            lcout => \transmit_module.video_signal_controller.VGA_X_8\,
            ltout => OPEN,
            carryin => \bfn_5_20_0_\,
            carryout => \transmit_module.video_signal_controller.n1852\,
            clk => \N__9423\,
            ce => 'H',
            sr => \N__6758\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i10_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6831\,
            in2 => \_gnd_net_\,
            in3 => \N__6802\,
            lcout => \transmit_module.video_signal_controller.VGA_X_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n1852\,
            carryout => \transmit_module.video_signal_controller.n1853\,
            clk => \N__9423\,
            ce => 'H',
            sr => \N__6758\
        );

    \transmit_module.video_signal_controller.VGA_X_275_276__i11_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6795\,
            in2 => \_gnd_net_\,
            in3 => \N__6799\,
            lcout => \transmit_module.video_signal_controller.VGA_X_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9423\,
            ce => 'H',
            sr => \N__6758\
        );

    \ADV_G__i3_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6709\,
            lcout => \ADV_G_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i3C_net\,
            ce => 'H',
            sr => \N__6882\
        );

    \ADV_B__i5_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6670\,
            lcout => \ADV_B_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i3C_net\,
            ce => 'H',
            sr => \N__6882\
        );

    \ADV_B__i1_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6604\,
            lcout => \ADV_B_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i3C_net\,
            ce => 'H',
            sr => \N__6882\
        );

    \ADV_G__i5_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6556\,
            lcout => \ADV_G_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i3C_net\,
            ce => 'H',
            sr => \N__6882\
        );

    \ADV_B__i8_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7035\,
            lcout => \ADV_B_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i3C_net\,
            ce => 'H',
            sr => \N__6882\
        );

    \ADV_B__i2_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6490\,
            lcout => \ADV_B_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i3C_net\,
            ce => 'H',
            sr => \N__6882\
        );

    \ADV_G__i8_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7261\,
            lcout => \ADV_G_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i3C_net\,
            ce => 'H',
            sr => \N__6882\
        );

    \ADV_G__i2_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7207\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ADV_G_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i2C_net\,
            ce => 'H',
            sr => \N__6889\
        );

    \ADV_G__i6_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7167\,
            lcout => \ADV_G_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i2C_net\,
            ce => 'H',
            sr => \N__6889\
        );

    \ADV_B__i7_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7111\,
            lcout => \ADV_B_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i2C_net\,
            ce => 'H',
            sr => \N__6889\
        );

    \ADV_R__i8_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7036\,
            lcout => \ADV_R_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i2C_net\,
            ce => 'H',
            sr => \N__6889\
        );

    \ADV_B__i3_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6976\,
            lcout => \ADV_B_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_G__i2C_net\,
            ce => 'H',
            sr => \N__6889\
        );

    \transmit_module.Y_DELTA_PATTERN_i3_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7312\,
            lcout => \transmit_module.Y_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9449\,
            ce => \N__9070\,
            sr => \N__8960\
        );

    \transmit_module.Y_DELTA_PATTERN_i99_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7886\,
            lcout => \transmit_module.Y_DELTA_PATTERN_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9449\,
            ce => \N__9070\,
            sr => \N__8960\
        );

    \transmit_module.Y_DELTA_PATTERN_i5_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7927\,
            lcout => \transmit_module.Y_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9449\,
            ce => \N__9070\,
            sr => \N__8960\
        );

    \transmit_module.Y_DELTA_PATTERN_i4_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7318\,
            lcout => \transmit_module.Y_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9449\,
            ce => \N__9070\,
            sr => \N__8960\
        );

    \transmit_module.Y_DELTA_PATTERN_i2_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7306\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9332\,
            ce => \N__9116\,
            sr => \N__8994\
        );

    \transmit_module.Y_DELTA_PATTERN_i1_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7300\,
            lcout => \transmit_module.Y_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9332\,
            ce => \N__9116\,
            sr => \N__8994\
        );

    \receive_module.rx_counter.i3_3_lut_4_lut_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__8067\,
            in1 => \N__8092\,
            in2 => \N__8119\,
            in3 => \N__8050\,
            lcout => \receive_module.rx_counter.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i444_2_lut_rep_17_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8048\,
            in2 => \_gnd_net_\,
            in3 => \N__8066\,
            lcout => \receive_module.rx_counter.n2153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8021\,
            in2 => \_gnd_net_\,
            in3 => \N__8143\,
            lcout => \receive_module.rx_counter.n7_adj_574\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__8113\,
            in1 => \N__7833\,
            in2 => \N__8146\,
            in3 => \N__8163\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n2063_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_4_lut_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__7402\,
            in1 => \N__7987\,
            in2 => \N__7276\,
            in3 => \N__8090\,
            lcout => \receive_module.rx_counter.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_18_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7832\,
            in2 => \_gnd_net_\,
            in3 => \N__8162\,
            lcout => \receive_module.rx_counter.n2007\,
            ltout => \receive_module.rx_counter.n2007_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_adj_20_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__8144\,
            in1 => \N__8089\,
            in2 => \N__7408\,
            in3 => \N__8114\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n2069_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8020\,
            in1 => \N__7988\,
            in2 => \N__7405\,
            in3 => \N__7401\,
            lcout => \receive_module.rx_counter.n2071\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i32_1_lut_rep_12_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7867\,
            lcout => n2148,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i6_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7336\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9531\,
            ce => \N__7650\,
            sr => \N__8977\
        );

    \transmit_module.ADDR_Y_COMPONENT__i7_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8571\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9531\,
            ce => \N__7650\,
            sr => \N__8977\
        );

    \transmit_module.BRAM_ADDR__i5_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__8445\,
            in1 => \N__7504\,
            in2 => \N__8555\,
            in3 => \N__7363\,
            lcout => \transmit_module.BRAM_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9569\,
            ce => \N__8316\,
            sr => \N__8998\
        );

    \transmit_module.BRAM_ADDR__i1_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__7357\,
            in1 => \N__8537\,
            in2 => \N__7543\,
            in3 => \N__8443\,
            lcout => \transmit_module.BRAM_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9569\,
            ce => \N__8316\,
            sr => \N__8998\
        );

    \transmit_module.BRAM_ADDR__i6_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__8446\,
            in1 => \N__7351\,
            in2 => \N__8556\,
            in3 => \N__7342\,
            lcout => \transmit_module.BRAM_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9569\,
            ce => \N__8316\,
            sr => \N__8998\
        );

    \transmit_module.BRAM_ADDR__i3_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__8444\,
            in1 => \N__7417\,
            in2 => \N__8554\,
            in3 => \N__7324\,
            lcout => \transmit_module.BRAM_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9569\,
            ce => \N__8316\,
            sr => \N__8998\
        );

    \transmit_module.ADDR_Y_COMPONENT__i1_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7555\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9462\,
            ce => \N__7645\,
            sr => \N__8975\
        );

    \transmit_module.ADDR_Y_COMPONENT__i10_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7534\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9462\,
            ce => \N__7645\,
            sr => \N__8975\
        );

    \transmit_module.ADDR_Y_COMPONENT__i5_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7516\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9462\,
            ce => \N__7645\,
            sr => \N__8975\
        );

    \transmit_module.ADDR_Y_COMPONENT__i13_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9462\,
            ce => \N__7645\,
            sr => \N__8975\
        );

    \transmit_module.ADDR_Y_COMPONENT__i8_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7495\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9541\,
            ce => \N__7649\,
            sr => \N__8968\
        );

    \transmit_module.ADDR_Y_COMPONENT__i11_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7474\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9541\,
            ce => \N__7649\,
            sr => \N__8968\
        );

    \transmit_module.ADDR_Y_COMPONENT__i0_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7452\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9541\,
            ce => \N__7649\,
            sr => \N__8968\
        );

    \transmit_module.ADDR_Y_COMPONENT__i3_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7432\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9541\,
            ce => \N__7649\,
            sr => \N__8968\
        );

    \transmit_module.ADDR_Y_COMPONENT__i12_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7696\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9541\,
            ce => \N__7649\,
            sr => \N__8968\
        );

    \transmit_module.ADDR_Y_COMPONENT__i2_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7674\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9541\,
            ce => \N__7649\,
            sr => \N__8968\
        );

    \transmit_module.X_DELTA_PATTERN_i7_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7759\,
            lcout => \transmit_module.X_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9461\,
            ce => \N__8206\,
            sr => \N__9048\
        );

    \transmit_module.X_DELTA_PATTERN_i1_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7600\,
            lcout => \transmit_module.X_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9461\,
            ce => \N__8206\,
            sr => \N__9048\
        );

    \transmit_module.X_DELTA_PATTERN_i2_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7588\,
            lcout => \transmit_module.X_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9461\,
            ce => \N__8206\,
            sr => \N__9048\
        );

    \transmit_module.X_DELTA_PATTERN_i4_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7741\,
            lcout => \transmit_module.X_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9461\,
            ce => \N__8206\,
            sr => \N__9048\
        );

    \transmit_module.X_DELTA_PATTERN_i3_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7594\,
            lcout => \transmit_module.X_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9461\,
            ce => \N__8206\,
            sr => \N__9048\
        );

    \transmit_module.X_DELTA_PATTERN_i0_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7582\,
            lcout => \transmit_module.X_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9461\,
            ce => \N__8206\,
            sr => \N__9048\
        );

    \transmit_module.X_DELTA_PATTERN_i15_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7569\,
            lcout => \transmit_module.X_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8192\,
            sr => \N__9085\
        );

    \transmit_module.X_DELTA_PATTERN_i6_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7771\,
            lcout => \transmit_module.X_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8192\,
            sr => \N__9085\
        );

    \transmit_module.X_DELTA_PATTERN_i9_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8230\,
            lcout => \transmit_module.X_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8192\,
            sr => \N__9085\
        );

    \transmit_module.X_DELTA_PATTERN_i8_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7765\,
            lcout => \transmit_module.X_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8192\,
            sr => \N__9085\
        );

    \transmit_module.X_DELTA_PATTERN_i14_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7753\,
            lcout => \transmit_module.X_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8192\,
            sr => \N__9085\
        );

    \transmit_module.X_DELTA_PATTERN_i5_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7747\,
            lcout => \transmit_module.X_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8192\,
            sr => \N__9085\
        );

    \transmit_module.X_DELTA_PATTERN_i13_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7735\,
            lcout => \transmit_module.X_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8192\,
            sr => \N__9085\
        );

    \transmit_module.Y_DELTA_PATTERN_i32_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7729\,
            lcout => \transmit_module.Y_DELTA_PATTERN_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => \N__9099\,
            sr => \N__8843\
        );

    \transmit_module.Y_DELTA_PATTERN_i31_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7714\,
            lcout => \transmit_module.Y_DELTA_PATTERN_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => \N__9099\,
            sr => \N__8843\
        );

    \transmit_module.Y_DELTA_PATTERN_i29_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7702\,
            lcout => \transmit_module.Y_DELTA_PATTERN_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => \N__9099\,
            sr => \N__8843\
        );

    \transmit_module.Y_DELTA_PATTERN_i30_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7708\,
            lcout => \transmit_module.Y_DELTA_PATTERN_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => \N__9099\,
            sr => \N__8843\
        );

    \transmit_module.Y_DELTA_PATTERN_i17_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7804\,
            lcout => \transmit_module.Y_DELTA_PATTERN_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => \N__9109\,
            sr => \N__8950\
        );

    \transmit_module.Y_DELTA_PATTERN_i20_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7792\,
            lcout => \transmit_module.Y_DELTA_PATTERN_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => \N__9109\,
            sr => \N__8950\
        );

    \transmit_module.Y_DELTA_PATTERN_i19_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7816\,
            lcout => \transmit_module.Y_DELTA_PATTERN_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => \N__9109\,
            sr => \N__8950\
        );

    \transmit_module.Y_DELTA_PATTERN_i22_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7909\,
            lcout => \transmit_module.Y_DELTA_PATTERN_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => \N__9109\,
            sr => \N__8950\
        );

    \transmit_module.Y_DELTA_PATTERN_i18_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7810\,
            lcout => \transmit_module.Y_DELTA_PATTERN_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => \N__9109\,
            sr => \N__8950\
        );

    \transmit_module.Y_DELTA_PATTERN_i21_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7798\,
            lcout => \transmit_module.Y_DELTA_PATTERN_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => \N__9109\,
            sr => \N__8950\
        );

    \transmit_module.Y_DELTA_PATTERN_i16_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7786\,
            lcout => \transmit_module.Y_DELTA_PATTERN_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => \N__9109\,
            sr => \N__8950\
        );

    \transmit_module.Y_DELTA_PATTERN_i28_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7780\,
            lcout => \transmit_module.Y_DELTA_PATTERN_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9384\,
            ce => \N__9115\,
            sr => \N__8916\
        );

    \transmit_module.Y_DELTA_PATTERN_i26_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7939\,
            lcout => \transmit_module.Y_DELTA_PATTERN_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9384\,
            ce => \N__9115\,
            sr => \N__8916\
        );

    \transmit_module.Y_DELTA_PATTERN_i27_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7945\,
            lcout => \transmit_module.Y_DELTA_PATTERN_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9384\,
            ce => \N__9115\,
            sr => \N__8916\
        );

    \transmit_module.Y_DELTA_PATTERN_i25_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7933\,
            lcout => \transmit_module.Y_DELTA_PATTERN_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9384\,
            ce => \N__9115\,
            sr => \N__8916\
        );

    \transmit_module.Y_DELTA_PATTERN_i6_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9604\,
            lcout => \transmit_module.Y_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9447\,
            ce => \N__9110\,
            sr => \N__8964\
        );

    \transmit_module.Y_DELTA_PATTERN_i24_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7921\,
            lcout => \transmit_module.Y_DELTA_PATTERN_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9447\,
            ce => \N__9110\,
            sr => \N__8964\
        );

    \transmit_module.Y_DELTA_PATTERN_i23_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7915\,
            lcout => \transmit_module.Y_DELTA_PATTERN_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9447\,
            ce => \N__9110\,
            sr => \N__8964\
        );

    \transmit_module.Y_DELTA_PATTERN_i0_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7900\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9280\,
            ce => \N__9117\,
            sr => \N__8978\
        );

    \receive_module.rx_counter.i281_3_lut_3_lut_3_lut_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__9924\,
            in1 => \N__7862\,
            in2 => \_gnd_net_\,
            in3 => \N__7840\,
            lcout => \receive_module.rx_counter.n752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_HS_50_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7863\,
            lcout => \receive_module.rx_counter.old_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.Y__i0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7834\,
            in2 => \_gnd_net_\,
            in3 => \N__7819\,
            lcout => \receive_module.rx_counter.Y_0\,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \receive_module.rx_counter.n1836\,
            clk => \N__9861\,
            ce => \N__7966\,
            sr => \N__8635\
        );

    \receive_module.rx_counter.Y__i1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8164\,
            in2 => \_gnd_net_\,
            in3 => \N__8149\,
            lcout => \receive_module.rx_counter.Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1836\,
            carryout => \receive_module.rx_counter.n1837\,
            clk => \N__9861\,
            ce => \N__7966\,
            sr => \N__8635\
        );

    \receive_module.rx_counter.Y__i2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8145\,
            in2 => \_gnd_net_\,
            in3 => \N__8122\,
            lcout => \receive_module.rx_counter.Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1837\,
            carryout => \receive_module.rx_counter.n1838\,
            clk => \N__9861\,
            ce => \N__7966\,
            sr => \N__8635\
        );

    \receive_module.rx_counter.Y__i3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8118\,
            in2 => \_gnd_net_\,
            in3 => \N__8095\,
            lcout => \receive_module.rx_counter.Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1838\,
            carryout => \receive_module.rx_counter.n1839\,
            clk => \N__9861\,
            ce => \N__7966\,
            sr => \N__8635\
        );

    \receive_module.rx_counter.Y__i4_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8091\,
            in2 => \_gnd_net_\,
            in3 => \N__8071\,
            lcout => \receive_module.rx_counter.Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1839\,
            carryout => \receive_module.rx_counter.n1840\,
            clk => \N__9861\,
            ce => \N__7966\,
            sr => \N__8635\
        );

    \receive_module.rx_counter.Y__i5_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8068\,
            in2 => \_gnd_net_\,
            in3 => \N__8053\,
            lcout => \receive_module.rx_counter.Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1840\,
            carryout => \receive_module.rx_counter.n1841\,
            clk => \N__9861\,
            ce => \N__7966\,
            sr => \N__8635\
        );

    \receive_module.rx_counter.Y__i6_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8049\,
            in2 => \_gnd_net_\,
            in3 => \N__8032\,
            lcout => \receive_module.rx_counter.Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1841\,
            carryout => \receive_module.rx_counter.n1842\,
            clk => \N__9861\,
            ce => \N__7966\,
            sr => \N__8635\
        );

    \receive_module.rx_counter.Y__i7_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8025\,
            in2 => \_gnd_net_\,
            in3 => \N__8002\,
            lcout => \receive_module.rx_counter.Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1842\,
            carryout => \receive_module.rx_counter.n1843\,
            clk => \N__9861\,
            ce => \N__7966\,
            sr => \N__8635\
        );

    \receive_module.rx_counter.Y__i8_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7992\,
            in2 => \_gnd_net_\,
            in3 => \N__7999\,
            lcout => \receive_module.rx_counter.Y_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9862\,
            ce => \N__7965\,
            sr => \N__8640\
        );

    \transmit_module.BRAM_ADDR__i7_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__8557\,
            in1 => \N__8596\,
            in2 => \N__8584\,
            in3 => \N__8442\,
            lcout => \transmit_module.BRAM_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9570\,
            ce => \N__8320\,
            sr => \N__8990\
        );

    \transmit_module.video_signal_controller.i960_3_lut_4_lut_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__8550\,
            in1 => \N__8464\,
            in2 => \N__8455\,
            in3 => \N__8441\,
            lcout => \transmit_module.BRAM_ADDR_13_N_257_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i13_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8251\,
            in1 => \N__8329\,
            in2 => \_gnd_net_\,
            in3 => \N__8304\,
            lcout => \DEBUG_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9532\,
            ce => 'H',
            sr => \N__8992\
        );

    \transmit_module.X_DELTA_PATTERN_i10_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8224\,
            lcout => \transmit_module.X_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9471\,
            ce => \N__8205\,
            sr => \N__9086\
        );

    \transmit_module.X_DELTA_PATTERN_i11_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8212\,
            lcout => \transmit_module.X_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9471\,
            ce => \N__8205\,
            sr => \N__9086\
        );

    \transmit_module.X_DELTA_PATTERN_i12_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8218\,
            lcout => \transmit_module.X_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9471\,
            ce => \N__8205\,
            sr => \N__9086\
        );

    \transmit_module.Y_DELTA_PATTERN_i15_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8176\,
            lcout => \transmit_module.Y_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9460\,
            ce => \N__9084\,
            sr => \N__8991\
        );

    \transmit_module.Y_DELTA_PATTERN_i14_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8170\,
            lcout => \transmit_module.Y_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9460\,
            ce => \N__9084\,
            sr => \N__8991\
        );

    \transmit_module.Y_DELTA_PATTERN_i13_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9634\,
            lcout => \transmit_module.Y_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9460\,
            ce => \N__9084\,
            sr => \N__8991\
        );

    \transmit_module.Y_DELTA_PATTERN_i12_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9628\,
            lcout => \transmit_module.Y_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9460\,
            ce => \N__9084\,
            sr => \N__8991\
        );

    \transmit_module.Y_DELTA_PATTERN_i9_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9610\,
            lcout => \transmit_module.Y_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9383\,
            ce => \N__9114\,
            sr => \N__8993\
        );

    \transmit_module.Y_DELTA_PATTERN_i11_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9622\,
            lcout => \transmit_module.Y_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9383\,
            ce => \N__9114\,
            sr => \N__8993\
        );

    \transmit_module.Y_DELTA_PATTERN_i10_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9616\,
            lcout => \transmit_module.Y_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9383\,
            ce => \N__9114\,
            sr => \N__8993\
        );

    \transmit_module.Y_DELTA_PATTERN_i7_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9592\,
            lcout => \transmit_module.Y_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9360\,
            ce => \N__9121\,
            sr => \N__8979\
        );

    \transmit_module.Y_DELTA_PATTERN_i8_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9598\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9360\,
            ce => \N__9121\,
            sr => \N__8979\
        );

    \receive_module.rx_counter.FRAME_COUNTER_273__i0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9673\,
            in2 => \_gnd_net_\,
            in3 => \N__8650\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_0\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \receive_module.rx_counter.n1865\,
            clk => \N__9860\,
            ce => \N__9709\,
            sr => \N__9949\
        );

    \receive_module.rx_counter.FRAME_COUNTER_273__i1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9685\,
            in2 => \_gnd_net_\,
            in3 => \N__8647\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1865\,
            carryout => \receive_module.rx_counter.n1866\,
            clk => \N__9860\,
            ce => \N__9709\,
            sr => \N__9949\
        );

    \receive_module.rx_counter.FRAME_COUNTER_273__i2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9721\,
            in2 => \_gnd_net_\,
            in3 => \N__9766\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1866\,
            carryout => \receive_module.rx_counter.n1867\,
            clk => \N__9860\,
            ce => \N__9709\,
            sr => \N__9949\
        );

    \receive_module.rx_counter.FRAME_COUNTER_273__i3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9661\,
            in2 => \_gnd_net_\,
            in3 => \N__9763\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1867\,
            carryout => \receive_module.rx_counter.n1868\,
            clk => \N__9860\,
            ce => \N__9709\,
            sr => \N__9949\
        );

    \receive_module.rx_counter.FRAME_COUNTER_273__i4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9733\,
            in2 => \_gnd_net_\,
            in3 => \N__9760\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n1868\,
            carryout => \receive_module.rx_counter.n1869\,
            clk => \N__9860\,
            ce => \N__9709\,
            sr => \N__9949\
        );

    \receive_module.rx_counter.FRAME_COUNTER_273__i5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9697\,
            in2 => \_gnd_net_\,
            in3 => \N__9757\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9860\,
            ce => \N__9709\,
            sr => \N__9949\
        );

    \receive_module.rx_counter.PULSE_1HZ_48_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9744\,
            in2 => \_gnd_net_\,
            in3 => \N__9640\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9857\,
            ce => \N__9708\,
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9732\,
            in2 => \_gnd_net_\,
            in3 => \N__9720\,
            lcout => \receive_module.rx_counter.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i435_2_lut_rep_14_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__9932\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9880\,
            lcout => \receive_module.rx_counter.n2150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1950_2_lut_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9696\,
            in2 => \_gnd_net_\,
            in3 => \N__9684\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n2113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_4_lut_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__9672\,
            in1 => \N__9660\,
            in2 => \N__9649\,
            in3 => \N__9646\,
            lcout => \receive_module.rx_counter.n11\,
            ltout => \receive_module.rx_counter.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1077_2_lut_3_lut_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__9931\,
            in1 => \_gnd_net_\,
            in2 => \N__9952\,
            in3 => \N__9879\,
            lcout => \receive_module.rx_counter.n1328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_VS_51_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9930\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.rx_counter.old_VS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9871\,
            lcout => \GB_BUFFER_TVP_CLK_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
