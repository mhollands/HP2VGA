// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Sat Sep 29 12:22:35 2018
//
// Verilog Description of module main
//

module main (DEBUG, TVP_CLK, TVP_HSYNC, TVP_VSYNC, TVP_VIDEO, LED, 
            ADV_HSYNC, ADV_VSYNC, ADV_R, ADV_G, ADV_B, ADV_CLK, 
            ADV_SYNC_N, ADV_BLANK_N) /* synthesis syn_module_defined=1 */ ;   // ../main.v(1[8:12])
    output [7:0]DEBUG;   // ../main.v(2[19:24])
    input TVP_CLK;   // ../main.v(3[13:20])
    input TVP_HSYNC;   // ../main.v(4[13:22])
    input TVP_VSYNC;   // ../main.v(5[13:22])
    input [9:0]TVP_VIDEO;   // ../main.v(6[19:28])
    output LED;   // ../main.v(7[14:17])
    output ADV_HSYNC;   // ../main.v(8[14:23])
    output ADV_VSYNC;   // ../main.v(9[14:23])
    output [7:0]ADV_R;   // ../main.v(10[20:25])
    output [7:0]ADV_G;   // ../main.v(11[20:25])
    output [7:0]ADV_B;   // ../main.v(12[20:25])
    output ADV_CLK;   // ../main.v(13[14:21])
    output ADV_SYNC_N;   // ../main.v(14[14:24])
    output ADV_BLANK_N;   // ../main.v(15[14:25])
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    
    wire GND_net, VCC_net, TVP_HSYNC_c, TVP_VSYNC_c, TVP_VIDEO_c_9, 
        TVP_VIDEO_c_8, TVP_VIDEO_c_7, TVP_VIDEO_c_6, TVP_VIDEO_c_5, 
        TVP_VIDEO_c_4, TVP_VIDEO_c_3, TVP_VIDEO_c_2, LED_c, ADV_HSYNC_c, 
        ADV_VSYNC_c, ADV_B_c, n1792, n1793, n1794, n1795, n1796, 
        n1797, n1798, RX_TX_SYNC;
    wire [13:0]RX_ADDR;   // ../main.v(28[14:21])
    
    wire RX_WE;
    wire [13:0]TX_ADDR;   // ../main.v(51[14:21])
    wire [7:0]TX_DATA;   // ../main.v(52[13:20])
    
    wire RX_TX_SYNC_BUFF, n27, n28, n22, n20, n18, n21, n26, 
        n25, n24, n23, n19;
    
    VCC i2 (.Y(VCC_net));
    INPUT_BUFFER sync_buffer (.RX_TX_SYNC(RX_TX_SYNC), .ADV_CLK_c(ADV_CLK_c), 
            .RX_TX_SYNC_BUFF(RX_TX_SYNC_BUFF)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(73[15:90])
    TX transmit_module (.ADV_CLK_c(ADV_CLK_c), .ADV_VSYNC_c(ADV_VSYNC_c), 
       .ADV_HSYNC_c(ADV_HSYNC_c), .n28(n28), .GND_net(GND_net), .TX_DATA({TX_DATA}), 
       .ADV_B_c(ADV_B_c), .n26(n26), .n1792(n1792), .n27(n27), .n1793(n1793), 
       .n1794(n1794), .n1795(n1795), .n1796(n1796), .n1797(n1797), .n18(n18), 
       .n25(n25), .n19(n19), .n20(n20), .n21(n21), .\TX_ADDR[13] (TX_ADDR[13]), 
       .\TX_ADDR[12] (TX_ADDR[12]), .n22(n22), .n24(n24), .n23(n23), 
       .\TX_ADDR[11] (TX_ADDR[11]), .n1798(n1798), .VCC_net(VCC_net), 
       .RX_TX_SYNC_BUFF(RX_TX_SYNC_BUFF)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(58[5] 71[26])
    SB_IO ADV_B_pad_2 (.PACKAGE_PIN(ADV_B[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1796));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_2.PULLUP = 1'b0;
    defparam ADV_B_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_1 (.PACKAGE_PIN(ADV_B[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1797));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_1.PULLUP = 1'b0;
    defparam ADV_B_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_4 (.PACKAGE_PIN(ADV_B[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1794));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_4.PULLUP = 1'b0;
    defparam ADV_B_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_5 (.PACKAGE_PIN(ADV_B[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1793));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_5.PULLUP = 1'b0;
    defparam ADV_B_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_1 (.PACKAGE_PIN(ADV_R[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1797));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_1.PULLUP = 1'b0;
    defparam ADV_R_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_2 (.PACKAGE_PIN(ADV_R[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1796));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_2.PULLUP = 1'b0;
    defparam ADV_R_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_3 (.PACKAGE_PIN(ADV_R[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1795));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_3.PULLUP = 1'b0;
    defparam ADV_R_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_4 (.PACKAGE_PIN(ADV_R[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1794));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_4.PULLUP = 1'b0;
    defparam ADV_R_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_5 (.PACKAGE_PIN(ADV_R[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1793));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_5.PULLUP = 1'b0;
    defparam ADV_R_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_6 (.PACKAGE_PIN(ADV_R[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1792));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_6.PULLUP = 1'b0;
    defparam ADV_R_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_6 (.PACKAGE_PIN(ADV_B[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1792));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_6.PULLUP = 1'b0;
    defparam ADV_B_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_7 (.PACKAGE_PIN(ADV_B[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_7.PULLUP = 1'b0;
    defparam ADV_B_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_0 (.PACKAGE_PIN(ADV_G[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1798));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_0.PULLUP = 1'b0;
    defparam ADV_G_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_7 (.PACKAGE_PIN(ADV_R[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_7.PULLUP = 1'b0;
    defparam ADV_R_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_VSYNC_pad (.PACKAGE_PIN(ADV_VSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_VSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_VSYNC_pad.PIN_TYPE = 6'b011001;
    defparam ADV_VSYNC_pad.PULLUP = 1'b0;
    defparam ADV_VSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_VSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_HSYNC_pad (.PACKAGE_PIN(ADV_HSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_HSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_HSYNC_pad.PIN_TYPE = 6'b011001;
    defparam ADV_HSYNC_pad.PULLUP = 1'b0;
    defparam ADV_HSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_HSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_0 (.PACKAGE_PIN(DEBUG[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_0.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_0.PULLUP = 1'b0;
    defparam DEBUG_pad_0.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_1 (.PACKAGE_PIN(DEBUG[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_1.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_1.PULLUP = 1'b0;
    defparam DEBUG_pad_1.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_2 (.PACKAGE_PIN(DEBUG[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_2.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_2.PULLUP = 1'b0;
    defparam DEBUG_pad_2.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_3 (.PACKAGE_PIN(DEBUG[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_3.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_3.PULLUP = 1'b0;
    defparam DEBUG_pad_3.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_4 (.PACKAGE_PIN(DEBUG[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_4.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_4.PULLUP = 1'b0;
    defparam DEBUG_pad_4.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_1 (.PACKAGE_PIN(ADV_G[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1797));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_1.PULLUP = 1'b0;
    defparam ADV_G_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_2 (.PACKAGE_PIN(ADV_G[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1796));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_2.PULLUP = 1'b0;
    defparam ADV_G_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_3 (.PACKAGE_PIN(ADV_G[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1795));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_3.PULLUP = 1'b0;
    defparam ADV_G_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_4 (.PACKAGE_PIN(ADV_G[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1794));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_4.PULLUP = 1'b0;
    defparam ADV_G_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_5 (.PACKAGE_PIN(ADV_G[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1793));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_5.PULLUP = 1'b0;
    defparam ADV_G_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_6 (.PACKAGE_PIN(ADV_G[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1792));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_6.PULLUP = 1'b0;
    defparam ADV_G_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_7 (.PACKAGE_PIN(ADV_G[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_7.PULLUP = 1'b0;
    defparam ADV_G_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_0 (.PACKAGE_PIN(ADV_R[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1798));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_0.PULLUP = 1'b0;
    defparam ADV_R_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_6 (.PACKAGE_PIN(DEBUG[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_6.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_6.PULLUP = 1'b0;
    defparam DEBUG_pad_6.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_7 (.PACKAGE_PIN(DEBUG[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_7.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_7.PULLUP = 1'b0;
    defparam DEBUG_pad_7.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_5 (.PACKAGE_PIN(DEBUG[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_5.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_5.PULLUP = 1'b0;
    defparam DEBUG_pad_5.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_2 (.PACKAGE_PIN(TVP_VIDEO[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_2));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_2.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_2.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_2.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_3 (.PACKAGE_PIN(ADV_B[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1795));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_3.PULLUP = 1'b0;
    defparam ADV_B_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_3 (.PACKAGE_PIN(TVP_VIDEO[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_3));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_3.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_3.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_3.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_4 (.PACKAGE_PIN(TVP_VIDEO[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_4));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_4.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_4.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_4.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_5 (.PACKAGE_PIN(TVP_VIDEO[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_5));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_5.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_5.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_5.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_6 (.PACKAGE_PIN(TVP_VIDEO[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_6));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_6.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_6.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_6.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_7 (.PACKAGE_PIN(TVP_VIDEO[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_7));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_7.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_7.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_7.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_8 (.PACKAGE_PIN(TVP_VIDEO[8]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_8));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_8.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_8.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_8.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_8.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_9 (.PACKAGE_PIN(TVP_VIDEO[9]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_9));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_9.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_9.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_9.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_9.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VSYNC_pad (.PACKAGE_PIN(TVP_VSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VSYNC_pad.PIN_TYPE = 6'b000001;
    defparam TVP_VSYNC_pad.PULLUP = 1'b0;
    defparam TVP_VSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_VSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_HSYNC_pad (.PACKAGE_PIN(TVP_HSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_HSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_HSYNC_pad.PIN_TYPE = 6'b000001;
    defparam TVP_HSYNC_pad.PULLUP = 1'b0;
    defparam TVP_HSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_HSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO TVP_CLK_pad (.PACKAGE_PIN(TVP_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(TVP_CLK_c));   // ../main.v(3[13:20])
    defparam TVP_CLK_pad.PIN_TYPE = 6'b000001;
    defparam TVP_CLK_pad.PULLUP = 1'b0;
    defparam TVP_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_BLANK_N_pad (.PACKAGE_PIN(ADV_BLANK_N), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_BLANK_N_pad.PIN_TYPE = 6'b011001;
    defparam ADV_BLANK_N_pad.PULLUP = 1'b0;
    defparam ADV_BLANK_N_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_BLANK_N_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_SYNC_N_pad (.PACKAGE_PIN(ADV_SYNC_N), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_SYNC_N_pad.PIN_TYPE = 6'b011001;
    defparam ADV_SYNC_N_pad.PULLUP = 1'b0;
    defparam ADV_SYNC_N_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_SYNC_N_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_CLK_pad (.PACKAGE_PIN(ADV_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(ADV_CLK_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_CLK_pad.PIN_TYPE = 6'b011001;
    defparam ADV_CLK_pad.PULLUP = 1'b0;
    defparam ADV_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_0 (.PACKAGE_PIN(ADV_B[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1798));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_0.PULLUP = 1'b0;
    defparam ADV_B_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_0.IO_STANDARD = "SB_LVCMOS";
    RX receive_module (.RX_ADDR({RX_ADDR}), .GND_net(GND_net), .RX_WE(RX_WE), 
       .TVP_VSYNC_c(TVP_VSYNC_c), .TVP_CLK_c(TVP_CLK_c), .VCC_net(VCC_net), 
       .TVP_HSYNC_c(TVP_HSYNC_c), .RX_TX_SYNC(RX_TX_SYNC), .LED_c(LED_c)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(37[5] 48[29])
    GND i1 (.Y(GND_net));
    RAM line_buffer (.TX_DATA({TX_DATA}), .ADV_CLK_c(ADV_CLK_c), .\TX_ADDR[12] (TX_ADDR[12]), 
        .\TX_ADDR[13] (TX_ADDR[13]), .\TX_ADDR[11] (TX_ADDR[11]), .GND_net(GND_net), 
        .RX_ADDR({RX_ADDR}), .n28(n28), .n27(n27), .n26(n26), .n25(n25), 
        .n24(n24), .n23(n23), .n22(n22), .n21(n21), .n20(n20), .n19(n19), 
        .n18(n18), .TVP_VIDEO_c_8(TVP_VIDEO_c_8), .TVP_VIDEO_c_9(TVP_VIDEO_c_9), 
        .TVP_CLK_c(TVP_CLK_c), .VCC_net(VCC_net), .TVP_VIDEO_c_6(TVP_VIDEO_c_6), 
        .TVP_VIDEO_c_7(TVP_VIDEO_c_7), .TVP_VIDEO_c_4(TVP_VIDEO_c_4), .TVP_VIDEO_c_5(TVP_VIDEO_c_5), 
        .TVP_VIDEO_c_2(TVP_VIDEO_c_2), .TVP_VIDEO_c_3(TVP_VIDEO_c_3), .RX_WE(RX_WE)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(83[6] 89[21])
    TX_PLL tx_pll (.TVP_CLK_c(TVP_CLK_c), .VCC_net(VCC_net), .GND_net(GND_net), 
           .ADV_CLK_c(ADV_CLK_c)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(20[9] 24[27])
    
endmodule
//
// Verilog Description of module INPUT_BUFFER
//

module INPUT_BUFFER (RX_TX_SYNC, ADV_CLK_c, RX_TX_SYNC_BUFF) /* synthesis syn_module_defined=1 */ ;
    input RX_TX_SYNC;
    input ADV_CLK_c;
    output RX_TX_SYNC_BUFF;
    
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    wire [1:0]BUFFER;   // ../input_buffer.v(7[24:30])
    
    SB_DFFN BUFFER_i0 (.Q(BUFFER[0]), .C(ADV_CLK_c), .D(RX_TX_SYNC));   // ../input_buffer.v(9[9] 12[5])
    SB_DFFN WIRE_OUT_8 (.Q(RX_TX_SYNC_BUFF), .C(ADV_CLK_c), .D(BUFFER[1]));   // ../input_buffer.v(9[9] 12[5])
    SB_DFFN BUFFER_i1 (.Q(BUFFER[1]), .C(ADV_CLK_c), .D(BUFFER[0]));   // ../input_buffer.v(9[9] 12[5])
    
endmodule
//
// Verilog Description of module TX
//

module TX (ADV_CLK_c, ADV_VSYNC_c, ADV_HSYNC_c, n28, GND_net, TX_DATA, 
           ADV_B_c, n26, n1792, n27, n1793, n1794, n1795, n1796, 
           n1797, n18, n25, n19, n20, n21, \TX_ADDR[13] , \TX_ADDR[12] , 
           n22, n24, n23, \TX_ADDR[11] , n1798, VCC_net, RX_TX_SYNC_BUFF) /* synthesis syn_module_defined=1 */ ;
    input ADV_CLK_c;
    output ADV_VSYNC_c;
    output ADV_HSYNC_c;
    output n28;
    input GND_net;
    input [7:0]TX_DATA;
    output ADV_B_c;
    output n26;
    output n1792;
    output n27;
    output n1793;
    output n1794;
    output n1795;
    output n1796;
    output n1797;
    output n18;
    output n25;
    output n19;
    output n20;
    output n21;
    output \TX_ADDR[13] ;
    output \TX_ADDR[12] ;
    output n22;
    output n24;
    output n23;
    output \TX_ADDR[11] ;
    output n1798;
    input VCC_net;
    input RX_TX_SYNC_BUFF;
    
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    wire [99:0]Y_DELTA_PATTERN;   // ../tx.v(61[16:31])
    
    wire n3797, n2147, old_VGA_HS;
    wire [13:0]TX_ADDR;   // ../main.v(51[14:21])
    wire [13:0]ADDR_Y_COMPONENT;   // ../tx.v(62[16:32])
    wire [13:0]n102;
    
    wire n2354;
    wire [13:0]n118;
    
    wire VGA_VISIBLE;
    wire [13:0]n133;
    
    wire n3787, n3261, n3270, n3269, n3262, n3260, n3798;
    wire [13:0]BRAM_ADDR_13__N_282;
    
    wire n2061, n2039, n2093, n3268, n3267, n3259, n3258, n3266, 
        n3265;
    wire [15:0]X_DELTA_PATTERN;   // ../tx.v(60[16:31])
    
    wire n3264, n3263, VGA_VISIBLE_Y;
    
    SB_DFFESR Y_DELTA_PATTERN_i94 (.Q(Y_DELTA_PATTERN[94]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[95]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i93 (.Q(Y_DELTA_PATTERN[93]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[94]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFF old_VGA_HS_40 (.Q(old_VGA_HS), .C(ADV_CLK_c), .D(ADV_HSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i0 (.Q(TX_ADDR[0]), .C(ADV_CLK_c), .D(n28));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i92 (.Q(Y_DELTA_PATTERN[92]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[93]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i91 (.Q(Y_DELTA_PATTERN[91]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[92]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i90 (.Q(Y_DELTA_PATTERN[90]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[91]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_12_i3_3_lut (.I0(ADDR_Y_COMPONENT[2]), .I1(TX_ADDR[2]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[2]));   // ../tx.v(83[30:81])
    defparam mux_12_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR VGA_R__i8 (.Q(ADV_B_c), .C(ADV_CLK_c), .D(TX_DATA[7]), .R(n2354));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_14_i3_3_lut (.I0(TX_ADDR[2]), .I1(n118[2]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[2]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1601_4_lut (.I0(n133[2]), .I1(ADV_VSYNC_c), .I2(n102[2]), 
            .I3(n3787), .O(n26));   // ../tx.v(68[12] 94[8])
    defparam i1601_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS Y_DELTA_PATTERN_i89 (.Q(Y_DELTA_PATTERN[89]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[90]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_12_i2_3_lut (.I0(ADDR_Y_COMPONENT[1]), .I1(TX_ADDR[1]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[1]));   // ../tx.v(83[30:81])
    defparam mux_12_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_13_6_lut (.I0(GND_net), .I1(TX_ADDR[4]), .I2(GND_net), 
            .I3(n3261), .O(n118[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR VGA_R__i7 (.Q(n1792), .C(ADV_CLK_c), .D(TX_DATA[6]), .R(n2354));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_14_i2_3_lut (.I0(TX_ADDR[1]), .I1(n118[1]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[1]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1600_4_lut (.I0(n133[1]), .I1(ADV_VSYNC_c), .I2(n102[1]), 
            .I3(n3787), .O(n27));   // ../tx.v(68[12] 94[8])
    defparam i1600_4_lut.LUT_INIT = 16'h3022;
    SB_DFFSR VGA_R__i6 (.Q(n1793), .C(ADV_CLK_c), .D(TX_DATA[5]), .R(n2354));   // ../tx.v(68[12] 94[8])
    SB_DFFSR VGA_R__i5 (.Q(n1794), .C(ADV_CLK_c), .D(TX_DATA[4]), .R(n2354));   // ../tx.v(68[12] 94[8])
    SB_DFFSR VGA_R__i4 (.Q(n1795), .C(ADV_CLK_c), .D(TX_DATA[3]), .R(n2354));   // ../tx.v(68[12] 94[8])
    SB_DFFSR VGA_R__i3 (.Q(n1796), .C(ADV_CLK_c), .D(TX_DATA[2]), .R(n2354));   // ../tx.v(68[12] 94[8])
    SB_DFFSR VGA_R__i2 (.Q(n1797), .C(ADV_CLK_c), .D(TX_DATA[1]), .R(n2354));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i10 (.Q(TX_ADDR[10]), .C(ADV_CLK_c), .D(n18));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_12_i4_3_lut (.I0(ADDR_Y_COMPONENT[3]), .I1(TX_ADDR[3]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[3]));   // ../tx.v(83[30:81])
    defparam mux_12_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i4_3_lut (.I0(TX_ADDR[3]), .I1(n118[3]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[3]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1602_4_lut (.I0(n133[3]), .I1(ADV_VSYNC_c), .I2(n102[3]), 
            .I3(n3787), .O(n25));   // ../tx.v(68[12] 94[8])
    defparam i1602_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i5_3_lut (.I0(ADDR_Y_COMPONENT[4]), .I1(TX_ADDR[4]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[4]));   // ../tx.v(83[30:81])
    defparam mux_12_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_12_i1_3_lut (.I0(ADDR_Y_COMPONENT[0]), .I1(TX_ADDR[0]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[0]));   // ../tx.v(83[30:81])
    defparam mux_12_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i1_3_lut (.I0(TX_ADDR[0]), .I1(n118[0]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[0]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1595_4_lut (.I0(n133[0]), .I1(ADV_VSYNC_c), .I2(n102[0]), 
            .I3(n3787), .O(n28));   // ../tx.v(68[12] 94[8])
    defparam i1595_4_lut.LUT_INIT = 16'h3022;
    SB_DFF BRAM_ADDR__i9 (.Q(TX_ADDR[9]), .C(ADV_CLK_c), .D(n19));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i98 (.Q(Y_DELTA_PATTERN[98]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[99]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i8 (.Q(TX_ADDR[8]), .C(ADV_CLK_c), .D(n20));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i7 (.Q(TX_ADDR[7]), .C(ADV_CLK_c), .D(n21));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_14_i5_3_lut (.I0(TX_ADDR[4]), .I1(n118[4]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[4]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_13_15_lut (.I0(GND_net), .I1(\TX_ADDR[13] ), .I2(GND_net), 
            .I3(n3270), .O(n118[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_14_lut (.I0(GND_net), .I1(\TX_ADDR[12] ), .I2(GND_net), 
            .I3(n3269), .O(n118[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_6 (.CI(n3261), .I0(TX_ADDR[4]), .I1(GND_net), .CO(n3262));
    SB_DFF BRAM_ADDR__i6 (.Q(TX_ADDR[6]), .C(ADV_CLK_c), .D(n22));   // ../tx.v(68[12] 94[8])
    SB_LUT4 i1603_4_lut (.I0(n133[4]), .I1(ADV_VSYNC_c), .I2(n102[4]), 
            .I3(n3787), .O(n24));   // ../tx.v(68[12] 94[8])
    defparam i1603_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESR Y_DELTA_PATTERN_i88 (.Q(Y_DELTA_PATTERN[88]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[89]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i5 (.Q(TX_ADDR[5]), .C(ADV_CLK_c), .D(n23));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i4 (.Q(TX_ADDR[4]), .C(ADV_CLK_c), .D(n24));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i3 (.Q(TX_ADDR[3]), .C(ADV_CLK_c), .D(n25));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_12_i6_3_lut (.I0(ADDR_Y_COMPONENT[5]), .I1(TX_ADDR[5]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[5]));   // ../tx.v(83[30:81])
    defparam mux_12_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_13_5_lut (.I0(GND_net), .I1(TX_ADDR[3]), .I2(GND_net), 
            .I3(n3260), .O(n118[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i6_3_lut (.I0(TX_ADDR[5]), .I1(n118[5]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[5]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1604_4_lut (.I0(n133[5]), .I1(ADV_VSYNC_c), .I2(n102[5]), 
            .I3(n3787), .O(n23));   // ../tx.v(68[12] 94[8])
    defparam i1604_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS Y_DELTA_PATTERN_i87 (.Q(Y_DELTA_PATTERN[87]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[88]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i86 (.Q(Y_DELTA_PATTERN[86]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[87]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_12_i7_3_lut (.I0(ADDR_Y_COMPONENT[6]), .I1(TX_ADDR[6]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[6]));   // ../tx.v(83[30:81])
    defparam mux_12_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS Y_DELTA_PATTERN_i85 (.Q(Y_DELTA_PATTERN[85]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[86]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i84 (.Q(Y_DELTA_PATTERN[84]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[85]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i83 (.Q(Y_DELTA_PATTERN[83]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[84]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i2 (.Q(TX_ADDR[2]), .C(ADV_CLK_c), .D(n26));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i82 (.Q(Y_DELTA_PATTERN[82]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[83]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFF BRAM_ADDR__i1 (.Q(TX_ADDR[1]), .C(ADV_CLK_c), .D(n27));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i81 (.Q(Y_DELTA_PATTERN[81]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[82]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i80 (.Q(Y_DELTA_PATTERN[80]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[81]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i79 (.Q(Y_DELTA_PATTERN[79]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[80]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_14_i7_3_lut (.I0(TX_ADDR[6]), .I1(n118[6]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[6]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR Y_DELTA_PATTERN_i78 (.Q(Y_DELTA_PATTERN[78]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[79]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_LUT4 i1605_4_lut (.I0(n133[6]), .I1(ADV_VSYNC_c), .I2(n102[6]), 
            .I3(n3787), .O(n22));   // ../tx.v(68[12] 94[8])
    defparam i1605_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS Y_DELTA_PATTERN_i97 (.Q(Y_DELTA_PATTERN[97]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[98]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i77 (.Q(Y_DELTA_PATTERN[77]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[78]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i96 (.Q(Y_DELTA_PATTERN[96]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[97]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_12_i8_3_lut (.I0(ADDR_Y_COMPONENT[7]), .I1(TX_ADDR[7]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[7]));   // ../tx.v(83[30:81])
    defparam mux_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS Y_DELTA_PATTERN_i76 (.Q(Y_DELTA_PATTERN[76]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[77]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i75 (.Q(Y_DELTA_PATTERN[75]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[76]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i74 (.Q(Y_DELTA_PATTERN[74]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[75]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i73 (.Q(Y_DELTA_PATTERN[73]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[74]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i72 (.Q(Y_DELTA_PATTERN[72]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[73]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i71 (.Q(Y_DELTA_PATTERN[71]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[72]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i70 (.Q(Y_DELTA_PATTERN[70]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[71]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i69 (.Q(Y_DELTA_PATTERN[69]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[70]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i68 (.Q(Y_DELTA_PATTERN[68]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[69]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i67 (.Q(Y_DELTA_PATTERN[67]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[68]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i66 (.Q(Y_DELTA_PATTERN[66]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[67]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i65 (.Q(Y_DELTA_PATTERN[65]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[66]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i64 (.Q(Y_DELTA_PATTERN[64]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[65]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i63 (.Q(Y_DELTA_PATTERN[63]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[64]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i62 (.Q(Y_DELTA_PATTERN[62]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[63]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i61 (.Q(Y_DELTA_PATTERN[61]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[62]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i60 (.Q(Y_DELTA_PATTERN[60]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[61]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i59 (.Q(Y_DELTA_PATTERN[59]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[60]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i58 (.Q(Y_DELTA_PATTERN[58]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[59]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i57 (.Q(Y_DELTA_PATTERN[57]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[58]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i56 (.Q(Y_DELTA_PATTERN[56]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[57]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i55 (.Q(Y_DELTA_PATTERN[55]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[56]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i54 (.Q(Y_DELTA_PATTERN[54]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[55]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i53 (.Q(Y_DELTA_PATTERN[53]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[54]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i52 (.Q(Y_DELTA_PATTERN[52]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[53]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i51 (.Q(Y_DELTA_PATTERN[51]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[52]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i50 (.Q(Y_DELTA_PATTERN[50]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[51]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i49 (.Q(Y_DELTA_PATTERN[49]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[50]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i48 (.Q(Y_DELTA_PATTERN[48]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[49]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i47 (.Q(Y_DELTA_PATTERN[47]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[48]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i46 (.Q(Y_DELTA_PATTERN[46]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[47]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i45 (.Q(Y_DELTA_PATTERN[45]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[46]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i44 (.Q(Y_DELTA_PATTERN[44]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[45]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i43 (.Q(Y_DELTA_PATTERN[43]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[44]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i42 (.Q(Y_DELTA_PATTERN[42]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[43]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i41 (.Q(Y_DELTA_PATTERN[41]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[42]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i40 (.Q(Y_DELTA_PATTERN[40]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[41]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i39 (.Q(Y_DELTA_PATTERN[39]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[40]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i38 (.Q(Y_DELTA_PATTERN[38]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[39]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i37 (.Q(Y_DELTA_PATTERN[37]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[38]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i36 (.Q(Y_DELTA_PATTERN[36]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[37]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i35 (.Q(Y_DELTA_PATTERN[35]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[36]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i34 (.Q(Y_DELTA_PATTERN[34]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[35]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i33 (.Q(Y_DELTA_PATTERN[33]), .C(ADV_CLK_c), 
            .E(n3798), .D(Y_DELTA_PATTERN[34]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i32 (.Q(Y_DELTA_PATTERN[32]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[33]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i31 (.Q(Y_DELTA_PATTERN[31]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[32]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i30 (.Q(Y_DELTA_PATTERN[30]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[31]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i29 (.Q(Y_DELTA_PATTERN[29]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[30]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i28 (.Q(Y_DELTA_PATTERN[28]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[29]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i27 (.Q(Y_DELTA_PATTERN[27]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[28]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i26 (.Q(Y_DELTA_PATTERN[26]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[27]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i25 (.Q(Y_DELTA_PATTERN[25]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[26]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i24 (.Q(Y_DELTA_PATTERN[24]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[25]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i23 (.Q(Y_DELTA_PATTERN[23]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[24]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i22 (.Q(Y_DELTA_PATTERN[22]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[23]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i21 (.Q(Y_DELTA_PATTERN[21]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[22]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i20 (.Q(Y_DELTA_PATTERN[20]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[21]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i19 (.Q(Y_DELTA_PATTERN[19]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[20]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i18 (.Q(Y_DELTA_PATTERN[18]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[19]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i17 (.Q(Y_DELTA_PATTERN[17]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[18]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i16 (.Q(Y_DELTA_PATTERN[16]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[17]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i15 (.Q(Y_DELTA_PATTERN[15]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[16]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i14 (.Q(Y_DELTA_PATTERN[14]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[15]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i13 (.Q(Y_DELTA_PATTERN[13]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[14]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i12 (.Q(Y_DELTA_PATTERN[12]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[13]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i11 (.Q(Y_DELTA_PATTERN[11]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[12]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i10 (.Q(Y_DELTA_PATTERN[10]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[11]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i9 (.Q(Y_DELTA_PATTERN[9]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[10]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i8 (.Q(Y_DELTA_PATTERN[8]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[9]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i7 (.Q(Y_DELTA_PATTERN[7]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[8]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i6 (.Q(Y_DELTA_PATTERN[6]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[7]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i5 (.Q(Y_DELTA_PATTERN[5]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[6]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i4 (.Q(Y_DELTA_PATTERN[4]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[5]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i3 (.Q(Y_DELTA_PATTERN[3]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[4]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_LUT4 mux_14_i8_3_lut (.I0(TX_ADDR[7]), .I1(n118[7]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[7]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1606_4_lut (.I0(n133[7]), .I1(ADV_VSYNC_c), .I2(n102[7]), 
            .I3(n3787), .O(n21));   // ../tx.v(68[12] 94[8])
    defparam i1606_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i9_3_lut (.I0(ADDR_Y_COMPONENT[8]), .I1(TX_ADDR[8]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[8]));   // ../tx.v(83[30:81])
    defparam mux_12_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i9_3_lut (.I0(TX_ADDR[8]), .I1(n118[8]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[8]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1607_4_lut (.I0(n133[8]), .I1(ADV_VSYNC_c), .I2(n102[8]), 
            .I3(n3787), .O(n20));   // ../tx.v(68[12] 94[8])
    defparam i1607_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i10_3_lut (.I0(ADDR_Y_COMPONENT[9]), .I1(TX_ADDR[9]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[9]));   // ../tx.v(83[30:81])
    defparam mux_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i10_3_lut (.I0(TX_ADDR[9]), .I1(n118[9]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[9]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1608_4_lut (.I0(n133[9]), .I1(ADV_VSYNC_c), .I2(n102[9]), 
            .I3(n3787), .O(n19));   // ../tx.v(68[12] 94[8])
    defparam i1608_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_18_i14_3_lut (.I0(n118[13]), .I1(ADDR_Y_COMPONENT[13]), 
            .I2(n3787), .I3(GND_net), .O(BRAM_ADDR_13__N_282[13]));   // ../tx.v(85[22] 90[16])
    defparam mux_18_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_18_i13_3_lut (.I0(n118[12]), .I1(ADDR_Y_COMPONENT[12]), 
            .I2(n3787), .I3(GND_net), .O(BRAM_ADDR_13__N_282[12]));   // ../tx.v(85[22] 90[16])
    defparam mux_18_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_12_i11_3_lut (.I0(ADDR_Y_COMPONENT[10]), .I1(TX_ADDR[10]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n102[10]));   // ../tx.v(83[30:81])
    defparam mux_12_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i11_3_lut (.I0(TX_ADDR[10]), .I1(n118[10]), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n133[10]));   // ../tx.v(86[17] 89[20])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1609_4_lut (.I0(n133[10]), .I1(ADV_VSYNC_c), .I2(n102[10]), 
            .I3(n3787), .O(n18));   // ../tx.v(68[12] 94[8])
    defparam i1609_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_3_lut (.I0(n3787), .I1(ADV_VSYNC_c), .I2(Y_DELTA_PATTERN[0]), 
            .I3(GND_net), .O(n2061));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1613_4_lut (.I0(ADV_VSYNC_c), .I1(VGA_VISIBLE), .I2(Y_DELTA_PATTERN[0]), 
            .I3(n3787), .O(n2039));
    defparam i1613_4_lut.LUT_INIT = 16'hafee;
    SB_LUT4 mux_18_i12_3_lut (.I0(n118[11]), .I1(ADDR_Y_COMPONENT[11]), 
            .I2(n3787), .I3(GND_net), .O(BRAM_ADDR_13__N_282[11]));   // ../tx.v(85[22] 90[16])
    defparam mux_18_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(n3787), .I1(ADV_VSYNC_c), .I2(VGA_VISIBLE), 
            .I3(GND_net), .O(n2093));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_13_14 (.CI(n3269), .I0(\TX_ADDR[12] ), .I1(GND_net), 
            .CO(n3270));
    SB_LUT4 add_13_13_lut (.I0(GND_net), .I1(\TX_ADDR[11] ), .I2(GND_net), 
            .I3(n3268), .O(n118[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_5 (.CI(n3260), .I0(TX_ADDR[3]), .I1(GND_net), .CO(n3261));
    SB_CARRY add_13_13 (.CI(n3268), .I0(\TX_ADDR[11] ), .I1(GND_net), 
            .CO(n3269));
    SB_LUT4 add_13_12_lut (.I0(GND_net), .I1(TX_ADDR[10]), .I2(GND_net), 
            .I3(n3267), .O(n118[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_4_lut (.I0(GND_net), .I1(TX_ADDR[2]), .I2(GND_net), 
            .I3(n3259), .O(n118[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_12 (.CI(n3267), .I0(TX_ADDR[10]), .I1(GND_net), .CO(n3268));
    SB_CARRY add_13_4 (.CI(n3259), .I0(TX_ADDR[2]), .I1(GND_net), .CO(n3260));
    SB_LUT4 add_13_3_lut (.I0(GND_net), .I1(TX_ADDR[1]), .I2(GND_net), 
            .I3(n3258), .O(n118[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_3 (.CI(n3258), .I0(TX_ADDR[1]), .I1(GND_net), .CO(n3259));
    SB_LUT4 add_13_11_lut (.I0(GND_net), .I1(TX_ADDR[9]), .I2(GND_net), 
            .I3(n3266), .O(n118[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_11 (.CI(n3266), .I0(TX_ADDR[9]), .I1(GND_net), .CO(n3267));
    SB_LUT4 add_13_10_lut (.I0(GND_net), .I1(TX_ADDR[8]), .I2(GND_net), 
            .I3(n3265), .O(n118[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_2_lut (.I0(GND_net), .I1(TX_ADDR[0]), .I2(X_DELTA_PATTERN[0]), 
            .I3(GND_net), .O(n118[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_2 (.CI(GND_net), .I0(TX_ADDR[0]), .I1(X_DELTA_PATTERN[0]), 
            .CO(n3258));
    SB_CARRY add_13_10 (.CI(n3265), .I0(TX_ADDR[8]), .I1(GND_net), .CO(n3266));
    SB_LUT4 add_13_9_lut (.I0(GND_net), .I1(TX_ADDR[7]), .I2(GND_net), 
            .I3(n3264), .O(n118[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_9 (.CI(n3264), .I0(TX_ADDR[7]), .I1(GND_net), .CO(n3265));
    SB_LUT4 add_13_8_lut (.I0(GND_net), .I1(TX_ADDR[6]), .I2(GND_net), 
            .I3(n3263), .O(n118[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_8 (.CI(n3263), .I0(TX_ADDR[6]), .I1(GND_net), .CO(n3264));
    SB_LUT4 add_13_7_lut (.I0(GND_net), .I1(TX_ADDR[5]), .I2(GND_net), 
            .I3(n3262), .O(n118[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_7 (.CI(n3262), .I0(TX_ADDR[5]), .I1(GND_net), .CO(n3263));
    SB_DFFESS Y_DELTA_PATTERN_i0 (.Q(Y_DELTA_PATTERN[0]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[1]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i0 (.Q(X_DELTA_PATTERN[0]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[1]), .S(n2147));   // ../tx.v(68[12] 94[8])
    SB_DFFESR BRAM_ADDR__rep_1_i0 (.Q(\TX_ADDR[11] ), .C(ADV_CLK_c), .E(n2039), 
            .D(BRAM_ADDR_13__N_282[11]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i0 (.Q(ADDR_Y_COMPONENT[0]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[0]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFSR VGA_R__i1 (.Q(n1798), .C(ADV_CLK_c), .D(TX_DATA[0]), .R(n2354));   // ../tx.v(68[12] 94[8])
    SB_DFFESR Y_DELTA_PATTERN_i2 (.Q(Y_DELTA_PATTERN[2]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[3]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i1 (.Q(Y_DELTA_PATTERN[1]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[2]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i15 (.Q(X_DELTA_PATTERN[15]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[0]), .S(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESR X_DELTA_PATTERN_i14 (.Q(X_DELTA_PATTERN[14]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[15]), .R(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i13 (.Q(X_DELTA_PATTERN[13]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[14]), .S(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESR X_DELTA_PATTERN_i12 (.Q(X_DELTA_PATTERN[12]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[13]), .R(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i11 (.Q(X_DELTA_PATTERN[11]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[12]), .S(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESR X_DELTA_PATTERN_i10 (.Q(X_DELTA_PATTERN[10]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[11]), .R(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i9 (.Q(X_DELTA_PATTERN[9]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[10]), .S(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESR X_DELTA_PATTERN_i8 (.Q(X_DELTA_PATTERN[8]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[9]), .R(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i7 (.Q(X_DELTA_PATTERN[7]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[8]), .S(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i6 (.Q(X_DELTA_PATTERN[6]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[7]), .S(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESR X_DELTA_PATTERN_i5 (.Q(X_DELTA_PATTERN[5]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[6]), .R(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i4 (.Q(X_DELTA_PATTERN[4]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[5]), .S(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESR X_DELTA_PATTERN_i3 (.Q(X_DELTA_PATTERN[3]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[4]), .R(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESS X_DELTA_PATTERN_i2 (.Q(X_DELTA_PATTERN[2]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[3]), .S(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESR X_DELTA_PATTERN_i1 (.Q(X_DELTA_PATTERN[1]), .C(ADV_CLK_c), 
            .E(n2093), .D(X_DELTA_PATTERN[2]), .R(n3797));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i13 (.Q(ADDR_Y_COMPONENT[13]), .C(ADV_CLK_c), 
            .E(n2061), .D(\TX_ADDR[13] ), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i12 (.Q(ADDR_Y_COMPONENT[12]), .C(ADV_CLK_c), 
            .E(n2061), .D(\TX_ADDR[12] ), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i11 (.Q(ADDR_Y_COMPONENT[11]), .C(ADV_CLK_c), 
            .E(n2061), .D(\TX_ADDR[11] ), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i10 (.Q(ADDR_Y_COMPONENT[10]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[10]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i9 (.Q(ADDR_Y_COMPONENT[9]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[9]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i8 (.Q(ADDR_Y_COMPONENT[8]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[8]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i7 (.Q(ADDR_Y_COMPONENT[7]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[7]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i6 (.Q(ADDR_Y_COMPONENT[6]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[6]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i5 (.Q(ADDR_Y_COMPONENT[5]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[5]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i4 (.Q(ADDR_Y_COMPONENT[4]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[4]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i3 (.Q(ADDR_Y_COMPONENT[3]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[3]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i2 (.Q(ADDR_Y_COMPONENT[2]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[2]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR ADDR_Y_COMPONENT__i1 (.Q(ADDR_Y_COMPONENT[1]), .C(ADV_CLK_c), 
            .E(n2061), .D(TX_ADDR[1]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR BRAM_ADDR__i12 (.Q(\TX_ADDR[12] ), .C(ADV_CLK_c), .E(n2039), 
            .D(BRAM_ADDR_13__N_282[12]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESR BRAM_ADDR__i13 (.Q(\TX_ADDR[13] ), .C(ADV_CLK_c), .E(n2039), 
            .D(BRAM_ADDR_13__N_282[13]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_LUT4 i246_2_lut_4_lut (.I0(ADV_HSYNC_c), .I1(VGA_VISIBLE_Y), .I2(old_VGA_HS), 
            .I3(ADV_VSYNC_c), .O(n2147));   // ../tx.v(80[16:63])
    defparam i246_2_lut_4_lut.LUT_INIT = 16'hff40;
    SB_LUT4 i2_3_lut_rep_20 (.I0(ADV_HSYNC_c), .I1(VGA_VISIBLE_Y), .I2(old_VGA_HS), 
            .I3(GND_net), .O(n3787));   // ../tx.v(80[16:63])
    defparam i2_3_lut_rep_20.LUT_INIT = 16'h4040;
    SB_LUT4 i246_2_lut_4_lut_rep_31 (.I0(ADV_HSYNC_c), .I1(VGA_VISIBLE_Y), 
            .I2(old_VGA_HS), .I3(ADV_VSYNC_c), .O(n3798));   // ../tx.v(80[16:63])
    defparam i246_2_lut_4_lut_rep_31.LUT_INIT = 16'hff40;
    SB_LUT4 i246_2_lut_4_lut_rep_30 (.I0(ADV_HSYNC_c), .I1(VGA_VISIBLE_Y), 
            .I2(old_VGA_HS), .I3(ADV_VSYNC_c), .O(n3797));   // ../tx.v(80[16:63])
    defparam i246_2_lut_4_lut_rep_30.LUT_INIT = 16'hff40;
    SB_DFFESR Y_DELTA_PATTERN_i99 (.Q(Y_DELTA_PATTERN[99]), .C(ADV_CLK_c), 
            .E(n3797), .D(Y_DELTA_PATTERN[0]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    SB_DFFESS Y_DELTA_PATTERN_i95 (.Q(Y_DELTA_PATTERN[95]), .C(ADV_CLK_c), 
            .E(n2147), .D(Y_DELTA_PATTERN[96]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 94[8])
    VGA_CONTROL video_signal_controller (.GND_net(GND_net), .ADV_CLK_c(ADV_CLK_c), 
            .VCC_net(VCC_net), .VGA_VISIBLE_Y(VGA_VISIBLE_Y), .VGA_VISIBLE(VGA_VISIBLE), 
            .ADV_HSYNC_c(ADV_HSYNC_c), .ADV_VSYNC_c(ADV_VSYNC_c), .RX_TX_SYNC_BUFF(RX_TX_SYNC_BUFF), 
            .n2354(n2354)) /* synthesis syn_module_defined=1 */ ;   // ../tx.v(44[17] 58[67])
    
endmodule
//
// Verilog Description of module VGA_CONTROL
//

module VGA_CONTROL (GND_net, ADV_CLK_c, VCC_net, VGA_VISIBLE_Y, VGA_VISIBLE, 
            ADV_HSYNC_c, ADV_VSYNC_c, RX_TX_SYNC_BUFF, n2354) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input ADV_CLK_c;
    input VCC_net;
    output VGA_VISIBLE_Y;
    output VGA_VISIBLE;
    output ADV_HSYNC_c;
    output ADV_VSYNC_c;
    input RX_TX_SYNC_BUFF;
    output n2354;
    
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    wire [11:0]n229;
    wire [11:0]VGA_X;   // ../vga_control.v(54[16:21])
    
    wire n3285, n3286, n3789, n1983, n3467, n18;
    wire [11:0]n249;
    
    wire n2010;
    wire [11:0]VGA_Y;   // ../vga_control.v(54[23:28])
    
    wire n2361, n3284, n3291, n3292, n3279, n7, VGA_VISIBLE_N_578, 
        n3486, VGA_VISIBLE_N_573, VGA_VISIBLE_Y_N_581, n3485, n3299, 
        VGA_HS_N_567, VGA_VS_N_570, n3300, n2, n3577, n3283, n3290, 
        n3785, n3786, n7_adj_615, n8, n2886, n2926, n3794, n3626, 
        n3614, n18_adj_616, n3632, n2876, n3788, n4, n4_adj_617, 
        n3618, n3282, n3294, n3295, n3293, n3296, n3297, n3298, 
        n3289, n3281, n3288, n3280, n3287;
    
    SB_LUT4 add_35_9_lut (.I0(GND_net), .I1(VGA_X[7]), .I2(GND_net), .I3(n3285), 
            .O(n229[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_35_9 (.CI(n3285), .I0(VGA_X[7]), .I1(GND_net), .CO(n3286));
    SB_LUT4 i483_4_lut (.I0(n3789), .I1(VGA_X[8]), .I2(n1983), .I3(n3467), 
            .O(n18));
    defparam i483_4_lut.LUT_INIT = 16'hc8c0;
    SB_DFFESR VGA_Y_i8 (.Q(VGA_Y[8]), .C(ADV_CLK_c), .E(n2010), .D(n249[8]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_LUT4 add_35_8_lut (.I0(GND_net), .I1(VGA_X[6]), .I2(GND_net), .I3(n3284), 
            .O(n229[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_42_4 (.CI(n3291), .I0(VGA_Y[2]), .I1(GND_net), .CO(n3292));
    SB_CARRY add_35_2 (.CI(VCC_net), .I0(VGA_X[0]), .I1(GND_net), .CO(n3279));
    SB_CARRY add_35_8 (.CI(n3284), .I0(VGA_X[6]), .I1(GND_net), .CO(n3285));
    SB_LUT4 i4_4_lut (.I0(n7), .I1(VGA_VISIBLE_N_578), .I2(VGA_X[11]), 
            .I3(n3486), .O(VGA_VISIBLE_N_573));
    defparam i4_4_lut.LUT_INIT = 16'h0008;
    SB_DFF VGA_VISIBLE_Y_64 (.Q(VGA_VISIBLE_Y), .C(ADV_CLK_c), .D(VGA_VISIBLE_Y_N_581));   // ../vga_control.v(69[12] 98[8])
    SB_LUT4 i1_2_lut (.I0(VGA_Y[10]), .I1(VGA_Y[11]), .I2(GND_net), .I3(GND_net), 
            .O(n3485));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_42_12_lut (.I0(GND_net), .I1(VGA_Y[10]), .I2(GND_net), 
            .I3(n3299), .O(n249[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF VGA_VISIBLE_65 (.Q(VGA_VISIBLE), .C(ADV_CLK_c), .D(VGA_VISIBLE_N_573));   // ../vga_control.v(69[12] 98[8])
    SB_DFF VGA_HS_66 (.Q(ADV_HSYNC_c), .C(ADV_CLK_c), .D(VGA_HS_N_567));   // ../vga_control.v(69[12] 98[8])
    SB_DFF VGA_VS_67 (.Q(ADV_VSYNC_c), .C(ADV_CLK_c), .D(VGA_VS_N_570));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i0 (.Q(VGA_X[0]), .C(ADV_CLK_c), .D(n229[0]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i1 (.Q(VGA_X[1]), .C(ADV_CLK_c), .D(n229[1]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i2 (.Q(VGA_X[2]), .C(ADV_CLK_c), .D(n229[2]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i3 (.Q(VGA_X[3]), .C(ADV_CLK_c), .D(n229[3]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i4 (.Q(VGA_X[4]), .C(ADV_CLK_c), .D(n229[4]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i5 (.Q(VGA_X[5]), .C(ADV_CLK_c), .D(n229[5]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i6 (.Q(VGA_X[6]), .C(ADV_CLK_c), .D(n229[6]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i7 (.Q(VGA_X[7]), .C(ADV_CLK_c), .D(n229[7]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i8 (.Q(VGA_X[8]), .C(ADV_CLK_c), .D(n229[8]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i9 (.Q(VGA_X[9]), .C(ADV_CLK_c), .D(n229[9]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i10 (.Q(VGA_X[10]), .C(ADV_CLK_c), .D(n229[10]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_DFFSR VGA_X_i11 (.Q(VGA_X[11]), .C(ADV_CLK_c), .D(n229[11]), .R(n2010));   // ../vga_control.v(69[12] 98[8])
    SB_CARRY add_42_12 (.CI(n3299), .I0(VGA_Y[10]), .I1(GND_net), .CO(n3300));
    SB_LUT4 i2_4_lut (.I0(VGA_Y[6]), .I1(VGA_Y[5]), .I2(VGA_Y[4]), .I3(n2), 
            .O(n3577));   // ../vga_control.v(54[23:28])
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 add_35_7_lut (.I0(GND_net), .I1(VGA_X[5]), .I2(GND_net), .I3(n3283), 
            .O(n229[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR VGA_Y_i7 (.Q(VGA_Y[7]), .C(ADV_CLK_c), .E(n2010), .D(n249[7]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_LUT4 add_42_3_lut (.I0(GND_net), .I1(VGA_Y[1]), .I2(GND_net), .I3(n3290), 
            .O(n249[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR VGA_Y_i6 (.Q(VGA_Y[6]), .C(ADV_CLK_c), .E(n2010), .D(n249[6]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_LUT4 i1_2_lut_adj_23 (.I0(VGA_X[4]), .I1(VGA_X[3]), .I2(GND_net), 
            .I3(GND_net), .O(n3467));
    defparam i1_2_lut_adj_23.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n3577), .I1(n3485), .I2(VGA_Y[9]), .I3(n3785), 
            .O(n3486));
    defparam i1_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_4_lut (.I0(VGA_X[11]), .I1(VGA_X[10]), .I2(VGA_X[9]), 
            .I3(n18), .O(n7));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h333e;
    SB_DFFESR VGA_Y_i11 (.Q(VGA_Y[11]), .C(ADV_CLK_c), .E(n2010), .D(n249[11]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_DFFESR VGA_Y_i10 (.Q(VGA_Y[10]), .C(ADV_CLK_c), .E(n2010), .D(n249[10]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_LUT4 i1_4_lut_adj_24 (.I0(n3485), .I1(VGA_Y[4]), .I2(n3786), .I3(VGA_Y[3]), 
            .O(n7_adj_615));
    defparam i1_4_lut_adj_24.LUT_INIT = 16'heeea;
    SB_DFFESR VGA_Y_i9 (.Q(VGA_Y[9]), .C(ADV_CLK_c), .E(n2010), .D(n249[9]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_LUT4 i1136_2_lut (.I0(n2010), .I1(RX_TX_SYNC_BUFF), .I2(GND_net), 
            .I3(GND_net), .O(n2361));   // ../vga_control.v(69[12] 98[8])
    defparam i1136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(VGA_Y[6]), .I1(n7_adj_615), .I2(VGA_Y[5]), .I3(n8), 
            .O(VGA_VISIBLE_N_578));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 VGA_VISIBLE_N_578_I_0_2_lut (.I0(VGA_VISIBLE_N_578), .I1(n3486), 
            .I2(GND_net), .I3(GND_net), .O(VGA_VISIBLE_Y_N_581));   // ../vga_control.v(72[26:101])
    defparam VGA_VISIBLE_N_578_I_0_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1693_4_lut (.I0(n2886), .I1(VGA_X[8]), .I2(n1983), .I3(n3467), 
            .O(n2926));
    defparam i1693_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i1699_4_lut (.I0(n2926), .I1(VGA_X[11]), .I2(VGA_X[10]), .I3(VGA_X[9]), 
            .O(n2010));
    defparam i1699_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_3_lut_rep_27 (.I0(VGA_X[11]), .I1(VGA_X[10]), .I2(VGA_X[9]), 
            .I3(GND_net), .O(n3794));
    defparam i2_3_lut_rep_27.LUT_INIT = 16'hfefe;
    SB_LUT4 i1120_1_lut (.I0(VGA_VISIBLE), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2354));   // ../vga_control.v(69[12] 98[8])
    defparam i1120_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2300_2_lut (.I0(VGA_Y[4]), .I1(VGA_Y[8]), .I2(GND_net), .I3(GND_net), 
            .O(n3626));
    defparam i2300_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2288_2_lut (.I0(VGA_Y[9]), .I1(VGA_Y[6]), .I2(GND_net), .I3(GND_net), 
            .O(n3614));
    defparam i2288_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut (.I0(VGA_Y[1]), .I1(n3626), .I2(VGA_Y[3]), .I3(VGA_Y[0]), 
            .O(n18_adj_616));
    defparam i7_4_lut.LUT_INIT = 16'h0302;
    SB_LUT4 i2306_4_lut (.I0(VGA_Y[7]), .I1(VGA_Y[5]), .I2(VGA_Y[11]), 
            .I3(VGA_Y[2]), .O(n3632));
    defparam i2306_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n3632), .I1(VGA_Y[10]), .I2(n18_adj_616), .I3(n3614), 
            .O(VGA_VS_N_570));
    defparam i10_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1643_2_lut (.I0(VGA_X[0]), .I1(VGA_X[1]), .I2(GND_net), .I3(GND_net), 
            .O(n2876));
    defparam i1643_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_25 (.I0(n3788), .I1(VGA_X[2]), .I2(VGA_X[3]), 
            .I3(n2876), .O(n4));   // ../vga_control.v(75[49:87])
    defparam i1_4_lut_adj_25.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_26 (.I0(VGA_X[7]), .I1(VGA_X[3]), .I2(VGA_X[5]), 
            .I3(VGA_X[4]), .O(n4_adj_617));
    defparam i1_4_lut_adj_26.LUT_INIT = 16'hfaea;
    SB_LUT4 i2292_4_lut (.I0(VGA_X[4]), .I1(n3794), .I2(VGA_X[7]), .I3(n4), 
            .O(n3618));
    defparam i2292_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2357_4_lut (.I0(VGA_X[6]), .I1(n3618), .I2(VGA_X[8]), .I3(n4_adj_617), 
            .O(VGA_HS_N_567));   // ../vga_control.v(75[19:88])
    defparam i2357_4_lut.LUT_INIT = 16'hfcfd;
    SB_CARRY add_35_7 (.CI(n3283), .I0(VGA_X[5]), .I1(GND_net), .CO(n3284));
    SB_LUT4 add_35_6_lut (.I0(GND_net), .I1(VGA_X[4]), .I2(GND_net), .I3(n3282), 
            .O(n229[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_42_3 (.CI(n3290), .I0(VGA_Y[1]), .I1(GND_net), .CO(n3291));
    SB_CARRY add_42_7 (.CI(n3294), .I0(VGA_Y[5]), .I1(GND_net), .CO(n3295));
    SB_LUT4 add_42_2_lut (.I0(GND_net), .I1(VGA_Y[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n249[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_35_6 (.CI(n3282), .I0(VGA_X[4]), .I1(GND_net), .CO(n3283));
    SB_CARRY add_42_2 (.CI(VCC_net), .I0(VGA_Y[0]), .I1(GND_net), .CO(n3290));
    SB_LUT4 add_42_6_lut (.I0(GND_net), .I1(VGA_Y[4]), .I2(GND_net), .I3(n3293), 
            .O(n249[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_42_9 (.CI(n3296), .I0(VGA_Y[7]), .I1(GND_net), .CO(n3297));
    SB_LUT4 add_42_11_lut (.I0(GND_net), .I1(VGA_Y[9]), .I2(GND_net), 
            .I3(n3298), .O(n249[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_35_13_lut (.I0(GND_net), .I1(VGA_X[11]), .I2(GND_net), 
            .I3(n3289), .O(n229[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_42_6 (.CI(n3293), .I0(VGA_Y[4]), .I1(GND_net), .CO(n3294));
    SB_LUT4 add_42_8_lut (.I0(GND_net), .I1(VGA_Y[6]), .I2(GND_net), .I3(n3295), 
            .O(n249[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_35_5_lut (.I0(GND_net), .I1(VGA_X[3]), .I2(GND_net), .I3(n3281), 
            .O(n229[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_42_11 (.CI(n3298), .I0(VGA_Y[9]), .I1(GND_net), .CO(n3299));
    SB_CARRY add_35_5 (.CI(n3281), .I0(VGA_X[3]), .I1(GND_net), .CO(n3282));
    SB_LUT4 add_35_12_lut (.I0(GND_net), .I1(VGA_X[10]), .I2(GND_net), 
            .I3(n3288), .O(n229[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_42_5_lut (.I0(GND_net), .I1(VGA_Y[3]), .I2(GND_net), .I3(n3292), 
            .O(n249[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_42_8 (.CI(n3295), .I0(VGA_Y[6]), .I1(GND_net), .CO(n3296));
    SB_LUT4 add_42_10_lut (.I0(GND_net), .I1(VGA_Y[8]), .I2(GND_net), 
            .I3(n3297), .O(n249[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_35_4_lut (.I0(GND_net), .I1(VGA_X[2]), .I2(GND_net), .I3(n3280), 
            .O(n229[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_35_12 (.CI(n3288), .I0(VGA_X[10]), .I1(GND_net), .CO(n3289));
    SB_CARRY add_35_4 (.CI(n3280), .I0(VGA_X[2]), .I1(GND_net), .CO(n3281));
    SB_LUT4 add_35_11_lut (.I0(GND_net), .I1(VGA_X[9]), .I2(GND_net), 
            .I3(n3287), .O(n229[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_42_5 (.CI(n3292), .I0(VGA_Y[3]), .I1(GND_net), .CO(n3293));
    SB_CARRY add_35_11 (.CI(n3287), .I0(VGA_X[9]), .I1(GND_net), .CO(n3288));
    SB_LUT4 add_42_4_lut (.I0(GND_net), .I1(VGA_Y[2]), .I2(GND_net), .I3(n3291), 
            .O(n249[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_42_7_lut (.I0(GND_net), .I1(VGA_Y[5]), .I2(GND_net), .I3(n3294), 
            .O(n249[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_42_10 (.CI(n3297), .I0(VGA_Y[8]), .I1(GND_net), .CO(n3298));
    SB_LUT4 add_35_3_lut (.I0(GND_net), .I1(VGA_X[1]), .I2(GND_net), .I3(n3279), 
            .O(n229[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_35_3 (.CI(n3279), .I0(VGA_X[1]), .I1(GND_net), .CO(n3280));
    SB_LUT4 add_35_10_lut (.I0(GND_net), .I1(VGA_X[8]), .I2(GND_net), 
            .I3(n3286), .O(n229[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_42_9_lut (.I0(GND_net), .I1(VGA_Y[7]), .I2(GND_net), .I3(n3296), 
            .O(n249[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_42_13_lut (.I0(GND_net), .I1(VGA_Y[11]), .I2(GND_net), 
            .I3(n3300), .O(n249[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_42_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR VGA_Y_i5 (.Q(VGA_Y[5]), .C(ADV_CLK_c), .E(n2010), .D(n249[5]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_DFFESR VGA_Y_i4 (.Q(VGA_Y[4]), .C(ADV_CLK_c), .E(n2010), .D(n249[4]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_DFFESR VGA_Y_i3 (.Q(VGA_Y[3]), .C(ADV_CLK_c), .E(n2010), .D(n249[3]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_DFFESR VGA_Y_i2 (.Q(VGA_Y[2]), .C(ADV_CLK_c), .E(n2010), .D(n249[2]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_DFFESR VGA_Y_i1 (.Q(VGA_Y[1]), .C(ADV_CLK_c), .E(n2010), .D(n249[1]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_DFFESR VGA_Y_i0 (.Q(VGA_Y[0]), .C(ADV_CLK_c), .E(n2010), .D(n249[0]), 
            .R(n2361));   // ../vga_control.v(69[12] 98[8])
    SB_LUT4 add_35_2_lut (.I0(GND_net), .I1(VGA_X[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_35_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_35_10 (.CI(n3286), .I0(VGA_X[8]), .I1(GND_net), .CO(n3287));
    SB_LUT4 i1653_2_lut_3_lut (.I0(VGA_X[1]), .I1(VGA_X[2]), .I2(VGA_X[0]), 
            .I3(GND_net), .O(n2886));
    defparam i1653_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i495_2_lut_rep_22 (.I0(VGA_X[1]), .I1(VGA_X[2]), .I2(GND_net), 
            .I3(GND_net), .O(n3789));
    defparam i495_2_lut_rep_22.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut (.I0(VGA_X[5]), .I1(VGA_X[6]), .I2(VGA_X[7]), 
            .I3(GND_net), .O(n1983));   // ../vga_control.v(75[49:87])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_rep_21 (.I0(VGA_X[5]), .I1(VGA_X[6]), .I2(GND_net), 
            .I3(GND_net), .O(n3788));   // ../vga_control.v(75[49:87])
    defparam i1_2_lut_rep_21.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_27 (.I0(VGA_Y[2]), .I1(VGA_Y[1]), .I2(VGA_Y[3]), 
            .I3(GND_net), .O(n2));   // ../vga_control.v(54[23:28])
    defparam i1_2_lut_3_lut_adj_27.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_rep_19 (.I0(VGA_Y[2]), .I1(VGA_Y[1]), .I2(GND_net), 
            .I3(GND_net), .O(n3786));   // ../vga_control.v(54[23:28])
    defparam i1_2_lut_rep_19.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_3_lut (.I0(VGA_Y[7]), .I1(VGA_Y[8]), .I2(VGA_Y[9]), 
            .I3(GND_net), .O(n8));   // ../vga_control.v(54[23:28])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_rep_18 (.I0(VGA_Y[7]), .I1(VGA_Y[8]), .I2(GND_net), 
            .I3(GND_net), .O(n3785));   // ../vga_control.v(54[23:28])
    defparam i1_2_lut_rep_18.LUT_INIT = 16'heeee;
    
endmodule
//
// Verilog Description of module RX
//

module RX (RX_ADDR, GND_net, RX_WE, TVP_VSYNC_c, TVP_CLK_c, VCC_net, 
           TVP_HSYNC_c, RX_TX_SYNC, LED_c) /* synthesis syn_module_defined=1 */ ;
    output [13:0]RX_ADDR;
    input GND_net;
    output RX_WE;
    input TVP_VSYNC_c;
    input TVP_CLK_c;
    input VCC_net;
    input TVP_HSYNC_c;
    output RX_TX_SYNC;
    output LED_c;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    
    wire n3250, n3251, n3255, n3256;
    wire [13:0]n122;
    
    wire n2713, n2715, n3249, n2717, n3245, n3246, n2719, n2721, 
        n2723, n3795, n3793, n3254, n3247, n3248, n3253, n3252, 
        n3257, n2703, n2705, n2711, n2707, n2709;
    
    SB_CARRY add_12_8 (.CI(n3250), .I0(RX_ADDR[6]), .I1(GND_net), .CO(n3251));
    SB_CARRY add_12_13 (.CI(n3255), .I0(RX_ADDR[11]), .I1(GND_net), .CO(n3256));
    SB_LUT4 i1479_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[8]), 
            .I3(RX_ADDR[8]), .O(n2713));
    defparam i1479_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1481_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[9]), 
            .I3(RX_ADDR[9]), .O(n2715));
    defparam i1481_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(RX_ADDR[5]), .I2(GND_net), 
            .I3(n3249), .O(n122[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1483_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[10]), 
            .I3(RX_ADDR[10]), .O(n2717));
    defparam i1483_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_CARRY add_12_3 (.CI(n3245), .I0(RX_ADDR[1]), .I1(GND_net), .CO(n3246));
    SB_LUT4 i1485_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[0]), 
            .I3(RX_ADDR[0]), .O(n2719));
    defparam i1485_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1487_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[1]), 
            .I3(RX_ADDR[1]), .O(n2721));
    defparam i1487_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1489_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[2]), 
            .I3(RX_ADDR[2]), .O(n2723));
    defparam i1489_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i245_2_lut_rep_28 (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(GND_net), 
            .I3(GND_net), .O(n3795));
    defparam i245_2_lut_rep_28.LUT_INIT = 16'hbbbb;
    SB_DFFESR BRAM_ADDR__i11 (.Q(RX_ADDR[11]), .C(TVP_CLK_c), .E(n3795), 
            .D(n122[11]), .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_DFFESR BRAM_ADDR__i12 (.Q(RX_ADDR[12]), .C(TVP_CLK_c), .E(n3795), 
            .D(n122[12]), .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_DFFESR BRAM_ADDR__i13 (.Q(RX_ADDR[13]), .C(TVP_CLK_c), .E(n3795), 
            .D(n122[13]), .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(RX_ADDR[10]), .I2(GND_net), 
            .I3(n3254), .O(n122[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_5 (.CI(n3247), .I0(RX_ADDR[3]), .I1(GND_net), .CO(n3248));
    SB_CARRY add_12_7 (.CI(n3249), .I0(RX_ADDR[5]), .I1(GND_net), .CO(n3250));
    SB_CARRY add_12_12 (.CI(n3254), .I0(RX_ADDR[10]), .I1(GND_net), .CO(n3255));
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(RX_ADDR[2]), .I2(GND_net), 
            .I3(n3246), .O(n122[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(RX_ADDR[9]), .I2(GND_net), 
            .I3(n3253), .O(n122[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n3253), .I0(RX_ADDR[9]), .I1(GND_net), .CO(n3254));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(RX_ADDR[8]), .I2(GND_net), 
            .I3(n3252), .O(n122[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_10 (.CI(n3252), .I0(RX_ADDR[8]), .I1(GND_net), .CO(n3253));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(RX_ADDR[4]), .I2(GND_net), 
            .I3(n3248), .O(n122[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_6 (.CI(n3248), .I0(RX_ADDR[4]), .I1(GND_net), .CO(n3249));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(RX_ADDR[7]), .I2(GND_net), 
            .I3(n3251), .O(n122[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_9 (.CI(n3251), .I0(RX_ADDR[7]), .I1(GND_net), .CO(n3252));
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(RX_ADDR[6]), .I2(GND_net), 
            .I3(n3250), .O(n122[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_2 (.CI(VCC_net), .I0(RX_ADDR[0]), .I1(GND_net), .CO(n3245));
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(RX_ADDR[13]), .I2(GND_net), 
            .I3(n3257), .O(n122[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(RX_ADDR[12]), .I2(GND_net), 
            .I3(n3256), .O(n122[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_4 (.CI(n3246), .I0(RX_ADDR[2]), .I1(GND_net), .CO(n3247));
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(RX_ADDR[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n122[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n3256), .I0(RX_ADDR[12]), .I1(GND_net), .CO(n3257));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(RX_ADDR[1]), .I2(GND_net), 
            .I3(n3245), .O(n122[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(RX_ADDR[3]), .I2(GND_net), 
            .I3(n3247), .O(n122[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(RX_ADDR[11]), .I2(GND_net), 
            .I3(n3255), .O(n122[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR BRAM_ADDR__i2 (.Q(RX_ADDR[2]), .C(TVP_CLK_c), .D(n2723), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_DFFSR BRAM_ADDR__i1 (.Q(RX_ADDR[1]), .C(TVP_CLK_c), .D(n2721), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_DFFSR BRAM_ADDR__i0 (.Q(RX_ADDR[0]), .C(TVP_CLK_c), .D(n2719), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_DFFSR BRAM_ADDR__i10 (.Q(RX_ADDR[10]), .C(TVP_CLK_c), .D(n2717), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1469_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[3]), 
            .I3(RX_ADDR[3]), .O(n2703));
    defparam i1469_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i9 (.Q(RX_ADDR[9]), .C(TVP_CLK_c), .D(n2715), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1471_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[4]), 
            .I3(RX_ADDR[4]), .O(n2705));
    defparam i1471_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i8 (.Q(RX_ADDR[8]), .C(TVP_CLK_c), .D(n2713), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_DFFSR BRAM_ADDR__i7 (.Q(RX_ADDR[7]), .C(TVP_CLK_c), .D(n2711), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1473_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[5]), 
            .I3(RX_ADDR[5]), .O(n2707));
    defparam i1473_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i6 (.Q(RX_ADDR[6]), .C(TVP_CLK_c), .D(n2709), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1475_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[6]), 
            .I3(RX_ADDR[6]), .O(n2709));
    defparam i1475_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i5 (.Q(RX_ADDR[5]), .C(TVP_CLK_c), .D(n2707), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1477_3_lut_4_lut (.I0(RX_WE), .I1(TVP_VSYNC_c), .I2(n122[7]), 
            .I3(RX_ADDR[7]), .O(n2711));
    defparam i1477_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i4 (.Q(RX_ADDR[4]), .C(TVP_CLK_c), .D(n2705), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    SB_DFFSR BRAM_ADDR__i3 (.Q(RX_ADDR[3]), .C(TVP_CLK_c), .D(n2703), 
            .R(n3793));   // ../rx.v(51[12] 60[8])
    O_COUNTER rx_counter (.TVP_CLK_c(TVP_CLK_c), .GND_net(GND_net), .VCC_net(VCC_net), 
            .TVP_HSYNC_c(TVP_HSYNC_c), .TVP_VSYNC_c(TVP_VSYNC_c), .RX_WE(RX_WE), 
            .RX_TX_SYNC(RX_TX_SYNC), .LED_c(LED_c), .n3793(n3793)) /* synthesis syn_module_defined=1 */ ;   // ../rx.v(41[15] 49[41])
    
endmodule
//
// Verilog Description of module O_COUNTER
//

module O_COUNTER (TVP_CLK_c, GND_net, VCC_net, TVP_HSYNC_c, TVP_VSYNC_c, 
            RX_WE, RX_TX_SYNC, LED_c, n3793) /* synthesis syn_module_defined=1 */ ;
    input TVP_CLK_c;
    input GND_net;
    input VCC_net;
    input TVP_HSYNC_c;
    input TVP_VSYNC_c;
    output RX_WE;
    output RX_TX_SYNC;
    output LED_c;
    output n3793;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire [5:0]n29;
    
    wire n3792;
    wire [5:0]FRAME_COUNTER;   // ../o_counter.v(46[19:32])
    
    wire n2517, n3305;
    wire [9:0]X;   // ../o_counter.v(47[19:20])
    
    wire n3306;
    wire [9:0]n45;
    
    wire n3304, n6, n3534, n4, n3581;
    wire [8:0]n1;
    wire [8:0]Y;   // ../o_counter.v(48[19:20])
    
    wire old_HS, n5, n3548, n4_adj_604, n3575, n3278, n3307, n3308, 
        n3277, old_VS, O_VISIBLE_N_99, SYNC_N_114;
    wire [9:0]n79;
    
    wire n3790, n3551, n3791, n4_adj_606, n3271, n55_adj_607, n3302, 
        n3303, n3301, n3276, PULSE_1HZ_N_110, n7_adj_609, n3628, 
        n11, n2045, n10_adj_610, n14_adj_611, n3314, n3313, n3275, 
        n3274, n3273, n3272, n3312, n3311, n3310, n3309;
    
    SB_DFFESR FRAME_COUNTER_243__i0 (.Q(FRAME_COUNTER[0]), .C(TVP_CLK_c), 
            .E(n3792), .D(n29[0]), .R(n2517));   // ../o_counter.v(72[46:66])
    SB_CARRY X_242_add_4_7 (.CI(n3305), .I0(GND_net), .I1(X[5]), .CO(n3306));
    SB_LUT4 X_242_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(X[4]), 
            .I3(n3304), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2208_4_lut (.I0(X[3]), .I1(X[7]), .I2(n6), .I3(X[6]), .O(n3534));
    defparam i2208_4_lut.LUT_INIT = 16'hccc8;
    SB_DFFESR FRAME_COUNTER_243__i3 (.Q(FRAME_COUNTER[3]), .C(TVP_CLK_c), 
            .E(n3792), .D(n29[3]), .R(n2517));   // ../o_counter.v(72[46:66])
    SB_LUT4 i2_4_lut (.I0(X[7]), .I1(X[6]), .I2(X[5]), .I3(n4), .O(n3581));
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 add_5_2_lut (.I0(GND_net), .I1(Y[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF old_HS_51 (.Q(old_HS), .C(TVP_CLK_c), .D(TVP_HSYNC_c));   // ../o_counter.v(51[16] 84[12])
    SB_LUT4 i3_4_lut (.I0(n5), .I1(Y[8]), .I2(n3548), .I3(n4_adj_604), 
            .O(n3575));
    defparam i3_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 add_5_10_lut (.I0(GND_net), .I1(Y[8]), .I2(GND_net), .I3(n3278), 
            .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_242_add_4_9 (.CI(n3307), .I0(GND_net), .I1(X[7]), .CO(n3308));
    SB_LUT4 add_5_9_lut (.I0(GND_net), .I1(Y[7]), .I2(GND_net), .I3(n3277), 
            .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF old_VS_52 (.Q(old_VS), .C(TVP_CLK_c), .D(TVP_VSYNC_c));   // ../o_counter.v(51[16] 84[12])
    SB_CARRY X_242_add_4_6 (.CI(n3304), .I0(GND_net), .I1(X[4]), .CO(n3305));
    SB_DFF O_VISIBLE_53 (.Q(RX_WE), .C(TVP_CLK_c), .D(O_VISIBLE_N_99));   // ../o_counter.v(51[16] 84[12])
    SB_DFF SYNC_46 (.Q(RX_TX_SYNC), .C(TVP_CLK_c), .D(SYNC_N_114));   // ../o_counter.v(51[16] 84[12])
    SB_DFFSR X_242__i0 (.Q(n79[0]), .C(TVP_CLK_c), .D(n45[0]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_LUT4 i1_4_lut (.I0(n3551), .I1(Y[7]), .I2(n3791), .I3(Y[4]), 
            .O(n4_adj_606));
    defparam i1_4_lut.LUT_INIT = 16'hc8c0;
    SB_CARRY add_5_2 (.CI(VCC_net), .I0(Y[0]), .I1(GND_net), .CO(n3271));
    SB_LUT4 i59_4_lut (.I0(X[8]), .I1(n3581), .I2(X[9]), .I3(n3534), 
            .O(n55_adj_607));
    defparam i59_4_lut.LUT_INIT = 16'he0e5;
    SB_LUT4 i2363_4_lut (.I0(Y[8]), .I1(n55_adj_607), .I2(n4_adj_606), 
            .I3(n3575), .O(O_VISIBLE_N_99));
    defparam i2363_4_lut.LUT_INIT = 16'h1300;
    SB_CARRY X_242_add_4_4 (.CI(n3302), .I0(GND_net), .I1(n79[2]), .CO(n3303));
    SB_CARRY add_5_9 (.CI(n3277), .I0(Y[7]), .I1(GND_net), .CO(n3278));
    SB_LUT4 X_242_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(X[3]), 
            .I3(n3303), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 X_242_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(n79[1]), 
            .I3(n3301), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5_8_lut (.I0(GND_net), .I1(Y[6]), .I2(GND_net), .I3(n3276), 
            .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_242_add_4_3 (.CI(n3301), .I0(GND_net), .I1(n79[1]), .CO(n3302));
    SB_DFFE PULSE_1HZ_49 (.Q(LED_c), .C(TVP_CLK_c), .E(n3792), .D(PULSE_1HZ_N_110));   // ../o_counter.v(51[16] 84[12])
    SB_CARRY add_5_8 (.CI(n3276), .I0(Y[6]), .I1(GND_net), .CO(n3277));
    SB_LUT4 X_242_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n79[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_242_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n79[0]), .CO(n3301));
    SB_LUT4 i1_2_lut (.I0(FRAME_COUNTER[2]), .I1(FRAME_COUNTER[4]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_609));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2302_2_lut (.I0(FRAME_COUNTER[1]), .I1(FRAME_COUNTER[5]), .I2(GND_net), 
            .I3(GND_net), .O(n3628));
    defparam i2302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n3628), .I1(n7_adj_609), .I2(FRAME_COUNTER[3]), 
            .I3(FRAME_COUNTER[0]), .O(n11));
    defparam i5_4_lut.LUT_INIT = 16'hdfff;
    SB_LUT4 i1_2_lut_adj_18 (.I0(LED_c), .I1(n11), .I2(GND_net), .I3(GND_net), 
            .O(PULSE_1HZ_N_110));
    defparam i1_2_lut_adj_18.LUT_INIT = 16'h9999;
    SB_LUT4 i248_3_lut_3_lut_3_lut (.I0(TVP_VSYNC_c), .I1(old_HS), .I2(TVP_HSYNC_c), 
            .I3(GND_net), .O(n2045));   // ../o_counter.v(65[19:33])
    defparam i248_3_lut_3_lut_3_lut.LUT_INIT = 16'h5d5d;
    SB_LUT4 O_VS_I_0_1_lut_rep_26 (.I0(TVP_VSYNC_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3793));   // ../o_counter.v(65[19:33])
    defparam O_VS_I_0_1_lut_rep_26.LUT_INIT = 16'h5555;
    SB_LUT4 i1286_2_lut_3_lut (.I0(old_VS), .I1(TVP_VSYNC_c), .I2(n11), 
            .I3(GND_net), .O(n2517));   // ../o_counter.v(65[16] 75[19])
    defparam i1286_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i129_2_lut_rep_25 (.I0(old_VS), .I1(TVP_VSYNC_c), .I2(GND_net), 
            .I3(GND_net), .O(n3792));   // ../o_counter.v(65[16] 75[19])
    defparam i129_2_lut_rep_25.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut (.I0(Y[7]), .I1(Y[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_610));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(Y[8]), .I1(Y[2]), .I2(Y[1]), .I3(Y[3]), .O(n14_adj_611));
    defparam i6_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 FRAME_COUNTER_243_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[5]), 
            .I3(n3314), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_243_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 FRAME_COUNTER_243_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[4]), 
            .I3(n3313), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_243_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5_7_lut (.I0(GND_net), .I1(Y[5]), .I2(GND_net), .I3(n3275), 
            .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_242_add_4_5 (.CI(n3303), .I0(GND_net), .I1(X[3]), .CO(n3304));
    SB_CARRY add_5_7 (.CI(n3275), .I0(Y[5]), .I1(GND_net), .CO(n3276));
    SB_LUT4 add_5_6_lut (.I0(GND_net), .I1(Y[4]), .I2(GND_net), .I3(n3274), 
            .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5_6 (.CI(n3274), .I0(Y[4]), .I1(GND_net), .CO(n3275));
    SB_LUT4 add_5_5_lut (.I0(GND_net), .I1(Y[3]), .I2(GND_net), .I3(n3273), 
            .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5_5 (.CI(n3273), .I0(Y[3]), .I1(GND_net), .CO(n3274));
    SB_LUT4 X_242_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(X[6]), 
            .I3(n3306), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5_4_lut (.I0(GND_net), .I1(Y[2]), .I2(GND_net), .I3(n3272), 
            .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5_4 (.CI(n3272), .I0(Y[2]), .I1(GND_net), .CO(n3273));
    SB_LUT4 add_5_3_lut (.I0(GND_net), .I1(Y[1]), .I2(GND_net), .I3(n3271), 
            .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_242_add_4_8 (.CI(n3306), .I0(GND_net), .I1(X[6]), .CO(n3307));
    SB_LUT4 X_242_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(n79[2]), 
            .I3(n3302), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 X_242_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(X[5]), 
            .I3(n3305), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_243_add_4_6 (.CI(n3313), .I0(GND_net), .I1(FRAME_COUNTER[4]), 
            .CO(n3314));
    SB_LUT4 FRAME_COUNTER_243_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[3]), 
            .I3(n3312), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_243_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR X_242__i1 (.Q(n79[1]), .C(TVP_CLK_c), .D(n45[1]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_DFFSR X_242__i2 (.Q(n79[2]), .C(TVP_CLK_c), .D(n45[2]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_CARRY FRAME_COUNTER_243_add_4_5 (.CI(n3312), .I0(GND_net), .I1(FRAME_COUNTER[3]), 
            .CO(n3313));
    SB_LUT4 FRAME_COUNTER_243_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[2]), 
            .I3(n3311), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_243_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_243_add_4_4 (.CI(n3311), .I0(GND_net), .I1(FRAME_COUNTER[2]), 
            .CO(n3312));
    SB_CARRY add_5_3 (.CI(n3271), .I0(Y[1]), .I1(GND_net), .CO(n3272));
    SB_DFFSR X_242__i3 (.Q(X[3]), .C(TVP_CLK_c), .D(n45[3]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_DFFSR X_242__i4 (.Q(X[4]), .C(TVP_CLK_c), .D(n45[4]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_DFFSR X_242__i5 (.Q(X[5]), .C(TVP_CLK_c), .D(n45[5]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_DFFSR X_242__i6 (.Q(X[6]), .C(TVP_CLK_c), .D(n45[6]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_DFFSR X_242__i7 (.Q(X[7]), .C(TVP_CLK_c), .D(n45[7]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_DFFSR X_242__i8 (.Q(X[8]), .C(TVP_CLK_c), .D(n45[8]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_DFFSR X_242__i9 (.Q(X[9]), .C(TVP_CLK_c), .D(n45[9]), .R(n3790));   // ../o_counter.v(62[26:35])
    SB_LUT4 i2360_4_lut (.I0(Y[0]), .I1(n14_adj_611), .I2(n10_adj_610), 
            .I3(n3791), .O(SYNC_N_114));   // ../o_counter.v(53[21:33])
    defparam i2360_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut (.I0(Y[5]), .I1(Y[6]), .I2(Y[7]), .I3(GND_net), 
            .O(n5));   // ../o_counter.v(81[116:145])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i592_2_lut_rep_24 (.I0(Y[5]), .I1(Y[6]), .I2(GND_net), .I3(GND_net), 
            .O(n3791));   // ../o_counter.v(81[116:145])
    defparam i592_2_lut_rep_24.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_19 (.I0(X[5]), .I1(X[4]), .I2(GND_net), .I3(GND_net), 
            .O(n6));
    defparam i2_2_lut_adj_19.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_20 (.I0(Y[4]), .I1(Y[3]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_604));
    defparam i1_2_lut_adj_20.LUT_INIT = 16'h8888;
    SB_LUT4 i5_1_lut_rep_23 (.I0(TVP_HSYNC_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3790));   // ../o_counter.v(56[19:33])
    defparam i5_1_lut_rep_23.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(Y[1]), .I1(Y[0]), .I2(Y[2]), .I3(GND_net), 
            .O(n3548));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 FRAME_COUNTER_243_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[1]), 
            .I3(n3310), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_243_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_243_add_4_3 (.CI(n3310), .I0(GND_net), .I1(FRAME_COUNTER[1]), 
            .CO(n3311));
    SB_LUT4 FRAME_COUNTER_243_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[0]), 
            .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_243_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_243_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(FRAME_COUNTER[0]), 
            .CO(n3310));
    SB_LUT4 X_242_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(X[9]), 
            .I3(n3309), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR Y__i0 (.Q(Y[0]), .C(TVP_CLK_c), .E(n2045), .D(n1[0]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_DFFESR Y__i8 (.Q(Y[8]), .C(TVP_CLK_c), .E(n2045), .D(n1[8]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_LUT4 i2_4_lut_adj_21 (.I0(Y[2]), .I1(Y[3]), .I2(Y[0]), .I3(Y[1]), 
            .O(n3551));
    defparam i2_4_lut_adj_21.LUT_INIT = 16'hfeee;
    SB_LUT4 X_242_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(X[8]), 
            .I3(n3308), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_242_add_4_10 (.CI(n3308), .I0(GND_net), .I1(X[8]), .CO(n3309));
    SB_LUT4 i1_2_lut_adj_22 (.I0(X[4]), .I1(X[3]), .I2(GND_net), .I3(GND_net), 
            .O(n4));
    defparam i1_2_lut_adj_22.LUT_INIT = 16'heeee;
    SB_DFFESR Y__i7 (.Q(Y[7]), .C(TVP_CLK_c), .E(n2045), .D(n1[7]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_DFFESR Y__i6 (.Q(Y[6]), .C(TVP_CLK_c), .E(n2045), .D(n1[6]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_DFFESR Y__i5 (.Q(Y[5]), .C(TVP_CLK_c), .E(n2045), .D(n1[5]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_DFFESR Y__i4 (.Q(Y[4]), .C(TVP_CLK_c), .E(n2045), .D(n1[4]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_DFFESR Y__i3 (.Q(Y[3]), .C(TVP_CLK_c), .E(n2045), .D(n1[3]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_DFFESR Y__i2 (.Q(Y[2]), .C(TVP_CLK_c), .E(n2045), .D(n1[2]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_DFFESR Y__i1 (.Q(Y[1]), .C(TVP_CLK_c), .E(n2045), .D(n1[1]), 
            .R(n3793));   // ../o_counter.v(51[16] 84[12])
    SB_DFFESR FRAME_COUNTER_243__i5 (.Q(FRAME_COUNTER[5]), .C(TVP_CLK_c), 
            .E(n3792), .D(n29[5]), .R(n2517));   // ../o_counter.v(72[46:66])
    SB_DFFESR FRAME_COUNTER_243__i1 (.Q(FRAME_COUNTER[1]), .C(TVP_CLK_c), 
            .E(n3792), .D(n29[1]), .R(n2517));   // ../o_counter.v(72[46:66])
    SB_DFFESR FRAME_COUNTER_243__i4 (.Q(FRAME_COUNTER[4]), .C(TVP_CLK_c), 
            .E(n3792), .D(n29[4]), .R(n2517));   // ../o_counter.v(72[46:66])
    SB_LUT4 X_242_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(X[7]), 
            .I3(n3307), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam X_242_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR FRAME_COUNTER_243__i2 (.Q(FRAME_COUNTER[2]), .C(TVP_CLK_c), 
            .E(n3792), .D(n29[2]), .R(n2517));   // ../o_counter.v(72[46:66])
    
endmodule
//
// Verilog Description of module RAM
//

module RAM (TX_DATA, ADV_CLK_c, \TX_ADDR[12] , \TX_ADDR[13] , \TX_ADDR[11] , 
            GND_net, RX_ADDR, n28, n27, n26, n25, n24, n23, 
            n22, n21, n20, n19, n18, TVP_VIDEO_c_8, TVP_VIDEO_c_9, 
            TVP_CLK_c, VCC_net, TVP_VIDEO_c_6, TVP_VIDEO_c_7, TVP_VIDEO_c_4, 
            TVP_VIDEO_c_5, TVP_VIDEO_c_2, TVP_VIDEO_c_3, RX_WE) /* synthesis syn_module_defined=1 */ ;
    output [7:0]TX_DATA;
    input ADV_CLK_c;
    input \TX_ADDR[12] ;
    input \TX_ADDR[13] ;
    input \TX_ADDR[11] ;
    input GND_net;
    input [13:0]RX_ADDR;
    input n28;
    input n27;
    input n26;
    input n25;
    input n24;
    input n23;
    input n22;
    input n21;
    input n20;
    input n19;
    input n18;
    input TVP_VIDEO_c_8;
    input TVP_VIDEO_c_9;
    input TVP_CLK_c;
    input VCC_net;
    input TVP_VIDEO_c_6;
    input TVP_VIDEO_c_7;
    input TVP_VIDEO_c_4;
    input TVP_VIDEO_c_5;
    input TVP_VIDEO_c_2;
    input TVP_VIDEO_c_3;
    input RX_WE;
    
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire [7:0]dout_7__N_596;
    
    wire n3676, n3677, n3716, n3674, n3673, n534, n542, n3710, 
        n445, n437, n3713, n565, n573, n538, n546, n3704, n449, 
        n441, n3707, n501, n509, n3749, n3755, n505, n506, n516, 
        n438, n439, n451, n436, n434, n435, n503, n504, n537, 
        n548, n502, n499, n500, n535, n536, n448, n452, n533, 
        n531, n532, n446, n447, n569, n570, n580, n444, n442, 
        n443, n567, n568, n513, n514, n517, n566, n563, n564, 
        n511, n512, n545, n549, n510, n507, n508, n544, n3698, 
        n543, n577, n578, n581, n541, n539, n540, n575, n576, 
        n440, n574, n571, n572, n3701, n3646, n3647, n3722, 
        n3679, n3680, n3640, n3641, n3635, n3634, n3764, n3767, 
        n3758, n3761, n3752, n3746, n3737, n3692, n3740, n3743, 
        n3695, n3734, n3728;
    
    SB_DFF dout_i0 (.Q(TX_DATA[0]), .C(ADV_CLK_c), .D(dout_7__N_596[0]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 TX_ADDR_12__bdd_4_lut_2392 (.I0(\TX_ADDR[12] ), .I1(n3676), 
            .I2(n3677), .I3(\TX_ADDR[13] ), .O(n3716));
    defparam TX_ADDR_12__bdd_4_lut_2392.LUT_INIT = 16'he4aa;
    SB_LUT4 n3716_bdd_4_lut (.I0(n3716), .I1(n3674), .I2(n3673), .I3(\TX_ADDR[13] ), 
            .O(dout_7__N_596[2]));
    defparam n3716_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2402 (.I0(\TX_ADDR[11] ), .I1(n534), .I2(n542), 
            .I3(\TX_ADDR[12] ), .O(n3710));
    defparam TX_ADDR_11__bdd_4_lut_2402.LUT_INIT = 16'he4aa;
    SB_LUT4 n3710_bdd_4_lut (.I0(n3710), .I1(n445), .I2(n437), .I3(\TX_ADDR[12] ), 
            .O(n3713));
    defparam n3710_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2351_3_lut (.I0(n565), .I1(n573), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3677));
    defparam i2351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2383 (.I0(\TX_ADDR[11] ), .I1(n538), .I2(n546), 
            .I3(\TX_ADDR[12] ), .O(n3704));
    defparam TX_ADDR_11__bdd_4_lut_2383.LUT_INIT = 16'he4aa;
    SB_LUT4 n3704_bdd_4_lut (.I0(n3704), .I1(n449), .I2(n441), .I3(\TX_ADDR[12] ), 
            .O(n3707));
    defparam n3704_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2350_3_lut (.I0(n501), .I1(n509), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3676));
    defparam i2350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i172111_i1_3_lut (.I0(n3749), .I1(n3755), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_596[0]));
    defparam i172111_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_RAM2048x2 mem0 (.RDATA({n506, n505}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n516), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem0.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem0.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem0.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem0.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem0.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem0.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem0.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem0.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem0.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem8 (.RDATA({n439, n438}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n451), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem8.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem8.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem8.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem8.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem8.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem8.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem8.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem8.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem9 (.RDATA({n437, n436}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n451), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem9.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem9.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem9.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem9.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem9.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem9.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem9.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem9.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem10 (.RDATA({n435, n434}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n451), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem10.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem10.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem10.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem10.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem10.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem10.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem10.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem10.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem11 (.RDATA({n504, n503}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n516), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem11.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem11.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem11.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem11.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem11.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem11.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem11.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem11.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem11.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem1 (.RDATA({n538, n537}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n548), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem1.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem1.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem1.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem1.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem1.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem1.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem1.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem1.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem1.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem1.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem12 (.RDATA({n502, n501}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n516), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem12.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem12.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem12.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem12.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem12.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem12.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem12.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem13 (.RDATA({n500, n499}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n516), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem13.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem13.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem13.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem13.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem13.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem13.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem13.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem13.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem13.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem14 (.RDATA({n536, n535}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n548), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem14.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem14.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem14.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem14.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem14.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem14.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem14.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem14.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem14.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem14.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem2 (.RDATA({n449, n448}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n452), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem2.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem2.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem2.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem2.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem2.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem2.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem2.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem2.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    SB_RAM2048x2 mem15 (.RDATA({n534, n533}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n548), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem15.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem15.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem15.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem15.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem15.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem15.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem15.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem15.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem15.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem15.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem16 (.RDATA({n532, n531}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n548), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem16.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem16.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem16.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem16.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem16.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem16.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem16.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem16.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem16.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem16.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem17 (.RDATA({n447, n446}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n452), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem17.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem17.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem17.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem17.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem17.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem17.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem17.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem17.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    SB_RAM2048x2 mem3 (.RDATA({n570, n569}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n580), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem3.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem3.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem3.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem3.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem3.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem3.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem3.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem3.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem3.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem18 (.RDATA({n445, n444}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n452), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem18.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem18.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem18.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem18.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem18.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem18.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem18.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem18.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    SB_RAM2048x2 mem19 (.RDATA({n443, n442}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n452), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem19.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem19.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem19.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem19.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem19.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem19.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem19.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem19.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    SB_RAM2048x2 mem20 (.RDATA({n568, n567}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n580), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem20.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem20.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem20.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem20.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem20.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem20.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem20.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem20.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem20.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem4 (.RDATA({n514, n513}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n517), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem4.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem4.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem4.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem4.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem4.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem4.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem4.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem4.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem21 (.RDATA({n566, n565}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n580), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem21.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem21.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem21.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem21.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem21.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem21.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem21.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem21.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem21.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem22 (.RDATA({n564, n563}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n580), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem22.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem22.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem22.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem22.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem22.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem22.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem22.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem22.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem22.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem23 (.RDATA({n512, n511}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n517), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem23.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem23.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem23.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem23.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem23.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem23.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem23.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem23.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem5 (.RDATA({n546, n545}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n549), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem5.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem5.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem5.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem5.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem5.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem5.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem5.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem5.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem5.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem5.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem5.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem24 (.RDATA({n510, n509}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n517), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem24.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem24.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem24.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem24.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem24.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem24.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem24.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem24.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem25 (.RDATA({n508, n507}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n517), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem25.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem25.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem25.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem25.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem25.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem25.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem25.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem25.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2378 (.I0(\TX_ADDR[11] ), .I1(n536), .I2(n544), 
            .I3(\TX_ADDR[12] ), .O(n3698));
    defparam TX_ADDR_11__bdd_4_lut_2378.LUT_INIT = 16'he4aa;
    SB_RAM2048x2 mem26 (.RDATA({n544, n543}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n549), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem26.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem26.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem26.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem26.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem26.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem26.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem26.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem26.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem26.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem26.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem26.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem6 (.RDATA({n578, n577}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n581), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem6.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem6.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem6.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem6.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem6.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem6.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem6.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem6.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem6.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem6.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem6.INIT_E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    defparam mem6.INIT_F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    SB_RAM2048x2 mem27 (.RDATA({n542, n541}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n549), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem27.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem27.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem27.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem27.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem27.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem27.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem27.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem27.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem27.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem27.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem27.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem28 (.RDATA({n540, n539}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n549), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem28.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem28.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem28.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem28.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem28.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem28.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem28.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem28.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem28.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem28.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem28.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem29 (.RDATA({n576, n575}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n581), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_7, 
            TVP_VIDEO_c_6}));
    defparam mem29.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem29.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem29.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem29.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem29.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem29.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem29.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem29.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem29.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem29.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem29.INIT_E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    defparam mem29.INIT_F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    SB_RAM2048x2 mem7 (.RDATA({n441, n440}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n451), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_9, 
            TVP_VIDEO_c_8}));
    defparam mem7.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem7.INIT_5 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem7.INIT_6 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem7.INIT_7 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem7.INIT_8 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem7.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem7.INIT_E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem7.INIT_F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    SB_RAM2048x2 mem30 (.RDATA({n574, n573}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n581), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_5, 
            TVP_VIDEO_c_4}));
    defparam mem30.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem30.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem30.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem30.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem30.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem30.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem30.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem30.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem30.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem30.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem30.INIT_E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    defparam mem30.INIT_F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    SB_RAM2048x2 mem31 (.RDATA({n572, n571}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n581), .WADDR({RX_ADDR[10:0]}), .WDATA({TVP_VIDEO_c_3, 
            TVP_VIDEO_c_2}));
    defparam mem31.INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem31.INIT_1 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem31.INIT_2 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem31.INIT_3 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem31.INIT_4 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem31.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_9 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000;
    defparam mem31.INIT_A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem31.INIT_B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem31.INIT_C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem31.INIT_D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam mem31.INIT_E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    defparam mem31.INIT_F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    SB_LUT4 n3698_bdd_4_lut (.I0(n3698), .I1(n447), .I2(n439), .I3(\TX_ADDR[12] ), 
            .O(n3701));
    defparam n3698_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_12__bdd_4_lut_2397 (.I0(\TX_ADDR[12] ), .I1(n3646), 
            .I2(n3647), .I3(\TX_ADDR[13] ), .O(n3722));
    defparam TX_ADDR_12__bdd_4_lut_2397.LUT_INIT = 16'he4aa;
    SB_LUT4 i2347_3_lut (.I0(n436), .I1(n444), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3673));
    defparam i2347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2353_3_lut (.I0(n440), .I1(n448), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3679));
    defparam i2353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2354_3_lut (.I0(n537), .I1(n545), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3680));
    defparam i2354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2314_3_lut (.I0(n438), .I1(n446), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3640));
    defparam i2314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2315_3_lut (.I0(n535), .I1(n543), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3641));
    defparam i2315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2309_3_lut (.I0(n567), .I1(n575), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3635));
    defparam i2309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2308_3_lut (.I0(n503), .I1(n511), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3634));
    defparam i2308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2348_3_lut (.I0(n533), .I1(n541), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3674));
    defparam i2348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut (.I0(\TX_ADDR[11] ), .I1(n570), .I2(n578), 
            .I3(\TX_ADDR[12] ), .O(n3764));
    defparam TX_ADDR_11__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n3764_bdd_4_lut (.I0(n3764), .I1(n514), .I2(n506), .I3(\TX_ADDR[12] ), 
            .O(n3767));
    defparam n3764_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2427 (.I0(\TX_ADDR[11] ), .I1(n566), .I2(n574), 
            .I3(\TX_ADDR[12] ), .O(n3758));
    defparam TX_ADDR_11__bdd_4_lut_2427.LUT_INIT = 16'he4aa;
    SB_LUT4 n3758_bdd_4_lut (.I0(n3758), .I1(n510), .I2(n502), .I3(\TX_ADDR[12] ), 
            .O(n3761));
    defparam n3758_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i176332_i1_3_lut (.I0(n3707), .I1(n3767), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_596[7]));
    defparam i176332_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dout_i1 (.Q(TX_DATA[1]), .C(ADV_CLK_c), .D(dout_7__N_596[1]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i2 (.Q(TX_DATA[2]), .C(ADV_CLK_c), .D(dout_7__N_596[2]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i3 (.Q(TX_DATA[3]), .C(ADV_CLK_c), .D(dout_7__N_596[3]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i4 (.Q(TX_DATA[4]), .C(ADV_CLK_c), .D(dout_7__N_596[4]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i5 (.Q(TX_DATA[5]), .C(ADV_CLK_c), .D(dout_7__N_596[5]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i6 (.Q(TX_DATA[6]), .C(ADV_CLK_c), .D(dout_7__N_596[6]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i7 (.Q(TX_DATA[7]), .C(ADV_CLK_c), .D(dout_7__N_596[7]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2422 (.I0(\TX_ADDR[11] ), .I1(n563), .I2(n571), 
            .I3(\TX_ADDR[12] ), .O(n3752));
    defparam TX_ADDR_11__bdd_4_lut_2422.LUT_INIT = 16'he4aa;
    SB_LUT4 n3752_bdd_4_lut (.I0(n3752), .I1(n507), .I2(n499), .I3(\TX_ADDR[12] ), 
            .O(n3755));
    defparam n3752_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2417 (.I0(\TX_ADDR[11] ), .I1(n531), .I2(n539), 
            .I3(\TX_ADDR[12] ), .O(n3746));
    defparam TX_ADDR_11__bdd_4_lut_2417.LUT_INIT = 16'he4aa;
    SB_LUT4 n3746_bdd_4_lut (.I0(n3746), .I1(n442), .I2(n434), .I3(\TX_ADDR[12] ), 
            .O(n3749));
    defparam n3746_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i175126_i1_3_lut (.I0(n3701), .I1(n3737), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_596[5]));
    defparam i175126_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i173920_i1_3_lut (.I0(n3713), .I1(n3761), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_596[3]));
    defparam i173920_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2373 (.I0(\TX_ADDR[11] ), .I1(n564), .I2(n572), 
            .I3(\TX_ADDR[12] ), .O(n3692));
    defparam TX_ADDR_11__bdd_4_lut_2373.LUT_INIT = 16'he4aa;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2412 (.I0(\TX_ADDR[11] ), .I1(n532), .I2(n540), 
            .I3(\TX_ADDR[12] ), .O(n3740));
    defparam TX_ADDR_11__bdd_4_lut_2412.LUT_INIT = 16'he4aa;
    SB_LUT4 n3740_bdd_4_lut (.I0(n3740), .I1(n443), .I2(n435), .I3(\TX_ADDR[12] ), 
            .O(n3743));
    defparam n3740_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i172714_i1_3_lut (.I0(n3743), .I1(n3695), .I2(\TX_ADDR[13] ), 
            .I3(GND_net), .O(dout_7__N_596[1]));
    defparam i172714_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2407 (.I0(\TX_ADDR[11] ), .I1(n568), .I2(n576), 
            .I3(\TX_ADDR[12] ), .O(n3734));
    defparam TX_ADDR_11__bdd_4_lut_2407.LUT_INIT = 16'he4aa;
    SB_LUT4 i2321_3_lut (.I0(n569), .I1(n577), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3647));
    defparam i2321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2320_3_lut (.I0(n505), .I1(n513), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3646));
    defparam i2320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n3734_bdd_4_lut (.I0(n3734), .I1(n512), .I2(n504), .I3(\TX_ADDR[12] ), 
            .O(n3737));
    defparam n3734_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_12__bdd_4_lut (.I0(\TX_ADDR[12] ), .I1(n3634), .I2(n3635), 
            .I3(\TX_ADDR[13] ), .O(n3728));
    defparam TX_ADDR_12__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n3692_bdd_4_lut (.I0(n3692), .I1(n508), .I2(n500), .I3(\TX_ADDR[12] ), 
            .O(n3695));
    defparam n3692_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n3728_bdd_4_lut (.I0(n3728), .I1(n3641), .I2(n3640), .I3(\TX_ADDR[13] ), 
            .O(dout_7__N_596[4]));
    defparam n3728_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n3722_bdd_4_lut (.I0(n3722), .I1(n3680), .I2(n3679), .I3(\TX_ADDR[13] ), 
            .O(dout_7__N_596[6]));
    defparam n3722_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(RX_WE), .I1(RX_ADDR[13]), .I2(RX_ADDR[12]), 
            .I3(RX_ADDR[11]), .O(n580));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_11 (.I0(RX_WE), .I1(RX_ADDR[13]), .I2(RX_ADDR[12]), 
            .I3(RX_ADDR[11]), .O(n581));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_11.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_12 (.I0(RX_WE), .I1(RX_ADDR[13]), .I2(RX_ADDR[12]), 
            .I3(RX_ADDR[11]), .O(n517));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_12.LUT_INIT = 16'h0800;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.I0(RX_WE), .I1(RX_ADDR[13]), .I2(RX_ADDR[12]), 
            .I3(RX_ADDR[11]), .O(n516));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_13.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_14 (.I0(RX_WE), .I1(RX_ADDR[13]), .I2(RX_ADDR[11]), 
            .I3(RX_ADDR[12]), .O(n451));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_14.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_15 (.I0(RX_WE), .I1(RX_ADDR[13]), .I2(RX_ADDR[11]), 
            .I3(RX_ADDR[12]), .O(n548));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_15.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_16 (.I0(RX_WE), .I1(RX_ADDR[13]), .I2(RX_ADDR[11]), 
            .I3(RX_ADDR[12]), .O(n549));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_16.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_17 (.I0(RX_WE), .I1(RX_ADDR[13]), .I2(RX_ADDR[11]), 
            .I3(RX_ADDR[12]), .O(n452));   // ../ram.v(12[4:14])
    defparam i1_2_lut_3_lut_4_lut_adj_17.LUT_INIT = 16'h0020;
    
endmodule
//
// Verilog Description of module TX_PLL
//

module TX_PLL (TVP_CLK_c, VCC_net, GND_net, ADV_CLK_c) /* synthesis syn_module_defined=1 */ ;
    input TVP_CLK_c;
    input VCC_net;
    input GND_net;
    output ADV_CLK_c;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    
    SB_PLL40_CORE TX_PLL_inst (.REFERENCECLK(TVP_CLK_c), .PLLOUTCORE(ADV_CLK_c), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=17, LSE_LCOL=9, LSE_RCOL=27, LSE_LLINE=20, LSE_RLINE=24 */ ;   // ../main.v(20[9] 24[27])
    defparam TX_PLL_inst.FEEDBACK_PATH = "SIMPLE";
    defparam TX_PLL_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam TX_PLL_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam TX_PLL_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam TX_PLL_inst.FDA_FEEDBACK = 4'b0000;
    defparam TX_PLL_inst.FDA_RELATIVE = 4'b0000;
    defparam TX_PLL_inst.PLLOUT_SELECT = "GENCLK";
    defparam TX_PLL_inst.DIVR = 4'b0000;
    defparam TX_PLL_inst.DIVF = 7'b0100110;
    defparam TX_PLL_inst.DIVQ = 3'b100;
    defparam TX_PLL_inst.FILTER_RANGE = 3'b010;
    defparam TX_PLL_inst.ENABLE_ICEGATE = 1'b0;
    defparam TX_PLL_inst.TEST_MODE = 1'b0;
    defparam TX_PLL_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
