-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 30 2018 19:21:12

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    TVP_VIDEO : in std_logic_vector(9 downto 0);
    ADV_B : out std_logic_vector(7 downto 0);
    ADV_G : out std_logic_vector(7 downto 0);
    ADV_R : out std_logic_vector(7 downto 0);
    DEBUG : inout std_logic_vector(7 downto 0);
    TVP_CLK : in std_logic;
    ADV_CLK : out std_logic;
    TVP_HSYNC : in std_logic;
    ADV_HSYNC : out std_logic;
    TVP_VSYNC : in std_logic;
    ADV_VSYNC : out std_logic;
    ADV_BLANK_N : out std_logic;
    LED : out std_logic;
    ADV_SYNC_N : out std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \GB_BUFFER_DEBUG_c_2_c_THRU_CO\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_70\ : std_logic;
signal \TVP_VIDEO_c_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_71\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_35\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_34\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_72\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_90\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_89\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_88\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_36\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_81\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_80\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_37\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_79\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_66\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_69\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_68\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_67\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_48\ : std_logic;
signal \TVP_VIDEO_c_2\ : std_logic;
signal \line_buffer.n533\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_82\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_49\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_84\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_83\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_85\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_87\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_86\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_91\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_93\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_92\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_94\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_97\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_98\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_96\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_95\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_33\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_29\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_32\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_31\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_30\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_74\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_73\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_65\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_64\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_63\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_75\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_62\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_78\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_2\ : std_logic;
signal \LED_c\ : std_logic;
signal \DEBUG_c_1_c\ : std_logic;
signal \tvp_hs_buffer.BUFFER_0_0\ : std_logic;
signal \tvp_hs_buffer.BUFFER_1_0\ : std_logic;
signal \receive_module.rx_counter.n10\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \receive_module.rx_counter.n9_adj_612\ : std_logic;
signal \receive_module.rx_counter.n3147\ : std_logic;
signal \receive_module.rx_counter.n8_adj_611\ : std_logic;
signal \receive_module.rx_counter.n3148\ : std_logic;
signal \receive_module.rx_counter.n3149\ : std_logic;
signal \receive_module.rx_counter.n3150\ : std_logic;
signal \receive_module.rx_counter.n3151\ : std_logic;
signal \receive_module.rx_counter.n3152\ : std_logic;
signal \receive_module.rx_counter.n3153\ : std_logic;
signal \receive_module.rx_counter.n3154\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \receive_module.rx_counter.n3155\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_50\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_51\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_58\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_57\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_22\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_21\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_24\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_23\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_28\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_27\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_26\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_25\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_99\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_38\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_40\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_39\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_41\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_42\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_43\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_59\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_45\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_44\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_47\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_46\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_61\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_60\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_77\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_76\ : std_logic;
signal n24 : std_logic;
signal \TVP_VIDEO_c_4\ : std_logic;
signal \DEBUG_c_0_c\ : std_logic;
signal \INVTVP_VSYNC_buff_I_0.BUFFER_0__i1C_net\ : std_logic;
signal \TVP_VSYNC_buff_I_0.BUFFER_0_0\ : std_logic;
signal \INVTVP_VSYNC_buff_I_0.BUFFER_0__i2C_net\ : std_logic;
signal \receive_module.rx_counter.X_8\ : std_logic;
signal \receive_module.rx_counter.X_9\ : std_logic;
signal \receive_module.rx_counter.n3630\ : std_logic;
signal \TVP_VSYNC_buff_I_0.BUFFER_1_0\ : std_logic;
signal \INVTVP_VSYNC_buff_I_0.WIRE_OUT_0__9C_net\ : std_logic;
signal \line_buffer.n467\ : std_logic;
signal \receive_module.rx_counter.n4_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3400\ : std_logic;
signal \line_buffer.n565\ : std_logic;
signal \receive_module.rx_counter.X_5\ : std_logic;
signal \receive_module.rx_counter.X_4\ : std_logic;
signal \receive_module.rx_counter.X_3\ : std_logic;
signal \receive_module.rx_counter.X_6\ : std_logic;
signal \receive_module.rx_counter.n6_cascade_\ : std_logic;
signal \receive_module.rx_counter.X_7\ : std_logic;
signal \receive_module.rx_counter.n3385\ : std_logic;
signal \receive_module.rx_counter.old_HS\ : std_logic;
signal \TVP_HSYNC_buff\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \receive_module.n3091\ : std_logic;
signal \receive_module.n3092\ : std_logic;
signal \receive_module.n3093\ : std_logic;
signal \receive_module.n3094\ : std_logic;
signal \receive_module.n3095\ : std_logic;
signal \receive_module.n3096\ : std_logic;
signal \receive_module.n3097\ : std_logic;
signal \receive_module.n3098\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \receive_module.n3099\ : std_logic;
signal \receive_module.n3100\ : std_logic;
signal \receive_module.n3101\ : std_logic;
signal \receive_module.n3102\ : std_logic;
signal \receive_module.n3103\ : std_logic;
signal \receive_module.n3632\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_53\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_52\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_56\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_55\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_54\ : std_logic;
signal \transmit_module.video_signal_controller.n3629_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2901\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3125\ : std_logic;
signal \transmit_module.video_signal_controller.n3126\ : std_logic;
signal \transmit_module.video_signal_controller.n3127\ : std_logic;
signal \transmit_module.video_signal_controller.n3128\ : std_logic;
signal \transmit_module.video_signal_controller.n3129\ : std_logic;
signal \transmit_module.video_signal_controller.n3130\ : std_logic;
signal \transmit_module.video_signal_controller.n3131\ : std_logic;
signal \transmit_module.video_signal_controller.n3132\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3133\ : std_logic;
signal \transmit_module.video_signal_controller.n3134\ : std_logic;
signal \transmit_module.video_signal_controller.n3135\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_6\ : std_logic;
signal \receive_module.n131\ : std_logic;
signal \RX_ADDR_5\ : std_logic;
signal \receive_module.n130\ : std_logic;
signal \RX_ADDR_6\ : std_logic;
signal \receive_module.n129\ : std_logic;
signal \RX_ADDR_7\ : std_logic;
signal \receive_module.n128\ : std_logic;
signal \RX_ADDR_8\ : std_logic;
signal \receive_module.n127\ : std_logic;
signal \RX_ADDR_9\ : std_logic;
signal \receive_module.n136\ : std_logic;
signal \RX_ADDR_0\ : std_logic;
signal \receive_module.n135\ : std_logic;
signal \RX_ADDR_1\ : std_logic;
signal \line_buffer.n593\ : std_logic;
signal \line_buffer.n585\ : std_logic;
signal \receive_module.n126\ : std_logic;
signal \RX_ADDR_10\ : std_logic;
signal \receive_module.n133\ : std_logic;
signal \RX_ADDR_3\ : std_logic;
signal \receive_module.n132\ : std_logic;
signal \RX_ADDR_4\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_2\ : std_logic;
signal \RX_DATA_0\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \receive_module.rx_counter.n3156\ : std_logic;
signal \receive_module.rx_counter.n3157\ : std_logic;
signal \receive_module.rx_counter.n3158\ : std_logic;
signal \receive_module.rx_counter.n3159\ : std_logic;
signal \receive_module.rx_counter.n3160\ : std_logic;
signal \receive_module.rx_counter.n3623\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_4\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_2\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_5\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_1\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_0\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_3\ : std_logic;
signal \receive_module.rx_counter.n3473_cascade_\ : std_logic;
signal \receive_module.rx_counter.n7\ : std_logic;
signal \receive_module.rx_counter.n11\ : std_logic;
signal \receive_module.rx_counter.old_VS\ : std_logic;
signal \receive_module.rx_counter.n11_cascade_\ : std_logic;
signal \receive_module.rx_counter.n2529\ : std_logic;
signal \receive_module.rx_counter.n4_adj_605\ : std_logic;
signal \receive_module.rx_counter.n3422_cascade_\ : std_logic;
signal \receive_module.rx_counter.n55_adj_606\ : std_logic;
signal \receive_module.rx_counter.n3394\ : std_logic;
signal \receive_module.rx_counter.n5\ : std_logic;
signal \receive_module.rx_counter.n3413\ : std_logic;
signal \line_buffer.n596\ : std_logic;
signal \receive_module.rx_counter.n4_adj_604\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \receive_module.rx_counter.n3117\ : std_logic;
signal \receive_module.rx_counter.n3118\ : std_logic;
signal \receive_module.rx_counter.n3119\ : std_logic;
signal \receive_module.rx_counter.n3120\ : std_logic;
signal \receive_module.rx_counter.Y_5\ : std_logic;
signal \receive_module.rx_counter.n3121\ : std_logic;
signal \receive_module.rx_counter.Y_6\ : std_logic;
signal \receive_module.rx_counter.n3122\ : std_logic;
signal \receive_module.rx_counter.n3123\ : std_logic;
signal \receive_module.rx_counter.n3124\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \receive_module.rx_counter.n2063\ : std_logic;
signal \receive_module.n134\ : std_logic;
signal \TVP_VSYNC_buff\ : std_logic;
signal \RX_ADDR_2\ : std_logic;
signal \receive_module.n3631\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3136\ : std_logic;
signal \transmit_module.video_signal_controller.n3137\ : std_logic;
signal \transmit_module.video_signal_controller.n3138\ : std_logic;
signal \transmit_module.video_signal_controller.n3139\ : std_logic;
signal \transmit_module.video_signal_controller.n3140\ : std_logic;
signal \transmit_module.video_signal_controller.n3141\ : std_logic;
signal \transmit_module.video_signal_controller.n3142\ : std_logic;
signal \transmit_module.video_signal_controller.n3143\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3144\ : std_logic;
signal \transmit_module.video_signal_controller.n3145\ : std_logic;
signal \transmit_module.video_signal_controller.n3146\ : std_logic;
signal \line_buffer.n564\ : std_logic;
signal \transmit_module.video_signal_controller.n3624\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_2\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_1\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_0\ : std_logic;
signal \transmit_module.video_signal_controller.n2001\ : std_logic;
signal \transmit_module.video_signal_controller.n2917_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3313\ : std_logic;
signal \transmit_module.video_signal_controller.n2947_cascade_\ : std_logic;
signal \line_buffer.n522\ : std_logic;
signal \line_buffer.n530\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_3\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_5\ : std_logic;
signal \transmit_module.video_signal_controller.n18\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_9\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_10\ : std_logic;
signal \transmit_module.video_signal_controller.n4\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_7\ : std_logic;
signal \transmit_module.video_signal_controller.n3625_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_4\ : std_logic;
signal \line_buffer.n597\ : std_logic;
signal \line_buffer.n594\ : std_logic;
signal \line_buffer.n586\ : std_logic;
signal \line_buffer.n3591\ : std_logic;
signal \line_buffer.n468\ : std_logic;
signal n25 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_3\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_4\ : std_logic;
signal \receive_module.rx_counter.Y_4\ : std_logic;
signal \receive_module.rx_counter.Y_7\ : std_logic;
signal \receive_module.rx_counter.Y_1\ : std_logic;
signal \receive_module.rx_counter.Y_3\ : std_logic;
signal \receive_module.rx_counter.Y_2\ : std_logic;
signal \receive_module.rx_counter.Y_8\ : std_logic;
signal \receive_module.rx_counter.n10_adj_610\ : std_logic;
signal \receive_module.rx_counter.Y_0\ : std_logic;
signal \receive_module.rx_counter.n14_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3633\ : std_logic;
signal \RX_TX_SYNC\ : std_logic;
signal \sync_buffer.BUFFER_0_0\ : std_logic;
signal \RX_ADDR_12\ : std_logic;
signal \RX_WE\ : std_logic;
signal \RX_ADDR_13\ : std_logic;
signal \RX_ADDR_11\ : std_logic;
signal \line_buffer.n532\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_3\ : std_logic;
signal \RX_DATA_1\ : std_logic;
signal \sync_buffer.BUFFER_1_0\ : std_logic;
signal \RX_TX_SYNC_BUFF\ : std_logic;
signal \transmit_module.video_signal_controller.n2036\ : std_logic;
signal \transmit_module.video_signal_controller.n2378\ : std_logic;
signal \transmit_module.video_signal_controller.n49_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_1\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_0\ : std_logic;
signal \transmit_module.n113\ : std_logic;
signal \transmit_module.n142_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n45\ : std_logic;
signal \transmit_module.video_signal_controller.n3412\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_8\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_7\ : std_logic;
signal \transmit_module.video_signal_controller.n3626\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_6\ : std_logic;
signal \transmit_module.video_signal_controller.n3626_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_11\ : std_logic;
signal \transmit_module.n137_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_5\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_3\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_4\ : std_logic;
signal \transmit_module.video_signal_controller.n3628\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_9\ : std_logic;
signal \transmit_module.video_signal_controller.n3331\ : std_logic;
signal \transmit_module.video_signal_controller.n7_adj_618_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3622\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_VISIBLE_N_580_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_10\ : std_logic;
signal \transmit_module.video_signal_controller.n3477\ : std_logic;
signal \transmit_module.video_signal_controller.n16\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_2\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_8\ : std_logic;
signal \transmit_module.video_signal_controller.n3471\ : std_logic;
signal \transmit_module.video_signal_controller.n4_adj_617\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_6\ : std_logic;
signal \transmit_module.n144\ : std_logic;
signal \transmit_module.n3636\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_0\ : std_logic;
signal \transmit_module.old_VGA_HS\ : std_logic;
signal \transmit_module.VGA_VISIBLE_Y\ : std_logic;
signal \ADV_HSYNC_c\ : std_logic;
signal \transmit_module.n137\ : std_logic;
signal n18 : std_logic;
signal \transmit_module.n116\ : std_logic;
signal \transmit_module.n147\ : std_logic;
signal n28 : std_logic;
signal \transmit_module.n115\ : std_logic;
signal \transmit_module.n146\ : std_logic;
signal n27 : std_logic;
signal \DEBUG_c_3_c\ : std_logic;
signal \DEBUG_c_4_c\ : std_logic;
signal \DEBUG_c_5_c\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_7\ : std_logic;
signal \transmit_module.TX_ADDR_0\ : std_logic;
signal \transmit_module.n132\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \transmit_module.n131\ : std_logic;
signal \transmit_module.n3104\ : std_logic;
signal \transmit_module.n3105\ : std_logic;
signal \transmit_module.TX_ADDR_3\ : std_logic;
signal \transmit_module.n129\ : std_logic;
signal \transmit_module.n3106\ : std_logic;
signal \transmit_module.n3107\ : std_logic;
signal \transmit_module.n127\ : std_logic;
signal \transmit_module.n3108\ : std_logic;
signal \transmit_module.n3109\ : std_logic;
signal \transmit_module.n3110\ : std_logic;
signal \transmit_module.n3111\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \transmit_module.n3112\ : std_logic;
signal \transmit_module.n122\ : std_logic;
signal \transmit_module.n3113\ : std_logic;
signal \transmit_module.n3114\ : std_logic;
signal \transmit_module.n3115\ : std_logic;
signal \transmit_module.n3116\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_5\ : std_logic;
signal \transmit_module.TX_ADDR_5\ : std_logic;
signal \transmit_module.n111\ : std_logic;
signal \transmit_module.n111_cascade_\ : std_logic;
signal \transmit_module.n142\ : std_logic;
signal n23 : std_logic;
signal \transmit_module.video_signal_controller.VGA_VISIBLE_N_580\ : std_logic;
signal \transmit_module.video_signal_controller.n3333\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_11\ : std_logic;
signal \transmit_module.video_signal_controller.n7\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_10\ : std_logic;
signal \transmit_module.TX_ADDR_10\ : std_logic;
signal \transmit_module.n106\ : std_logic;
signal \transmit_module.n120\ : std_logic;
signal \transmit_module.n121\ : std_logic;
signal \transmit_module.n119\ : std_logic;
signal \transmit_module.n2057\ : std_logic;
signal \transmit_module.n124\ : std_logic;
signal \transmit_module.n126\ : std_logic;
signal \transmit_module.n123\ : std_logic;
signal \transmit_module.n125\ : std_logic;
signal n22 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_8\ : std_logic;
signal \transmit_module.TX_ADDR_8\ : std_logic;
signal n21 : std_logic;
signal \transmit_module.TX_ADDR_1\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_1\ : std_logic;
signal \transmit_module.n128\ : std_logic;
signal \transmit_module.n143\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \RX_DATA_3\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_5\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_5\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_6\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_6\ : std_logic;
signal \RX_DATA_4\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_7\ : std_logic;
signal \RX_DATA_5\ : std_logic;
signal \RX_DATA_6\ : std_logic;
signal \DEBUG_c_6_c\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_8\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_8\ : std_logic;
signal \transmit_module.n141\ : std_logic;
signal \transmit_module.n2167\ : std_logic;
signal \transmit_module.n140\ : std_logic;
signal \transmit_module.n130\ : std_logic;
signal \transmit_module.n145_cascade_\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_16\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_17\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_20\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_19\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_18\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_13\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_12\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_11\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.n108\ : std_logic;
signal \transmit_module.n139\ : std_logic;
signal n20 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_7\ : std_logic;
signal \transmit_module.TX_ADDR_7\ : std_logic;
signal \transmit_module.n109\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_6\ : std_logic;
signal \transmit_module.TX_ADDR_6\ : std_logic;
signal \transmit_module.n110\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_2\ : std_logic;
signal \transmit_module.TX_ADDR_2\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_9\ : std_logic;
signal \transmit_module.TX_ADDR_9\ : std_logic;
signal \transmit_module.n107\ : std_logic;
signal \transmit_module.n107_cascade_\ : std_logic;
signal \transmit_module.n138\ : std_logic;
signal n19 : std_logic;
signal \transmit_module.n114\ : std_logic;
signal \transmit_module.n145\ : std_logic;
signal n26 : std_logic;
signal \tvp_video_buffer.BUFFER_1_4\ : std_logic;
signal \RX_DATA_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.n3627\ : std_logic;
signal \line_buffer.n556\ : std_logic;
signal \line_buffer.n548\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.n112\ : std_logic;
signal \transmit_module.TX_ADDR_4\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_4\ : std_logic;
signal \transmit_module.n2069\ : std_logic;
signal \ADV_VSYNC_c\ : std_logic;
signal \line_buffer.n529\ : std_logic;
signal \line_buffer.n521\ : std_logic;
signal \line_buffer.n3500_cascade_\ : std_logic;
signal \line_buffer.n3501\ : std_logic;
signal \line_buffer.n3537_cascade_\ : std_logic;
signal \line_buffer.n464\ : std_logic;
signal \line_buffer.n456\ : std_logic;
signal \line_buffer.n3497\ : std_logic;
signal \line_buffer.n524\ : std_logic;
signal \line_buffer.n516\ : std_logic;
signal \line_buffer.n560\ : std_logic;
signal \line_buffer.n552\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.n2115\ : std_logic;
signal \transmit_module.n3635\ : std_logic;
signal \line_buffer.n463\ : std_logic;
signal \line_buffer.n455\ : std_logic;
signal \line_buffer.n3525\ : std_logic;
signal \line_buffer.n3524_cascade_\ : std_logic;
signal \line_buffer.n3521\ : std_logic;
signal \line_buffer.n3555_cascade_\ : std_logic;
signal \line_buffer.n3519\ : std_logic;
signal \line_buffer.n561\ : std_logic;
signal \line_buffer.n553\ : std_logic;
signal \line_buffer.n3498\ : std_logic;
signal \line_buffer.n587\ : std_logic;
signal \line_buffer.n579\ : std_logic;
signal n1814 : std_logic;
signal \TX_DATA_1\ : std_logic;
signal n1813 : std_logic;
signal \TX_DATA_5\ : std_logic;
signal n1809 : std_logic;
signal \TX_DATA_6\ : std_logic;
signal n1808 : std_logic;
signal \line_buffer.n528\ : std_logic;
signal \line_buffer.n520\ : std_logic;
signal \line_buffer.n3594\ : std_logic;
signal \line_buffer.n592\ : std_logic;
signal \line_buffer.n584\ : std_logic;
signal \line_buffer.n3489\ : std_logic;
signal \line_buffer.n3488\ : std_logic;
signal \line_buffer.n3561\ : std_logic;
signal \line_buffer.n591\ : std_logic;
signal \line_buffer.n583\ : std_logic;
signal \line_buffer.n523\ : std_logic;
signal \line_buffer.n515\ : std_logic;
signal \line_buffer.n3597\ : std_logic;
signal \line_buffer.n3600_cascade_\ : std_logic;
signal \TX_DATA_0\ : std_logic;
signal \transmit_module.VGA_VISIBLE\ : std_logic;
signal \TX_DATA_7\ : std_logic;
signal \ADV_B_c\ : std_logic;
signal \RX_DATA_7\ : std_logic;
signal \line_buffer.n465\ : std_logic;
signal \line_buffer.n457\ : std_logic;
signal \line_buffer.n3588\ : std_logic;
signal \line_buffer.n557\ : std_logic;
signal \line_buffer.n549\ : std_logic;
signal \line_buffer.n460\ : std_logic;
signal \line_buffer.n452\ : std_logic;
signal \line_buffer.n3549\ : std_logic;
signal \line_buffer.n3552_cascade_\ : std_logic;
signal \line_buffer.n527\ : std_logic;
signal \line_buffer.n519\ : std_logic;
signal \line_buffer.n3573\ : std_logic;
signal \line_buffer.n589\ : std_logic;
signal \line_buffer.n581\ : std_logic;
signal \line_buffer.n517\ : std_logic;
signal \line_buffer.n525\ : std_logic;
signal \line_buffer.n3603_cascade_\ : std_logic;
signal \line_buffer.n3606\ : std_logic;
signal \line_buffer.n462\ : std_logic;
signal \line_buffer.n454\ : std_logic;
signal \line_buffer.n3546_cascade_\ : std_logic;
signal \line_buffer.n3576\ : std_logic;
signal \line_buffer.n555\ : std_logic;
signal \line_buffer.n547\ : std_logic;
signal \line_buffer.n461\ : std_logic;
signal \line_buffer.n453\ : std_logic;
signal \line_buffer.n588\ : std_logic;
signal \line_buffer.n580\ : std_logic;
signal \line_buffer.n3522\ : std_logic;
signal \line_buffer.n458\ : std_logic;
signal \line_buffer.n450\ : std_logic;
signal \line_buffer.n3579\ : std_logic;
signal \line_buffer.n3582\ : std_logic;
signal \TX_DATA_2\ : std_logic;
signal n1812 : std_logic;
signal \TX_DATA_4\ : std_logic;
signal n1810 : std_logic;
signal \line_buffer.n554\ : std_logic;
signal \line_buffer.n562\ : std_logic;
signal \line_buffer.n3585\ : std_logic;
signal \line_buffer.n558\ : std_logic;
signal \line_buffer.n550\ : std_logic;
signal \TX_ADDR_13\ : std_logic;
signal \line_buffer.n3482\ : std_logic;
signal \line_buffer.n3567_cascade_\ : std_logic;
signal \line_buffer.n3483\ : std_logic;
signal \line_buffer.n559\ : std_logic;
signal \TX_ADDR_12\ : std_logic;
signal \line_buffer.n551\ : std_logic;
signal \line_buffer.n3543\ : std_logic;
signal \line_buffer.n582\ : std_logic;
signal \line_buffer.n590\ : std_logic;
signal \line_buffer.n3480\ : std_logic;
signal \TX_DATA_3\ : std_logic;
signal n1811 : std_logic;
signal \ADV_CLK_c\ : std_logic;
signal \transmit_module.n2367\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_9\ : std_logic;
signal \line_buffer.n526\ : std_logic;
signal \line_buffer.n518\ : std_logic;
signal \line_buffer.n3479\ : std_logic;
signal \DEBUG_c_7_c\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_9\ : std_logic;
signal \DEBUG_c_2_c\ : std_logic;
signal \line_buffer.n459\ : std_logic;
signal \line_buffer.n451\ : std_logic;
signal \TX_ADDR_11\ : std_logic;
signal \line_buffer.n3518\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \TVP_CLK_wire\ : std_logic;
signal \ADV_CLK_wire\ : std_logic;
signal \TVP_VIDEO_wire\ : std_logic_vector(9 downto 0);
signal \ADV_G_wire\ : std_logic_vector(7 downto 0);
signal \ADV_R_wire\ : std_logic_vector(7 downto 0);
signal \ADV_B_wire\ : std_logic_vector(7 downto 0);
signal \ADV_SYNC_N_wire\ : std_logic;
signal \ADV_BLANK_N_wire\ : std_logic;
signal \TVP_HSYNC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \ADV_HSYNC_wire\ : std_logic;
signal \TVP_VSYNC_wire\ : std_logic;
signal \ADV_VSYNC_wire\ : std_logic;
signal \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \line_buffer.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \TVP_CLK_wire\ <= TVP_CLK;
    ADV_CLK <= \ADV_CLK_wire\;
    \TVP_VIDEO_wire\ <= TVP_VIDEO;
    ADV_G <= \ADV_G_wire\;
    ADV_R <= \ADV_R_wire\;
    ADV_B <= \ADV_B_wire\;
    ADV_SYNC_N <= \ADV_SYNC_N_wire\;
    ADV_BLANK_N <= \ADV_BLANK_N_wire\;
    \TVP_HSYNC_wire\ <= TVP_HSYNC;
    LED <= \LED_wire\;
    ADV_HSYNC <= \ADV_HSYNC_wire\;
    \TVP_VSYNC_wire\ <= TVP_VSYNC;
    ADV_VSYNC <= \ADV_VSYNC_wire\;
    \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.n465\ <= \line_buffer.mem2_physical_RDATA_wire\(11);
    \line_buffer.n464\ <= \line_buffer.mem2_physical_RDATA_wire\(3);
    \line_buffer.mem2_physical_RADDR_wire\ <= \N__16186\&\N__18964\&\N__19420\&\N__17104\&\N__17374\&\N__16837\&\N__9121\&\N__14008\&\N__18712\&\N__15670\&\N__15922\;
    \line_buffer.mem2_physical_WADDR_wire\ <= \N__12349\&\N__10438\&\N__10681\&\N__10936\&\N__11194\&\N__11452\&\N__11833\&\N__12091\&\N__12892\&\N__9922\&\N__10183\;
    \line_buffer.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22154\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18559\&'0'&'0'&'0';
    \line_buffer.n552\ <= \line_buffer.mem14_physical_RDATA_wire\(11);
    \line_buffer.n551\ <= \line_buffer.mem14_physical_RDATA_wire\(3);
    \line_buffer.mem14_physical_RADDR_wire\ <= \N__16258\&\N__19036\&\N__19492\&\N__17176\&\N__17446\&\N__16909\&\N__9193\&\N__14080\&\N__18784\&\N__15742\&\N__15994\;
    \line_buffer.mem14_physical_WADDR_wire\ <= \N__12421\&\N__10510\&\N__10753\&\N__11008\&\N__11266\&\N__11524\&\N__11905\&\N__12163\&\N__12964\&\N__9994\&\N__10255\;
    \line_buffer.mem14_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem14_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17671\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17762\&'0'&'0'&'0';
    \line_buffer.n562\ <= \line_buffer.mem5_physical_RDATA_wire\(11);
    \line_buffer.n561\ <= \line_buffer.mem5_physical_RDATA_wire\(3);
    \line_buffer.mem5_physical_RADDR_wire\ <= \N__16189\&\N__18985\&\N__19435\&\N__17113\&\N__17377\&\N__16840\&\N__9124\&\N__13999\&\N__18721\&\N__15679\&\N__15937\;
    \line_buffer.mem5_physical_WADDR_wire\ <= \N__12340\&\N__10441\&\N__10696\&\N__10945\&\N__11203\&\N__11467\&\N__11830\&\N__12088\&\N__12913\&\N__9937\&\N__10192\;
    \line_buffer.mem5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22148\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18561\&'0'&'0'&'0';
    \line_buffer.n520\ <= \line_buffer.mem11_physical_RDATA_wire\(11);
    \line_buffer.n519\ <= \line_buffer.mem11_physical_RDATA_wire\(3);
    \line_buffer.mem11_physical_RADDR_wire\ <= \N__16294\&\N__19072\&\N__19528\&\N__17212\&\N__17482\&\N__16945\&\N__9229\&\N__14116\&\N__18820\&\N__15778\&\N__16030\;
    \line_buffer.mem11_physical_WADDR_wire\ <= \N__12457\&\N__10546\&\N__10789\&\N__11044\&\N__11302\&\N__11560\&\N__11941\&\N__12199\&\N__13000\&\N__10030\&\N__10291\;
    \line_buffer.mem11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem11_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17654\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17761\&'0'&'0'&'0';
    \line_buffer.n582\ <= \line_buffer.mem21_physical_RDATA_wire\(11);
    \line_buffer.n581\ <= \line_buffer.mem21_physical_RDATA_wire\(3);
    \line_buffer.mem21_physical_RADDR_wire\ <= \N__16162\&\N__18940\&\N__19396\&\N__17080\&\N__17350\&\N__16813\&\N__9097\&\N__13984\&\N__18688\&\N__15646\&\N__15898\;
    \line_buffer.mem21_physical_WADDR_wire\ <= \N__12325\&\N__10414\&\N__10657\&\N__10912\&\N__11170\&\N__11428\&\N__11809\&\N__12067\&\N__12868\&\N__9898\&\N__10159\;
    \line_buffer.mem21_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem21_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17911\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19755\&'0'&'0'&'0';
    \line_buffer.n518\ <= \line_buffer.mem12_physical_RDATA_wire\(11);
    \line_buffer.n517\ <= \line_buffer.mem12_physical_RDATA_wire\(3);
    \line_buffer.mem12_physical_RADDR_wire\ <= \N__16282\&\N__19060\&\N__19516\&\N__17200\&\N__17470\&\N__16933\&\N__9217\&\N__14104\&\N__18808\&\N__15766\&\N__16018\;
    \line_buffer.mem12_physical_WADDR_wire\ <= \N__12445\&\N__10534\&\N__10777\&\N__11032\&\N__11290\&\N__11548\&\N__11929\&\N__12187\&\N__12988\&\N__10018\&\N__10279\;
    \line_buffer.mem12_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem12_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17886\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19742\&'0'&'0'&'0';
    \line_buffer.n526\ <= \line_buffer.mem24_physical_RDATA_wire\(11);
    \line_buffer.n525\ <= \line_buffer.mem24_physical_RDATA_wire\(3);
    \line_buffer.mem24_physical_RADDR_wire\ <= \N__16309\&\N__19105\&\N__19555\&\N__17233\&\N__17497\&\N__16960\&\N__9244\&\N__14119\&\N__18841\&\N__15799\&\N__16057\;
    \line_buffer.mem24_physical_WADDR_wire\ <= \N__12460\&\N__10561\&\N__10816\&\N__11065\&\N__11323\&\N__11587\&\N__11950\&\N__12208\&\N__13033\&\N__10057\&\N__10312\;
    \line_buffer.mem24_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem24_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17882\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19765\&'0'&'0'&'0';
    \line_buffer.n554\ <= \line_buffer.mem1_physical_RDATA_wire\(11);
    \line_buffer.n553\ <= \line_buffer.mem1_physical_RDATA_wire\(3);
    \line_buffer.mem1_physical_RADDR_wire\ <= \N__16318\&\N__19096\&\N__19552\&\N__17236\&\N__17506\&\N__16969\&\N__9253\&\N__14135\&\N__18844\&\N__15802\&\N__16054\;
    \line_buffer.mem1_physical_WADDR_wire\ <= \N__12476\&\N__10570\&\N__10813\&\N__11068\&\N__11326\&\N__11584\&\N__11963\&\N__12221\&\N__13024\&\N__10054\&\N__10315\;
    \line_buffer.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22132\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18540\&'0'&'0'&'0';
    \line_buffer.n550\ <= \line_buffer.mem15_physical_RDATA_wire\(11);
    \line_buffer.n549\ <= \line_buffer.mem15_physical_RDATA_wire\(3);
    \line_buffer.mem15_physical_RADDR_wire\ <= \N__16246\&\N__19024\&\N__19480\&\N__17164\&\N__17434\&\N__16897\&\N__9181\&\N__14068\&\N__18772\&\N__15730\&\N__15982\;
    \line_buffer.mem15_physical_WADDR_wire\ <= \N__12409\&\N__10498\&\N__10741\&\N__10996\&\N__11254\&\N__11512\&\N__11893\&\N__12151\&\N__12952\&\N__9982\&\N__10243\;
    \line_buffer.mem15_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem15_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17913\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19770\&'0'&'0'&'0';
    \line_buffer.n558\ <= \line_buffer.mem27_physical_RDATA_wire\(11);
    \line_buffer.n557\ <= \line_buffer.mem27_physical_RDATA_wire\(3);
    \line_buffer.mem27_physical_RADDR_wire\ <= \N__16273\&\N__19069\&\N__19519\&\N__17197\&\N__17461\&\N__16924\&\N__9208\&\N__14083\&\N__18805\&\N__15763\&\N__16021\;
    \line_buffer.mem27_physical_WADDR_wire\ <= \N__12424\&\N__10525\&\N__10780\&\N__11029\&\N__11287\&\N__11551\&\N__11914\&\N__12172\&\N__12997\&\N__10021\&\N__10276\;
    \line_buffer.mem27_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem27_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17912\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19748\&'0'&'0'&'0';
    \line_buffer.n530\ <= \line_buffer.mem4_physical_RDATA_wire\(11);
    \line_buffer.n529\ <= \line_buffer.mem4_physical_RDATA_wire\(3);
    \line_buffer.mem4_physical_RADDR_wire\ <= \N__16201\&\N__18997\&\N__19447\&\N__17125\&\N__17389\&\N__16852\&\N__9136\&\N__14011\&\N__18733\&\N__15691\&\N__15949\;
    \line_buffer.mem4_physical_WADDR_wire\ <= \N__12352\&\N__10453\&\N__10708\&\N__10957\&\N__11215\&\N__11479\&\N__11842\&\N__12100\&\N__12925\&\N__9949\&\N__10204\;
    \line_buffer.mem4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22135\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18560\&'0'&'0'&'0';
    \line_buffer.n548\ <= \line_buffer.mem16_physical_RDATA_wire\(11);
    \line_buffer.n547\ <= \line_buffer.mem16_physical_RDATA_wire\(3);
    \line_buffer.mem16_physical_RADDR_wire\ <= \N__16234\&\N__19012\&\N__19468\&\N__17152\&\N__17422\&\N__16885\&\N__9169\&\N__14056\&\N__18760\&\N__15718\&\N__15970\;
    \line_buffer.mem16_physical_WADDR_wire\ <= \N__12397\&\N__10486\&\N__10729\&\N__10984\&\N__11242\&\N__11500\&\N__11881\&\N__12139\&\N__12940\&\N__9970\&\N__10231\;
    \line_buffer.mem16_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem16_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14334\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11716\&'0'&'0'&'0';
    \line_buffer.n590\ <= \line_buffer.mem30_physical_RDATA_wire\(11);
    \line_buffer.n589\ <= \line_buffer.mem30_physical_RDATA_wire\(3);
    \line_buffer.mem30_physical_RADDR_wire\ <= \N__16225\&\N__19021\&\N__19471\&\N__17149\&\N__17413\&\N__16876\&\N__9160\&\N__14035\&\N__18757\&\N__15715\&\N__15973\;
    \line_buffer.mem30_physical_WADDR_wire\ <= \N__12376\&\N__10477\&\N__10732\&\N__10981\&\N__11239\&\N__11503\&\N__11866\&\N__12124\&\N__12949\&\N__9973\&\N__10228\;
    \line_buffer.mem30_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem30_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17892\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19766\&'0'&'0'&'0';
    \line_buffer.n457\ <= \line_buffer.mem7_physical_RDATA_wire\(11);
    \line_buffer.n456\ <= \line_buffer.mem7_physical_RDATA_wire\(3);
    \line_buffer.mem7_physical_RADDR_wire\ <= \N__16165\&\N__18961\&\N__19411\&\N__17089\&\N__17353\&\N__16816\&\N__9100\&\N__13975\&\N__18697\&\N__15655\&\N__15913\;
    \line_buffer.mem7_physical_WADDR_wire\ <= \N__12316\&\N__10417\&\N__10672\&\N__10921\&\N__11179\&\N__11443\&\N__11806\&\N__12064\&\N__12889\&\N__9913\&\N__10168\;
    \line_buffer.mem7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem7_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22150\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18569\&'0'&'0'&'0';
    \line_buffer.n584\ <= \line_buffer.mem20_physical_RDATA_wire\(11);
    \line_buffer.n583\ <= \line_buffer.mem20_physical_RDATA_wire\(3);
    \line_buffer.mem20_physical_RADDR_wire\ <= \N__16174\&\N__18952\&\N__19408\&\N__17092\&\N__17362\&\N__16825\&\N__9109\&\N__13996\&\N__18700\&\N__15658\&\N__15910\;
    \line_buffer.mem20_physical_WADDR_wire\ <= \N__12337\&\N__10426\&\N__10669\&\N__10924\&\N__11182\&\N__11440\&\N__11821\&\N__12079\&\N__12880\&\N__9910\&\N__10171\;
    \line_buffer.mem20_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem20_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17672\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17788\&'0'&'0'&'0';
    \line_buffer.n516\ <= \line_buffer.mem13_physical_RDATA_wire\(11);
    \line_buffer.n515\ <= \line_buffer.mem13_physical_RDATA_wire\(3);
    \line_buffer.mem13_physical_RADDR_wire\ <= \N__16270\&\N__19048\&\N__19504\&\N__17188\&\N__17458\&\N__16921\&\N__9205\&\N__14092\&\N__18796\&\N__15754\&\N__16006\;
    \line_buffer.mem13_physical_WADDR_wire\ <= \N__12433\&\N__10522\&\N__10765\&\N__11020\&\N__11278\&\N__11536\&\N__11917\&\N__12175\&\N__12976\&\N__10006\&\N__10267\;
    \line_buffer.mem13_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem13_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14327\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11699\&'0'&'0'&'0';
    \line_buffer.n459\ <= \line_buffer.mem19_physical_RDATA_wire\(11);
    \line_buffer.n458\ <= \line_buffer.mem19_physical_RDATA_wire\(3);
    \line_buffer.mem19_physical_RADDR_wire\ <= \N__16198\&\N__18976\&\N__19432\&\N__17116\&\N__17386\&\N__16849\&\N__9133\&\N__14020\&\N__18724\&\N__15682\&\N__15934\;
    \line_buffer.mem19_physical_WADDR_wire\ <= \N__12361\&\N__10450\&\N__10693\&\N__10948\&\N__11206\&\N__11464\&\N__11845\&\N__12103\&\N__12904\&\N__9934\&\N__10195\;
    \line_buffer.mem19_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem19_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14335\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11717\&'0'&'0'&'0';
    \line_buffer.n528\ <= \line_buffer.mem23_physical_RDATA_wire\(11);
    \line_buffer.n527\ <= \line_buffer.mem23_physical_RDATA_wire\(3);
    \line_buffer.mem23_physical_RADDR_wire\ <= \N__16321\&\N__19112\&\N__19565\&\N__17245\&\N__17509\&\N__16972\&\N__9256\&\N__14131\&\N__18853\&\N__15811\&\N__16067\;
    \line_buffer.mem23_physical_WADDR_wire\ <= \N__12472\&\N__10573\&\N__10826\&\N__11077\&\N__11335\&\N__11597\&\N__11962\&\N__12220\&\N__13040\&\N__10067\&\N__10324\;
    \line_buffer.mem23_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem23_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17677\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17770\&'0'&'0'&'0';
    \line_buffer.n522\ <= \line_buffer.mem0_physical_RDATA_wire\(11);
    \line_buffer.n521\ <= \line_buffer.mem0_physical_RDATA_wire\(3);
    \line_buffer.mem0_physical_RADDR_wire\ <= \N__16325\&\N__19108\&\N__19564\&\N__17246\&\N__17513\&\N__16976\&\N__9260\&\N__14141\&\N__18854\&\N__15812\&\N__16066\;
    \line_buffer.mem0_physical_WADDR_wire\ <= \N__12482\&\N__10577\&\N__10825\&\N__11078\&\N__11336\&\N__11596\&\N__11969\&\N__12227\&\N__13036\&\N__10066\&\N__10325\;
    \line_buffer.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22133\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18558\&'0'&'0'&'0';
    \line_buffer.n560\ <= \line_buffer.mem26_physical_RDATA_wire\(11);
    \line_buffer.n559\ <= \line_buffer.mem26_physical_RDATA_wire\(3);
    \line_buffer.mem26_physical_RADDR_wire\ <= \N__16285\&\N__19081\&\N__19531\&\N__17209\&\N__17473\&\N__16936\&\N__9220\&\N__14095\&\N__18817\&\N__15775\&\N__16033\;
    \line_buffer.mem26_physical_WADDR_wire\ <= \N__12436\&\N__10537\&\N__10792\&\N__11041\&\N__11299\&\N__11563\&\N__11926\&\N__12184\&\N__13009\&\N__10033\&\N__10288\;
    \line_buffer.mem26_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem26_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17645\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17774\&'0'&'0'&'0';
    \line_buffer.n586\ <= \line_buffer.mem3_physical_RDATA_wire\(11);
    \line_buffer.n585\ <= \line_buffer.mem3_physical_RDATA_wire\(3);
    \line_buffer.mem3_physical_RADDR_wire\ <= \N__16237\&\N__19033\&\N__19483\&\N__17161\&\N__17425\&\N__16888\&\N__9172\&\N__14047\&\N__18769\&\N__15727\&\N__15985\;
    \line_buffer.mem3_physical_WADDR_wire\ <= \N__12388\&\N__10489\&\N__10744\&\N__10993\&\N__11251\&\N__11515\&\N__11878\&\N__12136\&\N__12961\&\N__9985\&\N__10240\;
    \line_buffer.mem3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22134\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18532\&'0'&'0'&'0';
    \line_buffer.n463\ <= \line_buffer.mem17_physical_RDATA_wire\(11);
    \line_buffer.n462\ <= \line_buffer.mem17_physical_RDATA_wire\(3);
    \line_buffer.mem17_physical_RADDR_wire\ <= \N__16222\&\N__19000\&\N__19456\&\N__17140\&\N__17410\&\N__16873\&\N__9157\&\N__14044\&\N__18748\&\N__15706\&\N__15958\;
    \line_buffer.mem17_physical_WADDR_wire\ <= \N__12385\&\N__10474\&\N__10717\&\N__10972\&\N__11230\&\N__11488\&\N__11869\&\N__12127\&\N__12928\&\N__9958\&\N__10219\;
    \line_buffer.mem17_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem17_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17658\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17775\&'0'&'0'&'0';
    \line_buffer.n588\ <= \line_buffer.mem31_physical_RDATA_wire\(11);
    \line_buffer.n587\ <= \line_buffer.mem31_physical_RDATA_wire\(3);
    \line_buffer.mem31_physical_RADDR_wire\ <= \N__16213\&\N__19009\&\N__19459\&\N__17137\&\N__17401\&\N__16864\&\N__9148\&\N__14023\&\N__18745\&\N__15703\&\N__15961\;
    \line_buffer.mem31_physical_WADDR_wire\ <= \N__12364\&\N__10465\&\N__10720\&\N__10969\&\N__11227\&\N__11491\&\N__11854\&\N__12112\&\N__12937\&\N__9961\&\N__10216\;
    \line_buffer.mem31_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem31_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14348\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11721\&'0'&'0'&'0';
    \line_buffer.n453\ <= \line_buffer.mem9_physical_RDATA_wire\(11);
    \line_buffer.n452\ <= \line_buffer.mem9_physical_RDATA_wire\(3);
    \line_buffer.mem9_physical_RADDR_wire\ <= \N__16141\&\N__18937\&\N__19387\&\N__17065\&\N__17329\&\N__16792\&\N__9076\&\N__13951\&\N__18673\&\N__15631\&\N__15889\;
    \line_buffer.mem9_physical_WADDR_wire\ <= \N__12291\&\N__10393\&\N__10648\&\N__10897\&\N__11155\&\N__11419\&\N__11781\&\N__12039\&\N__12865\&\N__9889\&\N__10144\;
    \line_buffer.mem9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem9_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17924\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19778\&'0'&'0'&'0';
    \line_buffer.n592\ <= \line_buffer.mem29_physical_RDATA_wire\(11);
    \line_buffer.n591\ <= \line_buffer.mem29_physical_RDATA_wire\(3);
    \line_buffer.mem29_physical_RADDR_wire\ <= \N__16249\&\N__19045\&\N__19495\&\N__17173\&\N__17437\&\N__16900\&\N__9184\&\N__14059\&\N__18781\&\N__15739\&\N__15997\;
    \line_buffer.mem29_physical_WADDR_wire\ <= \N__12400\&\N__10501\&\N__10756\&\N__11005\&\N__11263\&\N__11527\&\N__11890\&\N__12148\&\N__12973\&\N__9997\&\N__10252\;
    \line_buffer.mem29_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem29_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17673\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17769\&'0'&'0'&'0';
    \line_buffer.n594\ <= \line_buffer.mem6_physical_RDATA_wire\(11);
    \line_buffer.n593\ <= \line_buffer.mem6_physical_RDATA_wire\(3);
    \line_buffer.mem6_physical_RADDR_wire\ <= \N__16177\&\N__18973\&\N__19423\&\N__17101\&\N__17365\&\N__16828\&\N__9112\&\N__13987\&\N__18709\&\N__15667\&\N__15925\;
    \line_buffer.mem6_physical_WADDR_wire\ <= \N__12328\&\N__10429\&\N__10684\&\N__10933\&\N__11191\&\N__11455\&\N__11818\&\N__12076\&\N__12901\&\N__9925\&\N__10180\;
    \line_buffer.mem6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22149\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18568\&'0'&'0'&'0';
    \line_buffer.n451\ <= \line_buffer.mem10_physical_RDATA_wire\(11);
    \line_buffer.n450\ <= \line_buffer.mem10_physical_RDATA_wire\(3);
    \line_buffer.mem10_physical_RADDR_wire\ <= \N__16306\&\N__19084\&\N__19540\&\N__17224\&\N__17494\&\N__16957\&\N__9241\&\N__14128\&\N__18832\&\N__15790\&\N__16042\;
    \line_buffer.mem10_physical_WADDR_wire\ <= \N__12469\&\N__10558\&\N__10801\&\N__11056\&\N__11314\&\N__11572\&\N__11953\&\N__12211\&\N__13012\&\N__10042\&\N__10303\;
    \line_buffer.mem10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem10_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14339\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11698\&'0'&'0'&'0';
    \line_buffer.n580\ <= \line_buffer.mem22_physical_RDATA_wire\(11);
    \line_buffer.n579\ <= \line_buffer.mem22_physical_RDATA_wire\(3);
    \line_buffer.mem22_physical_RADDR_wire\ <= \N__16150\&\N__18928\&\N__19384\&\N__17068\&\N__17338\&\N__16801\&\N__9085\&\N__13972\&\N__18676\&\N__15634\&\N__15886\;
    \line_buffer.mem22_physical_WADDR_wire\ <= \N__12313\&\N__10402\&\N__10645\&\N__10900\&\N__11158\&\N__11416\&\N__11797\&\N__12055\&\N__12856\&\N__9886\&\N__10147\;
    \line_buffer.mem22_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem22_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14346\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11723\&'0'&'0'&'0';
    \line_buffer.n524\ <= \line_buffer.mem25_physical_RDATA_wire\(11);
    \line_buffer.n523\ <= \line_buffer.mem25_physical_RDATA_wire\(3);
    \line_buffer.mem25_physical_RADDR_wire\ <= \N__16297\&\N__19093\&\N__19543\&\N__17221\&\N__17485\&\N__16948\&\N__9232\&\N__14107\&\N__18829\&\N__15787\&\N__16045\;
    \line_buffer.mem25_physical_WADDR_wire\ <= \N__12448\&\N__10549\&\N__10804\&\N__11053\&\N__11311\&\N__11575\&\N__11938\&\N__12196\&\N__13021\&\N__10045\&\N__10300\;
    \line_buffer.mem25_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem25_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14347\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11712\&'0'&'0'&'0';
    \line_buffer.n455\ <= \line_buffer.mem8_physical_RDATA_wire\(11);
    \line_buffer.n454\ <= \line_buffer.mem8_physical_RDATA_wire\(3);
    \line_buffer.mem8_physical_RADDR_wire\ <= \N__16153\&\N__18949\&\N__19399\&\N__17077\&\N__17341\&\N__16804\&\N__9088\&\N__13963\&\N__18685\&\N__15643\&\N__15901\;
    \line_buffer.mem8_physical_WADDR_wire\ <= \N__12304\&\N__10405\&\N__10660\&\N__10909\&\N__11167\&\N__11431\&\N__11794\&\N__12052\&\N__12877\&\N__9901\&\N__10156\;
    \line_buffer.mem8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem8_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17687\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17789\&'0'&'0'&'0';
    \line_buffer.n556\ <= \line_buffer.mem28_physical_RDATA_wire\(11);
    \line_buffer.n555\ <= \line_buffer.mem28_physical_RDATA_wire\(3);
    \line_buffer.mem28_physical_RADDR_wire\ <= \N__16261\&\N__19057\&\N__19507\&\N__17185\&\N__17449\&\N__16912\&\N__9196\&\N__14071\&\N__18793\&\N__15751\&\N__16009\;
    \line_buffer.mem28_physical_WADDR_wire\ <= \N__12412\&\N__10513\&\N__10768\&\N__11017\&\N__11275\&\N__11539\&\N__11902\&\N__12160\&\N__12985\&\N__10009\&\N__10264\;
    \line_buffer.mem28_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem28_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14305\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11722\&'0'&'0'&'0';
    \line_buffer.n461\ <= \line_buffer.mem18_physical_RDATA_wire\(11);
    \line_buffer.n460\ <= \line_buffer.mem18_physical_RDATA_wire\(3);
    \line_buffer.mem18_physical_RADDR_wire\ <= \N__16210\&\N__18988\&\N__19444\&\N__17128\&\N__17398\&\N__16861\&\N__9145\&\N__14032\&\N__18736\&\N__15694\&\N__15946\;
    \line_buffer.mem18_physical_WADDR_wire\ <= \N__12373\&\N__10462\&\N__10705\&\N__10960\&\N__11218\&\N__11476\&\N__11857\&\N__12115\&\N__12916\&\N__9946\&\N__10207\;
    \line_buffer.mem18_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem18_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17920\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19777\&'0'&'0'&'0';

    \tx_pll.TX_PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0100110",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \ADV_CLK_c\,
            REFERENCECLK => \N__8399\,
            RESETB => \N__18070\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \line_buffer.mem2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem2_physical_RDATA_wire\,
            RADDR => \line_buffer.mem2_physical_RADDR_wire\,
            WADDR => \line_buffer.mem2_physical_WADDR_wire\,
            MASK => \line_buffer.mem2_physical_MASK_wire\,
            WDATA => \line_buffer.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23228\,
            RE => \N__18072\,
            WCLKE => 'H',
            WCLK => \N__24625\,
            WE => \N__14183\
        );

    \line_buffer.mem14_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem14_physical_RDATA_wire\,
            RADDR => \line_buffer.mem14_physical_RADDR_wire\,
            WADDR => \line_buffer.mem14_physical_WADDR_wire\,
            MASK => \line_buffer.mem14_physical_MASK_wire\,
            WDATA => \line_buffer.mem14_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23483\,
            RE => \N__18170\,
            WCLKE => 'H',
            WCLK => \N__24611\,
            WE => \N__13374\
        );

    \line_buffer.mem5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem5_physical_RDATA_wire\,
            RADDR => \line_buffer.mem5_physical_RADDR_wire\,
            WADDR => \line_buffer.mem5_physical_WADDR_wire\,
            MASK => \line_buffer.mem5_physical_MASK_wire\,
            WDATA => \line_buffer.mem5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22710\,
            RE => \N__18051\,
            WCLKE => 'H',
            WCLK => \N__24624\,
            WE => \N__9647\
        );

    \line_buffer.mem11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem11_physical_RDATA_wire\,
            RADDR => \line_buffer.mem11_physical_RADDR_wire\,
            WADDR => \line_buffer.mem11_physical_WADDR_wire\,
            MASK => \line_buffer.mem11_physical_MASK_wire\,
            WDATA => \line_buffer.mem11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23320\,
            RE => \N__18197\,
            WCLKE => 'H',
            WCLK => \N__24601\,
            WE => \N__14395\
        );

    \line_buffer.mem21_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem21_physical_RDATA_wire\,
            RADDR => \line_buffer.mem21_physical_RADDR_wire\,
            WADDR => \line_buffer.mem21_physical_WADDR_wire\,
            MASK => \line_buffer.mem21_physical_MASK_wire\,
            WDATA => \line_buffer.mem21_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23057\,
            RE => \N__18089\,
            WCLKE => 'H',
            WCLK => \N__24631\,
            WE => \N__12691\
        );

    \line_buffer.mem12_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem12_physical_RDATA_wire\,
            RADDR => \line_buffer.mem12_physical_RADDR_wire\,
            WADDR => \line_buffer.mem12_physical_WADDR_wire\,
            MASK => \line_buffer.mem12_physical_MASK_wire\,
            WDATA => \line_buffer.mem12_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23169\,
            RE => \N__18196\,
            WCLKE => 'H',
            WCLK => \N__24606\,
            WE => \N__14393\
        );

    \line_buffer.mem24_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem24_physical_RDATA_wire\,
            RADDR => \line_buffer.mem24_physical_RADDR_wire\,
            WADDR => \line_buffer.mem24_physical_WADDR_wire\,
            MASK => \line_buffer.mem24_physical_MASK_wire\,
            WDATA => \line_buffer.mem24_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23542\,
            RE => \N__18208\,
            WCLKE => 'H',
            WCLK => \N__24589\,
            WE => \N__8613\
        );

    \line_buffer.mem1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem1_physical_RDATA_wire\,
            RADDR => \line_buffer.mem1_physical_RADDR_wire\,
            WADDR => \line_buffer.mem1_physical_WADDR_wire\,
            MASK => \line_buffer.mem1_physical_MASK_wire\,
            WDATA => \line_buffer.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23427\,
            RE => \N__18213\,
            WCLKE => 'H',
            WCLK => \N__24585\,
            WE => \N__13400\
        );

    \line_buffer.mem15_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem15_physical_RDATA_wire\,
            RADDR => \line_buffer.mem15_physical_RADDR_wire\,
            WADDR => \line_buffer.mem15_physical_WADDR_wire\,
            MASK => \line_buffer.mem15_physical_MASK_wire\,
            WDATA => \line_buffer.mem15_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23426\,
            RE => \N__18141\,
            WCLKE => 'H',
            WCLK => \N__24613\,
            WE => \N__13392\
        );

    \line_buffer.mem27_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem27_physical_RDATA_wire\,
            RADDR => \line_buffer.mem27_physical_RADDR_wire\,
            WADDR => \line_buffer.mem27_physical_WADDR_wire\,
            MASK => \line_buffer.mem27_physical_MASK_wire\,
            WDATA => \line_buffer.mem27_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23517\,
            RE => \N__18185\,
            WCLKE => 'H',
            WCLK => \N__24607\,
            WE => \N__9618\
        );

    \line_buffer.mem4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem4_physical_RDATA_wire\,
            RADDR => \line_buffer.mem4_physical_RADDR_wire\,
            WADDR => \line_buffer.mem4_physical_WADDR_wire\,
            MASK => \line_buffer.mem4_physical_MASK_wire\,
            WDATA => \line_buffer.mem4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23318\,
            RE => \N__18094\,
            WCLKE => 'H',
            WCLK => \N__24622\,
            WE => \N__8615\
        );

    \line_buffer.mem16_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem16_physical_RDATA_wire\,
            RADDR => \line_buffer.mem16_physical_RADDR_wire\,
            WADDR => \line_buffer.mem16_physical_WADDR_wire\,
            MASK => \line_buffer.mem16_physical_MASK_wire\,
            WDATA => \line_buffer.mem16_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23429\,
            RE => \N__18140\,
            WCLKE => 'H',
            WCLK => \N__24616\,
            WE => \N__13399\
        );

    \line_buffer.mem30_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem30_physical_RDATA_wire\,
            RADDR => \line_buffer.mem30_physical_RADDR_wire\,
            WADDR => \line_buffer.mem30_physical_WADDR_wire\,
            MASK => \line_buffer.mem30_physical_MASK_wire\,
            WDATA => \line_buffer.mem30_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23440\,
            RE => \N__18125\,
            WCLKE => 'H',
            WCLK => \N__24617\,
            WE => \N__13485\
        );

    \line_buffer.mem7_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem7_physical_RDATA_wire\,
            RADDR => \line_buffer.mem7_physical_RADDR_wire\,
            WADDR => \line_buffer.mem7_physical_WADDR_wire\,
            MASK => \line_buffer.mem7_physical_MASK_wire\,
            WDATA => \line_buffer.mem7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23011\,
            RE => \N__18052\,
            WCLKE => 'H',
            WCLK => \N__24630\,
            WE => \N__9375\
        );

    \line_buffer.mem20_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem20_physical_RDATA_wire\,
            RADDR => \line_buffer.mem20_physical_RADDR_wire\,
            WADDR => \line_buffer.mem20_physical_WADDR_wire\,
            MASK => \line_buffer.mem20_physical_MASK_wire\,
            WDATA => \line_buffer.mem20_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23091\,
            RE => \N__18088\,
            WCLKE => 'H',
            WCLK => \N__24629\,
            WE => \N__12690\
        );

    \line_buffer.mem13_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem13_physical_RDATA_wire\,
            RADDR => \line_buffer.mem13_physical_RADDR_wire\,
            WADDR => \line_buffer.mem13_physical_WADDR_wire\,
            MASK => \line_buffer.mem13_physical_MASK_wire\,
            WDATA => \line_buffer.mem13_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22997\,
            RE => \N__18171\,
            WCLKE => 'H',
            WCLK => \N__24608\,
            WE => \N__14394\
        );

    \line_buffer.mem19_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem19_physical_RDATA_wire\,
            RADDR => \line_buffer.mem19_physical_RADDR_wire\,
            WADDR => \line_buffer.mem19_physical_WADDR_wire\,
            MASK => \line_buffer.mem19_physical_MASK_wire\,
            WDATA => \line_buffer.mem19_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23124\,
            RE => \N__18073\,
            WCLKE => 'H',
            WCLK => \N__24623\,
            WE => \N__14182\
        );

    \line_buffer.mem23_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem23_physical_RDATA_wire\,
            RADDR => \line_buffer.mem23_physical_RADDR_wire\,
            WADDR => \line_buffer.mem23_physical_WADDR_wire\,
            MASK => \line_buffer.mem23_physical_MASK_wire\,
            WDATA => \line_buffer.mem23_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23546\,
            RE => \N__18217\,
            WCLKE => 'H',
            WCLK => \N__24579\,
            WE => \N__8614\
        );

    \line_buffer.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem0_physical_RDATA_wire\,
            RADDR => \line_buffer.mem0_physical_RADDR_wire\,
            WADDR => \line_buffer.mem0_physical_WADDR_wire\,
            MASK => \line_buffer.mem0_physical_MASK_wire\,
            WDATA => \line_buffer.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23428\,
            RE => \N__18218\,
            WCLKE => 'H',
            WCLK => \N__24574\,
            WE => \N__14399\
        );

    \line_buffer.mem26_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem26_physical_RDATA_wire\,
            RADDR => \line_buffer.mem26_physical_RADDR_wire\,
            WADDR => \line_buffer.mem26_physical_WADDR_wire\,
            MASK => \line_buffer.mem26_physical_MASK_wire\,
            WDATA => \line_buffer.mem26_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23526\,
            RE => \N__18186\,
            WCLKE => 'H',
            WCLK => \N__24603\,
            WE => \N__9640\
        );

    \line_buffer.mem3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem3_physical_RDATA_wire\,
            RADDR => \line_buffer.mem3_physical_RADDR_wire\,
            WADDR => \line_buffer.mem3_physical_WADDR_wire\,
            MASK => \line_buffer.mem3_physical_MASK_wire\,
            WDATA => \line_buffer.mem3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23304\,
            RE => \N__18126\,
            WCLKE => 'H',
            WCLK => \N__24615\,
            WE => \N__12680\
        );

    \line_buffer.mem17_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem17_physical_RDATA_wire\,
            RADDR => \line_buffer.mem17_physical_RADDR_wire\,
            WADDR => \line_buffer.mem17_physical_WADDR_wire\,
            MASK => \line_buffer.mem17_physical_MASK_wire\,
            WDATA => \line_buffer.mem17_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23312\,
            RE => \N__18110\,
            WCLKE => 'H',
            WCLK => \N__24618\,
            WE => \N__14174\
        );

    \line_buffer.mem31_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem31_physical_RDATA_wire\,
            RADDR => \line_buffer.mem31_physical_RADDR_wire\,
            WADDR => \line_buffer.mem31_physical_WADDR_wire\,
            MASK => \line_buffer.mem31_physical_MASK_wire\,
            WDATA => \line_buffer.mem31_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23165\,
            RE => \N__18095\,
            WCLKE => 'H',
            WCLK => \N__24620\,
            WE => \N__13486\
        );

    \line_buffer.mem9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem9_physical_RDATA_wire\,
            RADDR => \line_buffer.mem9_physical_RADDR_wire\,
            WADDR => \line_buffer.mem9_physical_WADDR_wire\,
            MASK => \line_buffer.mem9_physical_MASK_wire\,
            WDATA => \line_buffer.mem9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22644\,
            RE => \N__18093\,
            WCLKE => 'H',
            WCLK => \N__24637\,
            WE => \N__9383\
        );

    \line_buffer.mem29_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem29_physical_RDATA_wire\,
            RADDR => \line_buffer.mem29_physical_RADDR_wire\,
            WADDR => \line_buffer.mem29_physical_WADDR_wire\,
            MASK => \line_buffer.mem29_physical_MASK_wire\,
            WDATA => \line_buffer.mem29_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23456\,
            RE => \N__18155\,
            WCLKE => 'H',
            WCLK => \N__24612\,
            WE => \N__13484\
        );

    \line_buffer.mem6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem6_physical_RDATA_wire\,
            RADDR => \line_buffer.mem6_physical_RADDR_wire\,
            WADDR => \line_buffer.mem6_physical_WADDR_wire\,
            MASK => \line_buffer.mem6_physical_MASK_wire\,
            WDATA => \line_buffer.mem6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23182\,
            RE => \N__18050\,
            WCLKE => 'H',
            WCLK => \N__24627\,
            WE => \N__13493\
        );

    \line_buffer.mem10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem10_physical_RDATA_wire\,
            RADDR => \line_buffer.mem10_physical_RADDR_wire\,
            WADDR => \line_buffer.mem10_physical_WADDR_wire\,
            MASK => \line_buffer.mem10_physical_MASK_wire\,
            WDATA => \line_buffer.mem10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23321\,
            RE => \N__18212\,
            WCLKE => 'H',
            WCLK => \N__24593\,
            WE => \N__9361\
        );

    \line_buffer.mem22_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem22_physical_RDATA_wire\,
            RADDR => \line_buffer.mem22_physical_RADDR_wire\,
            WADDR => \line_buffer.mem22_physical_WADDR_wire\,
            MASK => \line_buffer.mem22_physical_MASK_wire\,
            WDATA => \line_buffer.mem22_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22751\,
            RE => \N__18124\,
            WCLKE => 'H',
            WCLK => \N__24636\,
            WE => \N__12695\
        );

    \line_buffer.mem25_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem25_physical_RDATA_wire\,
            RADDR => \line_buffer.mem25_physical_RADDR_wire\,
            WADDR => \line_buffer.mem25_physical_WADDR_wire\,
            MASK => \line_buffer.mem25_physical_MASK_wire\,
            WDATA => \line_buffer.mem25_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23535\,
            RE => \N__18207\,
            WCLKE => 'H',
            WCLK => \N__24598\,
            WE => \N__8603\
        );

    \line_buffer.mem8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem8_physical_RDATA_wire\,
            RADDR => \line_buffer.mem8_physical_RADDR_wire\,
            WADDR => \line_buffer.mem8_physical_WADDR_wire\,
            MASK => \line_buffer.mem8_physical_MASK_wire\,
            WDATA => \line_buffer.mem8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22844\,
            RE => \N__18053\,
            WCLKE => 'H',
            WCLK => \N__24632\,
            WE => \N__9382\
        );

    \line_buffer.mem28_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem28_physical_RDATA_wire\,
            RADDR => \line_buffer.mem28_physical_RADDR_wire\,
            WADDR => \line_buffer.mem28_physical_WADDR_wire\,
            MASK => \line_buffer.mem28_physical_MASK_wire\,
            WDATA => \line_buffer.mem28_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22833\,
            RE => \N__18156\,
            WCLKE => 'H',
            WCLK => \N__24610\,
            WE => \N__9636\
        );

    \line_buffer.mem18_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem18_physical_RDATA_wire\,
            RADDR => \line_buffer.mem18_physical_RADDR_wire\,
            WADDR => \line_buffer.mem18_physical_WADDR_wire\,
            MASK => \line_buffer.mem18_physical_MASK_wire\,
            WDATA => \line_buffer.mem18_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23328\,
            RE => \N__18109\,
            WCLKE => 'H',
            WCLK => \N__24621\,
            WE => \N__14175\
        );

    \DEBUG_c_2_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__25254\,
            GLOBALBUFFEROUTPUT => \DEBUG_c_2_c\
        );

    \DEBUG_c_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25256\,
            DIN => \N__25255\,
            DOUT => \N__25254\,
            PACKAGEPIN => \TVP_CLK_wire\
        );

    \DEBUG_c_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25256\,
            PADOUT => \N__25255\,
            PADIN => \N__25254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25245\,
            DIN => \N__25244\,
            DOUT => \N__25243\,
            PACKAGEPIN => \ADV_CLK_wire\
        );

    \ADV_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25245\,
            PADOUT => \N__25244\,
            PADIN => \N__25243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22910\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25236\,
            DIN => \N__25235\,
            DOUT => \N__25234\,
            PACKAGEPIN => DEBUG(3)
        );

    \DEBUG_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25236\,
            PADOUT => \N__25235\,
            PADIN => \N__25234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15601\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25227\,
            DIN => \N__25226\,
            DOUT => \N__25225\,
            PACKAGEPIN => \TVP_VIDEO_wire\(2)
        );

    \TVP_VIDEO_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25227\,
            PADOUT => \N__25226\,
            PADIN => \N__25225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25218\,
            DIN => \N__25217\,
            DOUT => \N__25216\,
            PACKAGEPIN => \ADV_G_wire\(5)
        );

    \ADV_G_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25218\,
            PADOUT => \N__25217\,
            PADIN => \N__25216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21310\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25209\,
            DIN => \N__25208\,
            DOUT => \N__25207\,
            PACKAGEPIN => \ADV_R_wire\(3)
        );

    \ADV_R_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25209\,
            PADOUT => \N__25208\,
            PADIN => \N__25207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23592\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25200\,
            DIN => \N__25199\,
            DOUT => \N__25198\,
            PACKAGEPIN => \TVP_VIDEO_wire\(5)
        );

    \DEBUG_c_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25200\,
            PADOUT => \N__25199\,
            PADIN => \N__25198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25191\,
            DIN => \N__25190\,
            DOUT => \N__25189\,
            PACKAGEPIN => \ADV_R_wire\(0)
        );

    \ADV_R_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25191\,
            PADOUT => \N__25190\,
            PADIN => \N__25189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21431\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25182\,
            DIN => \N__25181\,
            DOUT => \N__25180\,
            PACKAGEPIN => DEBUG(2)
        );

    \DEBUG_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25182\,
            PADOUT => \N__25181\,
            PADIN => \N__25180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8395\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25173\,
            DIN => \N__25172\,
            DOUT => \N__25171\,
            PACKAGEPIN => \TVP_VIDEO_wire\(3)
        );

    \TVP_VIDEO_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25173\,
            PADOUT => \N__25172\,
            PADIN => \N__25171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25164\,
            DIN => \N__25163\,
            DOUT => \N__25162\,
            PACKAGEPIN => \ADV_G_wire\(4)
        );

    \ADV_G_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25164\,
            PADOUT => \N__25163\,
            PADIN => \N__25162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24140\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25155\,
            DIN => \N__25154\,
            DOUT => \N__25153\,
            PACKAGEPIN => \ADV_R_wire\(5)
        );

    \ADV_R_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25155\,
            PADOUT => \N__25154\,
            PADIN => \N__25153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21317\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25146\,
            DIN => \N__25145\,
            DOUT => \N__25144\,
            PACKAGEPIN => DEBUG(1)
        );

    \DEBUG_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25146\,
            PADOUT => \N__25145\,
            PADIN => \N__25144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25137\,
            DIN => \N__25136\,
            DOUT => \N__25135\,
            PACKAGEPIN => \TVP_VIDEO_wire\(8)
        );

    \DEBUG_c_6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25137\,
            PADOUT => \N__25136\,
            PADIN => \N__25135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_6_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25128\,
            DIN => \N__25127\,
            DOUT => \N__25126\,
            PACKAGEPIN => \ADV_B_wire\(1)
        );

    \ADV_B_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25128\,
            PADOUT => \N__25127\,
            PADIN => \N__25126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21355\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_SYNC_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25119\,
            DIN => \N__25118\,
            DOUT => \N__25117\,
            PACKAGEPIN => \ADV_SYNC_N_wire\
        );

    \ADV_SYNC_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25119\,
            PADOUT => \N__25118\,
            PADIN => \N__25117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25110\,
            DIN => \N__25109\,
            DOUT => \N__25108\,
            PACKAGEPIN => \ADV_B_wire\(6)
        );

    \ADV_B_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25110\,
            PADOUT => \N__25109\,
            PADIN => \N__25108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21855\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25101\,
            DIN => \N__25100\,
            DOUT => \N__25099\,
            PACKAGEPIN => DEBUG(6)
        );

    \DEBUG_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25101\,
            PADOUT => \N__25100\,
            PADIN => \N__25099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18470\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25092\,
            DIN => \N__25091\,
            DOUT => \N__25090\,
            PACKAGEPIN => \ADV_G_wire\(0)
        );

    \ADV_G_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25092\,
            PADOUT => \N__25091\,
            PADIN => \N__25090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21423\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25083\,
            DIN => \N__25082\,
            DOUT => \N__25081\,
            PACKAGEPIN => \ADV_R_wire\(1)
        );

    \ADV_R_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25083\,
            PADOUT => \N__25082\,
            PADIN => \N__25081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21373\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25074\,
            DIN => \N__25073\,
            DOUT => \N__25072\,
            PACKAGEPIN => DEBUG(5)
        );

    \DEBUG_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25074\,
            PADOUT => \N__25073\,
            PADIN => \N__25072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16592\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25065\,
            DIN => \N__25064\,
            DOUT => \N__25063\,
            PACKAGEPIN => \ADV_G_wire\(7)
        );

    \ADV_G_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25065\,
            PADOUT => \N__25064\,
            PADIN => \N__25063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22207\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25056\,
            DIN => \N__25055\,
            DOUT => \N__25054\,
            PACKAGEPIN => \ADV_R_wire\(6)
        );

    \ADV_R_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25056\,
            PADOUT => \N__25055\,
            PADIN => \N__25054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21869\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_BLANK_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25047\,
            DIN => \N__25046\,
            DOUT => \N__25045\,
            PACKAGEPIN => \ADV_BLANK_N_wire\
        );

    \ADV_BLANK_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25047\,
            PADOUT => \N__25046\,
            PADIN => \N__25045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18071\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25038\,
            DIN => \N__25037\,
            DOUT => \N__25036\,
            PACKAGEPIN => DEBUG(0)
        );

    \DEBUG_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25038\,
            PADOUT => \N__25037\,
            PADIN => \N__25036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9479\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25029\,
            DIN => \N__25028\,
            DOUT => \N__25027\,
            PACKAGEPIN => \ADV_B_wire\(2)
        );

    \ADV_B_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25029\,
            PADOUT => \N__25028\,
            PADIN => \N__25027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25020\,
            DIN => \N__25019\,
            DOUT => \N__25018\,
            PACKAGEPIN => \TVP_VIDEO_wire\(9)
        );

    \DEBUG_c_7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25020\,
            PADOUT => \N__25019\,
            PADIN => \N__25018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_7_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25011\,
            DIN => \N__25010\,
            DOUT => \N__25009\,
            PACKAGEPIN => \TVP_HSYNC_wire\
        );

    \DEBUG_c_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25011\,
            PADOUT => \N__25010\,
            PADIN => \N__25009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25002\,
            DIN => \N__25001\,
            DOUT => \N__25000\,
            PACKAGEPIN => \TVP_VIDEO_wire\(7)
        );

    \DEBUG_c_5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25002\,
            PADOUT => \N__25001\,
            PADIN => \N__25000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_5_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24993\,
            DIN => \N__24992\,
            DOUT => \N__24991\,
            PACKAGEPIN => \ADV_B_wire\(7)
        );

    \ADV_B_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24993\,
            PADOUT => \N__24992\,
            PADIN => \N__24991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22197\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24984\,
            DIN => \N__24983\,
            DOUT => \N__24982\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24984\,
            PADOUT => \N__24983\,
            PADIN => \N__24982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8816\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24975\,
            DIN => \N__24974\,
            DOUT => \N__24973\,
            PACKAGEPIN => \TVP_VIDEO_wire\(4)
        );

    \TVP_VIDEO_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24975\,
            PADOUT => \N__24974\,
            PADIN => \N__24973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24966\,
            DIN => \N__24965\,
            DOUT => \N__24964\,
            PACKAGEPIN => \ADV_G_wire\(3)
        );

    \ADV_G_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24966\,
            PADOUT => \N__24965\,
            PADIN => \N__24964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23606\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24957\,
            DIN => \N__24956\,
            DOUT => \N__24955\,
            PACKAGEPIN => \ADV_HSYNC_wire\
        );

    \ADV_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24957\,
            PADOUT => \N__24956\,
            PADIN => \N__24955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16379\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24948\,
            DIN => \N__24947\,
            DOUT => \N__24946\,
            PACKAGEPIN => \ADV_R_wire\(2)
        );

    \ADV_R_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24948\,
            PADOUT => \N__24947\,
            PADIN => \N__24946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24939\,
            DIN => \N__24938\,
            DOUT => \N__24937\,
            PACKAGEPIN => \TVP_VSYNC_wire\
        );

    \DEBUG_c_0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24939\,
            PADOUT => \N__24938\,
            PADIN => \N__24937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_0_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24930\,
            DIN => \N__24929\,
            DOUT => \N__24928\,
            PACKAGEPIN => \ADV_B_wire\(4)
        );

    \ADV_B_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24930\,
            PADOUT => \N__24929\,
            PADIN => \N__24928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24136\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24921\,
            DIN => \N__24920\,
            DOUT => \N__24919\,
            PACKAGEPIN => DEBUG(4)
        );

    \DEBUG_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24921\,
            PADOUT => \N__24920\,
            PADIN => \N__24919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15575\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24912\,
            DIN => \N__24911\,
            DOUT => \N__24910\,
            PACKAGEPIN => \ADV_G_wire\(6)
        );

    \ADV_G_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24912\,
            PADOUT => \N__24911\,
            PADIN => \N__24910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21862\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24903\,
            DIN => \N__24902\,
            DOUT => \N__24901\,
            PACKAGEPIN => \ADV_R_wire\(7)
        );

    \ADV_R_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24903\,
            PADOUT => \N__24902\,
            PADIN => \N__24901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22208\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24894\,
            DIN => \N__24893\,
            DOUT => \N__24892\,
            PACKAGEPIN => \ADV_B_wire\(3)
        );

    \ADV_B_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24894\,
            PADOUT => \N__24893\,
            PADIN => \N__24892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23602\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24885\,
            DIN => \N__24884\,
            DOUT => \N__24883\,
            PACKAGEPIN => \ADV_R_wire\(4)
        );

    \ADV_R_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24885\,
            PADOUT => \N__24884\,
            PADIN => \N__24883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24126\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24876\,
            DIN => \N__24875\,
            DOUT => \N__24874\,
            PACKAGEPIN => \ADV_B_wire\(0)
        );

    \ADV_B_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24876\,
            PADOUT => \N__24875\,
            PADIN => \N__24874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21430\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24867\,
            DIN => \N__24866\,
            DOUT => \N__24865\,
            PACKAGEPIN => \ADV_G_wire\(2)
        );

    \ADV_G_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24867\,
            PADOUT => \N__24866\,
            PADIN => \N__24865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22268\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24858\,
            DIN => \N__24857\,
            DOUT => \N__24856\,
            PACKAGEPIN => \ADV_VSYNC_wire\
        );

    \ADV_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24858\,
            PADOUT => \N__24857\,
            PADIN => \N__24856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20420\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_4_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24849\,
            DIN => \N__24848\,
            DOUT => \N__24847\,
            PACKAGEPIN => \TVP_VIDEO_wire\(6)
        );

    \DEBUG_c_4_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24849\,
            PADOUT => \N__24848\,
            PADIN => \N__24847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_4_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24840\,
            DIN => \N__24839\,
            DOUT => \N__24838\,
            PACKAGEPIN => \ADV_B_wire\(5)
        );

    \ADV_B_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24840\,
            PADOUT => \N__24839\,
            PADIN => \N__24838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21303\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24831\,
            DIN => \N__24830\,
            DOUT => \N__24829\,
            PACKAGEPIN => DEBUG(7)
        );

    \DEBUG_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24831\,
            PADOUT => \N__24830\,
            PADIN => \N__24829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24683\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24822\,
            DIN => \N__24821\,
            DOUT => \N__24820\,
            PACKAGEPIN => \ADV_G_wire\(1)
        );

    \ADV_G_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24822\,
            PADOUT => \N__24821\,
            PADIN => \N__24820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21377\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__6017\ : SRMux
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__24800\,
            I => \N__24793\
        );

    \I__6015\ : SRMux
    port map (
            O => \N__24799\,
            I => \N__24789\
        );

    \I__6014\ : SRMux
    port map (
            O => \N__24798\,
            I => \N__24786\
        );

    \I__6013\ : SRMux
    port map (
            O => \N__24797\,
            I => \N__24781\
        );

    \I__6012\ : SRMux
    port map (
            O => \N__24796\,
            I => \N__24778\
        );

    \I__6011\ : Span4Mux_h
    port map (
            O => \N__24793\,
            I => \N__24775\
        );

    \I__6010\ : SRMux
    port map (
            O => \N__24792\,
            I => \N__24772\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__24789\,
            I => \N__24769\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__24786\,
            I => \N__24766\
        );

    \I__6007\ : SRMux
    port map (
            O => \N__24785\,
            I => \N__24763\
        );

    \I__6006\ : SRMux
    port map (
            O => \N__24784\,
            I => \N__24760\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__24781\,
            I => \N__24751\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__24778\,
            I => \N__24751\
        );

    \I__6003\ : Span4Mux_h
    port map (
            O => \N__24775\,
            I => \N__24751\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__24772\,
            I => \N__24751\
        );

    \I__6001\ : Span4Mux_v
    port map (
            O => \N__24769\,
            I => \N__24748\
        );

    \I__6000\ : Span4Mux_v
    port map (
            O => \N__24766\,
            I => \N__24741\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__24763\,
            I => \N__24741\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__24760\,
            I => \N__24741\
        );

    \I__5997\ : Span4Mux_v
    port map (
            O => \N__24751\,
            I => \N__24738\
        );

    \I__5996\ : Sp12to4
    port map (
            O => \N__24748\,
            I => \N__24733\
        );

    \I__5995\ : Sp12to4
    port map (
            O => \N__24741\,
            I => \N__24733\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__24738\,
            I => \transmit_module.n2367\
        );

    \I__5993\ : Odrv12
    port map (
            O => \N__24733\,
            I => \transmit_module.n2367\
        );

    \I__5992\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24725\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__24725\,
            I => \N__24722\
        );

    \I__5990\ : Odrv4
    port map (
            O => \N__24722\,
            I => \tvp_video_buffer.BUFFER_1_9\
        );

    \I__5989\ : InMux
    port map (
            O => \N__24719\,
            I => \N__24716\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__24716\,
            I => \N__24713\
        );

    \I__5987\ : Span12Mux_h
    port map (
            O => \N__24713\,
            I => \N__24710\
        );

    \I__5986\ : Span12Mux_v
    port map (
            O => \N__24710\,
            I => \N__24707\
        );

    \I__5985\ : Odrv12
    port map (
            O => \N__24707\,
            I => \line_buffer.n526\
        );

    \I__5984\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24701\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__24701\,
            I => \N__24698\
        );

    \I__5982\ : Span4Mux_h
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__5981\ : Span4Mux_v
    port map (
            O => \N__24695\,
            I => \N__24692\
        );

    \I__5980\ : Odrv4
    port map (
            O => \N__24692\,
            I => \line_buffer.n518\
        );

    \I__5979\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24686\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__24686\,
            I => \line_buffer.n3479\
        );

    \I__5977\ : IoInMux
    port map (
            O => \N__24683\,
            I => \N__24680\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24677\
        );

    \I__5975\ : IoSpan4Mux
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__5974\ : Span4Mux_s0_h
    port map (
            O => \N__24674\,
            I => \N__24671\
        );

    \I__5973\ : Sp12to4
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__5972\ : Span12Mux_s11_h
    port map (
            O => \N__24668\,
            I => \N__24665\
        );

    \I__5971\ : Span12Mux_v
    port map (
            O => \N__24665\,
            I => \N__24661\
        );

    \I__5970\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24658\
        );

    \I__5969\ : Span12Mux_h
    port map (
            O => \N__24661\,
            I => \N__24655\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__24658\,
            I => \N__24652\
        );

    \I__5967\ : Odrv12
    port map (
            O => \N__24655\,
            I => \DEBUG_c_7_c\
        );

    \I__5966\ : Odrv4
    port map (
            O => \N__24652\,
            I => \DEBUG_c_7_c\
        );

    \I__5965\ : InMux
    port map (
            O => \N__24647\,
            I => \N__24644\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__24644\,
            I => \tvp_video_buffer.BUFFER_0_9\
        );

    \I__5963\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__24638\,
            I => \N__24633\
        );

    \I__5961\ : ClkMux
    port map (
            O => \N__24637\,
            I => \N__24419\
        );

    \I__5960\ : ClkMux
    port map (
            O => \N__24636\,
            I => \N__24419\
        );

    \I__5959\ : Glb2LocalMux
    port map (
            O => \N__24633\,
            I => \N__24419\
        );

    \I__5958\ : ClkMux
    port map (
            O => \N__24632\,
            I => \N__24419\
        );

    \I__5957\ : ClkMux
    port map (
            O => \N__24631\,
            I => \N__24419\
        );

    \I__5956\ : ClkMux
    port map (
            O => \N__24630\,
            I => \N__24419\
        );

    \I__5955\ : ClkMux
    port map (
            O => \N__24629\,
            I => \N__24419\
        );

    \I__5954\ : ClkMux
    port map (
            O => \N__24628\,
            I => \N__24419\
        );

    \I__5953\ : ClkMux
    port map (
            O => \N__24627\,
            I => \N__24419\
        );

    \I__5952\ : ClkMux
    port map (
            O => \N__24626\,
            I => \N__24419\
        );

    \I__5951\ : ClkMux
    port map (
            O => \N__24625\,
            I => \N__24419\
        );

    \I__5950\ : ClkMux
    port map (
            O => \N__24624\,
            I => \N__24419\
        );

    \I__5949\ : ClkMux
    port map (
            O => \N__24623\,
            I => \N__24419\
        );

    \I__5948\ : ClkMux
    port map (
            O => \N__24622\,
            I => \N__24419\
        );

    \I__5947\ : ClkMux
    port map (
            O => \N__24621\,
            I => \N__24419\
        );

    \I__5946\ : ClkMux
    port map (
            O => \N__24620\,
            I => \N__24419\
        );

    \I__5945\ : ClkMux
    port map (
            O => \N__24619\,
            I => \N__24419\
        );

    \I__5944\ : ClkMux
    port map (
            O => \N__24618\,
            I => \N__24419\
        );

    \I__5943\ : ClkMux
    port map (
            O => \N__24617\,
            I => \N__24419\
        );

    \I__5942\ : ClkMux
    port map (
            O => \N__24616\,
            I => \N__24419\
        );

    \I__5941\ : ClkMux
    port map (
            O => \N__24615\,
            I => \N__24419\
        );

    \I__5940\ : ClkMux
    port map (
            O => \N__24614\,
            I => \N__24419\
        );

    \I__5939\ : ClkMux
    port map (
            O => \N__24613\,
            I => \N__24419\
        );

    \I__5938\ : ClkMux
    port map (
            O => \N__24612\,
            I => \N__24419\
        );

    \I__5937\ : ClkMux
    port map (
            O => \N__24611\,
            I => \N__24419\
        );

    \I__5936\ : ClkMux
    port map (
            O => \N__24610\,
            I => \N__24419\
        );

    \I__5935\ : ClkMux
    port map (
            O => \N__24609\,
            I => \N__24419\
        );

    \I__5934\ : ClkMux
    port map (
            O => \N__24608\,
            I => \N__24419\
        );

    \I__5933\ : ClkMux
    port map (
            O => \N__24607\,
            I => \N__24419\
        );

    \I__5932\ : ClkMux
    port map (
            O => \N__24606\,
            I => \N__24419\
        );

    \I__5931\ : ClkMux
    port map (
            O => \N__24605\,
            I => \N__24419\
        );

    \I__5930\ : ClkMux
    port map (
            O => \N__24604\,
            I => \N__24419\
        );

    \I__5929\ : ClkMux
    port map (
            O => \N__24603\,
            I => \N__24419\
        );

    \I__5928\ : ClkMux
    port map (
            O => \N__24602\,
            I => \N__24419\
        );

    \I__5927\ : ClkMux
    port map (
            O => \N__24601\,
            I => \N__24419\
        );

    \I__5926\ : ClkMux
    port map (
            O => \N__24600\,
            I => \N__24419\
        );

    \I__5925\ : ClkMux
    port map (
            O => \N__24599\,
            I => \N__24419\
        );

    \I__5924\ : ClkMux
    port map (
            O => \N__24598\,
            I => \N__24419\
        );

    \I__5923\ : ClkMux
    port map (
            O => \N__24597\,
            I => \N__24419\
        );

    \I__5922\ : ClkMux
    port map (
            O => \N__24596\,
            I => \N__24419\
        );

    \I__5921\ : ClkMux
    port map (
            O => \N__24595\,
            I => \N__24419\
        );

    \I__5920\ : ClkMux
    port map (
            O => \N__24594\,
            I => \N__24419\
        );

    \I__5919\ : ClkMux
    port map (
            O => \N__24593\,
            I => \N__24419\
        );

    \I__5918\ : ClkMux
    port map (
            O => \N__24592\,
            I => \N__24419\
        );

    \I__5917\ : ClkMux
    port map (
            O => \N__24591\,
            I => \N__24419\
        );

    \I__5916\ : ClkMux
    port map (
            O => \N__24590\,
            I => \N__24419\
        );

    \I__5915\ : ClkMux
    port map (
            O => \N__24589\,
            I => \N__24419\
        );

    \I__5914\ : ClkMux
    port map (
            O => \N__24588\,
            I => \N__24419\
        );

    \I__5913\ : ClkMux
    port map (
            O => \N__24587\,
            I => \N__24419\
        );

    \I__5912\ : ClkMux
    port map (
            O => \N__24586\,
            I => \N__24419\
        );

    \I__5911\ : ClkMux
    port map (
            O => \N__24585\,
            I => \N__24419\
        );

    \I__5910\ : ClkMux
    port map (
            O => \N__24584\,
            I => \N__24419\
        );

    \I__5909\ : ClkMux
    port map (
            O => \N__24583\,
            I => \N__24419\
        );

    \I__5908\ : ClkMux
    port map (
            O => \N__24582\,
            I => \N__24419\
        );

    \I__5907\ : ClkMux
    port map (
            O => \N__24581\,
            I => \N__24419\
        );

    \I__5906\ : ClkMux
    port map (
            O => \N__24580\,
            I => \N__24419\
        );

    \I__5905\ : ClkMux
    port map (
            O => \N__24579\,
            I => \N__24419\
        );

    \I__5904\ : ClkMux
    port map (
            O => \N__24578\,
            I => \N__24419\
        );

    \I__5903\ : ClkMux
    port map (
            O => \N__24577\,
            I => \N__24419\
        );

    \I__5902\ : ClkMux
    port map (
            O => \N__24576\,
            I => \N__24419\
        );

    \I__5901\ : ClkMux
    port map (
            O => \N__24575\,
            I => \N__24419\
        );

    \I__5900\ : ClkMux
    port map (
            O => \N__24574\,
            I => \N__24419\
        );

    \I__5899\ : ClkMux
    port map (
            O => \N__24573\,
            I => \N__24419\
        );

    \I__5898\ : ClkMux
    port map (
            O => \N__24572\,
            I => \N__24419\
        );

    \I__5897\ : ClkMux
    port map (
            O => \N__24571\,
            I => \N__24419\
        );

    \I__5896\ : ClkMux
    port map (
            O => \N__24570\,
            I => \N__24419\
        );

    \I__5895\ : ClkMux
    port map (
            O => \N__24569\,
            I => \N__24419\
        );

    \I__5894\ : ClkMux
    port map (
            O => \N__24568\,
            I => \N__24419\
        );

    \I__5893\ : ClkMux
    port map (
            O => \N__24567\,
            I => \N__24419\
        );

    \I__5892\ : ClkMux
    port map (
            O => \N__24566\,
            I => \N__24419\
        );

    \I__5891\ : ClkMux
    port map (
            O => \N__24565\,
            I => \N__24419\
        );

    \I__5890\ : ClkMux
    port map (
            O => \N__24564\,
            I => \N__24419\
        );

    \I__5889\ : GlobalMux
    port map (
            O => \N__24419\,
            I => \N__24416\
        );

    \I__5888\ : gio2CtrlBuf
    port map (
            O => \N__24416\,
            I => \DEBUG_c_2_c\
        );

    \I__5887\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24410\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__24410\,
            I => \N__24407\
        );

    \I__5885\ : Span4Mux_h
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__5884\ : Odrv4
    port map (
            O => \N__24404\,
            I => \line_buffer.n459\
        );

    \I__5883\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__5881\ : Sp12to4
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__5880\ : Span12Mux_v
    port map (
            O => \N__24392\,
            I => \N__24389\
        );

    \I__5879\ : Odrv12
    port map (
            O => \N__24389\,
            I => \line_buffer.n451\
        );

    \I__5878\ : InMux
    port map (
            O => \N__24386\,
            I => \N__24381\
        );

    \I__5877\ : InMux
    port map (
            O => \N__24385\,
            I => \N__24374\
        );

    \I__5876\ : InMux
    port map (
            O => \N__24384\,
            I => \N__24370\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__24381\,
            I => \N__24364\
        );

    \I__5874\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24359\
        );

    \I__5873\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24359\
        );

    \I__5872\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24354\
        );

    \I__5871\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24351\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24348\
        );

    \I__5869\ : InMux
    port map (
            O => \N__24373\,
            I => \N__24345\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__24370\,
            I => \N__24332\
        );

    \I__5867\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24329\
        );

    \I__5866\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24326\
        );

    \I__5865\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24323\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__24364\,
            I => \N__24320\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24317\
        );

    \I__5862\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24314\
        );

    \I__5861\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24311\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__24354\,
            I => \N__24307\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__24351\,
            I => \N__24304\
        );

    \I__5858\ : Span4Mux_v
    port map (
            O => \N__24348\,
            I => \N__24299\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__24345\,
            I => \N__24299\
        );

    \I__5856\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24296\
        );

    \I__5855\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24291\
        );

    \I__5854\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24291\
        );

    \I__5853\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24285\
        );

    \I__5852\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24285\
        );

    \I__5851\ : InMux
    port map (
            O => \N__24339\,
            I => \N__24282\
        );

    \I__5850\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24279\
        );

    \I__5849\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24276\
        );

    \I__5848\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24273\
        );

    \I__5847\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24270\
        );

    \I__5846\ : Span4Mux_v
    port map (
            O => \N__24332\,
            I => \N__24265\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24265\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__24326\,
            I => \N__24262\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__24323\,
            I => \N__24254\
        );

    \I__5842\ : Span4Mux_h
    port map (
            O => \N__24320\,
            I => \N__24254\
        );

    \I__5841\ : Span4Mux_v
    port map (
            O => \N__24317\,
            I => \N__24254\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24251\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__24311\,
            I => \N__24248\
        );

    \I__5838\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24245\
        );

    \I__5837\ : Span4Mux_h
    port map (
            O => \N__24307\,
            I => \N__24242\
        );

    \I__5836\ : Span4Mux_v
    port map (
            O => \N__24304\,
            I => \N__24233\
        );

    \I__5835\ : Span4Mux_v
    port map (
            O => \N__24299\,
            I => \N__24233\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__24296\,
            I => \N__24233\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__24291\,
            I => \N__24233\
        );

    \I__5832\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24230\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__24285\,
            I => \N__24227\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__24282\,
            I => \N__24224\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__24279\,
            I => \N__24217\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__24276\,
            I => \N__24217\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__24273\,
            I => \N__24217\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__24270\,
            I => \N__24210\
        );

    \I__5825\ : Span4Mux_v
    port map (
            O => \N__24265\,
            I => \N__24210\
        );

    \I__5824\ : Span4Mux_h
    port map (
            O => \N__24262\,
            I => \N__24210\
        );

    \I__5823\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24207\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__24254\,
            I => \N__24202\
        );

    \I__5821\ : Span4Mux_v
    port map (
            O => \N__24251\,
            I => \N__24202\
        );

    \I__5820\ : Span4Mux_h
    port map (
            O => \N__24248\,
            I => \N__24197\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__24245\,
            I => \N__24197\
        );

    \I__5818\ : Span4Mux_v
    port map (
            O => \N__24242\,
            I => \N__24194\
        );

    \I__5817\ : Sp12to4
    port map (
            O => \N__24233\,
            I => \N__24189\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24189\
        );

    \I__5815\ : Span4Mux_h
    port map (
            O => \N__24227\,
            I => \N__24184\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__24224\,
            I => \N__24184\
        );

    \I__5813\ : Span12Mux_h
    port map (
            O => \N__24217\,
            I => \N__24181\
        );

    \I__5812\ : Span4Mux_h
    port map (
            O => \N__24210\,
            I => \N__24178\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__24207\,
            I => \TX_ADDR_11\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__24202\,
            I => \TX_ADDR_11\
        );

    \I__5809\ : Odrv4
    port map (
            O => \N__24197\,
            I => \TX_ADDR_11\
        );

    \I__5808\ : Odrv4
    port map (
            O => \N__24194\,
            I => \TX_ADDR_11\
        );

    \I__5807\ : Odrv12
    port map (
            O => \N__24189\,
            I => \TX_ADDR_11\
        );

    \I__5806\ : Odrv4
    port map (
            O => \N__24184\,
            I => \TX_ADDR_11\
        );

    \I__5805\ : Odrv12
    port map (
            O => \N__24181\,
            I => \TX_ADDR_11\
        );

    \I__5804\ : Odrv4
    port map (
            O => \N__24178\,
            I => \TX_ADDR_11\
        );

    \I__5803\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24158\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__24158\,
            I => \N__24155\
        );

    \I__5801\ : Odrv12
    port map (
            O => \N__24155\,
            I => \line_buffer.n3518\
        );

    \I__5800\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24149\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__24149\,
            I => \N__24146\
        );

    \I__5798\ : Span4Mux_v
    port map (
            O => \N__24146\,
            I => \N__24143\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__24143\,
            I => \TX_DATA_4\
        );

    \I__5796\ : IoInMux
    port map (
            O => \N__24140\,
            I => \N__24137\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__24137\,
            I => \N__24133\
        );

    \I__5794\ : IoInMux
    port map (
            O => \N__24136\,
            I => \N__24130\
        );

    \I__5793\ : IoSpan4Mux
    port map (
            O => \N__24133\,
            I => \N__24127\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__24123\
        );

    \I__5791\ : Span4Mux_s2_v
    port map (
            O => \N__24127\,
            I => \N__24120\
        );

    \I__5790\ : IoInMux
    port map (
            O => \N__24126\,
            I => \N__24117\
        );

    \I__5789\ : IoSpan4Mux
    port map (
            O => \N__24123\,
            I => \N__24114\
        );

    \I__5788\ : Sp12to4
    port map (
            O => \N__24120\,
            I => \N__24111\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__24117\,
            I => \N__24108\
        );

    \I__5786\ : Span4Mux_s0_v
    port map (
            O => \N__24114\,
            I => \N__24105\
        );

    \I__5785\ : Span12Mux_s7_v
    port map (
            O => \N__24111\,
            I => \N__24100\
        );

    \I__5784\ : Span12Mux_s7_h
    port map (
            O => \N__24108\,
            I => \N__24100\
        );

    \I__5783\ : Span4Mux_v
    port map (
            O => \N__24105\,
            I => \N__24097\
        );

    \I__5782\ : Span12Mux_h
    port map (
            O => \N__24100\,
            I => \N__24094\
        );

    \I__5781\ : Span4Mux_v
    port map (
            O => \N__24097\,
            I => \N__24091\
        );

    \I__5780\ : Odrv12
    port map (
            O => \N__24094\,
            I => n1810
        );

    \I__5779\ : Odrv4
    port map (
            O => \N__24091\,
            I => n1810
        );

    \I__5778\ : InMux
    port map (
            O => \N__24086\,
            I => \N__24083\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__24083\,
            I => \N__24080\
        );

    \I__5776\ : Span12Mux_h
    port map (
            O => \N__24080\,
            I => \N__24077\
        );

    \I__5775\ : Span12Mux_v
    port map (
            O => \N__24077\,
            I => \N__24074\
        );

    \I__5774\ : Odrv12
    port map (
            O => \N__24074\,
            I => \line_buffer.n554\
        );

    \I__5773\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24068\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24065\
        );

    \I__5771\ : Span12Mux_h
    port map (
            O => \N__24065\,
            I => \N__24062\
        );

    \I__5770\ : Span12Mux_h
    port map (
            O => \N__24062\,
            I => \N__24059\
        );

    \I__5769\ : Odrv12
    port map (
            O => \N__24059\,
            I => \line_buffer.n562\
        );

    \I__5768\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24053\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__24053\,
            I => \line_buffer.n3585\
        );

    \I__5766\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24047\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__24047\,
            I => \N__24044\
        );

    \I__5764\ : Span4Mux_v
    port map (
            O => \N__24044\,
            I => \N__24041\
        );

    \I__5763\ : Span4Mux_v
    port map (
            O => \N__24041\,
            I => \N__24038\
        );

    \I__5762\ : Sp12to4
    port map (
            O => \N__24038\,
            I => \N__24035\
        );

    \I__5761\ : Odrv12
    port map (
            O => \N__24035\,
            I => \line_buffer.n558\
        );

    \I__5760\ : InMux
    port map (
            O => \N__24032\,
            I => \N__24029\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__24026\
        );

    \I__5758\ : Span4Mux_v
    port map (
            O => \N__24026\,
            I => \N__24023\
        );

    \I__5757\ : Span4Mux_h
    port map (
            O => \N__24023\,
            I => \N__24020\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__24020\,
            I => \line_buffer.n550\
        );

    \I__5755\ : CascadeMux
    port map (
            O => \N__24017\,
            I => \N__24012\
        );

    \I__5754\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24005\
        );

    \I__5753\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24002\
        );

    \I__5752\ : InMux
    port map (
            O => \N__24012\,
            I => \N__23999\
        );

    \I__5751\ : InMux
    port map (
            O => \N__24011\,
            I => \N__23993\
        );

    \I__5750\ : InMux
    port map (
            O => \N__24010\,
            I => \N__23990\
        );

    \I__5749\ : CascadeMux
    port map (
            O => \N__24009\,
            I => \N__23987\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__24008\,
            I => \N__23983\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__24005\,
            I => \N__23980\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23975\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__23999\,
            I => \N__23975\
        );

    \I__5744\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23971\
        );

    \I__5743\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23968\
        );

    \I__5742\ : InMux
    port map (
            O => \N__23996\,
            I => \N__23965\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__23993\,
            I => \N__23960\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__23990\,
            I => \N__23960\
        );

    \I__5739\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23957\
        );

    \I__5738\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23954\
        );

    \I__5737\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23951\
        );

    \I__5736\ : Span4Mux_v
    port map (
            O => \N__23980\,
            I => \N__23946\
        );

    \I__5735\ : Span4Mux_h
    port map (
            O => \N__23975\,
            I => \N__23943\
        );

    \I__5734\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23940\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__23971\,
            I => \N__23937\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__23968\,
            I => \N__23928\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__23965\,
            I => \N__23928\
        );

    \I__5730\ : Span4Mux_h
    port map (
            O => \N__23960\,
            I => \N__23928\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__23957\,
            I => \N__23928\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__23954\,
            I => \N__23923\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23923\
        );

    \I__5726\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23920\
        );

    \I__5725\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23917\
        );

    \I__5724\ : Span4Mux_h
    port map (
            O => \N__23946\,
            I => \N__23914\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__23943\,
            I => \N__23911\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__23940\,
            I => \N__23902\
        );

    \I__5721\ : Span4Mux_v
    port map (
            O => \N__23937\,
            I => \N__23902\
        );

    \I__5720\ : Span4Mux_v
    port map (
            O => \N__23928\,
            I => \N__23902\
        );

    \I__5719\ : Span4Mux_h
    port map (
            O => \N__23923\,
            I => \N__23902\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__23920\,
            I => \N__23899\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__23917\,
            I => \TX_ADDR_13\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__23914\,
            I => \TX_ADDR_13\
        );

    \I__5715\ : Odrv4
    port map (
            O => \N__23911\,
            I => \TX_ADDR_13\
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__23902\,
            I => \TX_ADDR_13\
        );

    \I__5713\ : Odrv4
    port map (
            O => \N__23899\,
            I => \TX_ADDR_13\
        );

    \I__5712\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__23885\,
            I => \N__23882\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__23882\,
            I => \line_buffer.n3482\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__23879\,
            I => \line_buffer.n3567_cascade_\
        );

    \I__5708\ : InMux
    port map (
            O => \N__23876\,
            I => \N__23873\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__23873\,
            I => \line_buffer.n3483\
        );

    \I__5706\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23867\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__23867\,
            I => \N__23864\
        );

    \I__5704\ : Span4Mux_v
    port map (
            O => \N__23864\,
            I => \N__23861\
        );

    \I__5703\ : Span4Mux_v
    port map (
            O => \N__23861\,
            I => \N__23858\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__23858\,
            I => \N__23855\
        );

    \I__5701\ : Sp12to4
    port map (
            O => \N__23855\,
            I => \N__23852\
        );

    \I__5700\ : Odrv12
    port map (
            O => \N__23852\,
            I => \line_buffer.n559\
        );

    \I__5699\ : CascadeMux
    port map (
            O => \N__23849\,
            I => \N__23837\
        );

    \I__5698\ : CascadeMux
    port map (
            O => \N__23848\,
            I => \N__23834\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__23847\,
            I => \N__23828\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__23846\,
            I => \N__23823\
        );

    \I__5695\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23820\
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__23844\,
            I => \N__23813\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__23843\,
            I => \N__23810\
        );

    \I__5692\ : CascadeMux
    port map (
            O => \N__23842\,
            I => \N__23807\
        );

    \I__5691\ : CascadeMux
    port map (
            O => \N__23841\,
            I => \N__23803\
        );

    \I__5690\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23798\
        );

    \I__5689\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23798\
        );

    \I__5688\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23795\
        );

    \I__5687\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23792\
        );

    \I__5686\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23789\
        );

    \I__5685\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23784\
        );

    \I__5684\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23784\
        );

    \I__5683\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23780\
        );

    \I__5682\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23777\
        );

    \I__5681\ : InMux
    port map (
            O => \N__23823\,
            I => \N__23774\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__23820\,
            I => \N__23771\
        );

    \I__5679\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23768\
        );

    \I__5678\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23759\
        );

    \I__5677\ : InMux
    port map (
            O => \N__23817\,
            I => \N__23759\
        );

    \I__5676\ : InMux
    port map (
            O => \N__23816\,
            I => \N__23759\
        );

    \I__5675\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23759\
        );

    \I__5674\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23756\
        );

    \I__5673\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23753\
        );

    \I__5672\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23750\
        );

    \I__5671\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23747\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23742\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__23795\,
            I => \N__23742\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__23792\,
            I => \N__23737\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__23789\,
            I => \N__23737\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23734\
        );

    \I__5665\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23730\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23723\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__23777\,
            I => \N__23723\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__23774\,
            I => \N__23723\
        );

    \I__5661\ : Span4Mux_v
    port map (
            O => \N__23771\,
            I => \N__23712\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__23768\,
            I => \N__23712\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__23759\,
            I => \N__23712\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__23756\,
            I => \N__23712\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__23753\,
            I => \N__23712\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__23750\,
            I => \N__23707\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__23747\,
            I => \N__23707\
        );

    \I__5654\ : Span4Mux_h
    port map (
            O => \N__23742\,
            I => \N__23704\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__23737\,
            I => \N__23699\
        );

    \I__5652\ : Span4Mux_h
    port map (
            O => \N__23734\,
            I => \N__23699\
        );

    \I__5651\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23696\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__23730\,
            I => \N__23693\
        );

    \I__5649\ : Span4Mux_v
    port map (
            O => \N__23723\,
            I => \N__23686\
        );

    \I__5648\ : Span4Mux_h
    port map (
            O => \N__23712\,
            I => \N__23686\
        );

    \I__5647\ : Span4Mux_v
    port map (
            O => \N__23707\,
            I => \N__23686\
        );

    \I__5646\ : Span4Mux_h
    port map (
            O => \N__23704\,
            I => \N__23683\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__23699\,
            I => \N__23680\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__23696\,
            I => \TX_ADDR_12\
        );

    \I__5643\ : Odrv4
    port map (
            O => \N__23693\,
            I => \TX_ADDR_12\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__23686\,
            I => \TX_ADDR_12\
        );

    \I__5641\ : Odrv4
    port map (
            O => \N__23683\,
            I => \TX_ADDR_12\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__23680\,
            I => \TX_ADDR_12\
        );

    \I__5639\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__5636\ : Odrv4
    port map (
            O => \N__23660\,
            I => \line_buffer.n551\
        );

    \I__5635\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23654\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__23654\,
            I => \line_buffer.n3543\
        );

    \I__5633\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23648\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__23648\,
            I => \N__23645\
        );

    \I__5631\ : Span12Mux_h
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__5630\ : Span12Mux_v
    port map (
            O => \N__23642\,
            I => \N__23639\
        );

    \I__5629\ : Odrv12
    port map (
            O => \N__23639\,
            I => \line_buffer.n582\
        );

    \I__5628\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__5626\ : Span12Mux_h
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__5625\ : Odrv12
    port map (
            O => \N__23627\,
            I => \line_buffer.n590\
        );

    \I__5624\ : InMux
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__23621\,
            I => \line_buffer.n3480\
        );

    \I__5622\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__23609\,
            I => \TX_DATA_3\
        );

    \I__5618\ : IoInMux
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23599\
        );

    \I__5616\ : IoInMux
    port map (
            O => \N__23602\,
            I => \N__23596\
        );

    \I__5615\ : IoSpan4Mux
    port map (
            O => \N__23599\,
            I => \N__23593\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__23596\,
            I => \N__23589\
        );

    \I__5613\ : Span4Mux_s3_v
    port map (
            O => \N__23593\,
            I => \N__23586\
        );

    \I__5612\ : IoInMux
    port map (
            O => \N__23592\,
            I => \N__23583\
        );

    \I__5611\ : Span4Mux_s3_v
    port map (
            O => \N__23589\,
            I => \N__23580\
        );

    \I__5610\ : Sp12to4
    port map (
            O => \N__23586\,
            I => \N__23577\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__23583\,
            I => \N__23574\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__23580\,
            I => \N__23571\
        );

    \I__5607\ : Span12Mux_s11_v
    port map (
            O => \N__23577\,
            I => \N__23568\
        );

    \I__5606\ : Span12Mux_s8_h
    port map (
            O => \N__23574\,
            I => \N__23565\
        );

    \I__5605\ : Span4Mux_v
    port map (
            O => \N__23571\,
            I => \N__23562\
        );

    \I__5604\ : Span12Mux_h
    port map (
            O => \N__23568\,
            I => \N__23559\
        );

    \I__5603\ : Span12Mux_h
    port map (
            O => \N__23565\,
            I => \N__23556\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__23562\,
            I => \N__23553\
        );

    \I__5601\ : Odrv12
    port map (
            O => \N__23559\,
            I => n1811
        );

    \I__5600\ : Odrv12
    port map (
            O => \N__23556\,
            I => n1811
        );

    \I__5599\ : Odrv4
    port map (
            O => \N__23553\,
            I => n1811
        );

    \I__5598\ : ClkMux
    port map (
            O => \N__23546\,
            I => \N__23543\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__23543\,
            I => \N__23539\
        );

    \I__5596\ : ClkMux
    port map (
            O => \N__23542\,
            I => \N__23536\
        );

    \I__5595\ : Span4Mux_h
    port map (
            O => \N__23539\,
            I => \N__23530\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__23536\,
            I => \N__23530\
        );

    \I__5593\ : ClkMux
    port map (
            O => \N__23535\,
            I => \N__23527\
        );

    \I__5592\ : Span4Mux_v
    port map (
            O => \N__23530\,
            I => \N__23521\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__23527\,
            I => \N__23521\
        );

    \I__5590\ : ClkMux
    port map (
            O => \N__23526\,
            I => \N__23518\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__23521\,
            I => \N__23511\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__23518\,
            I => \N__23511\
        );

    \I__5587\ : ClkMux
    port map (
            O => \N__23517\,
            I => \N__23508\
        );

    \I__5586\ : ClkMux
    port map (
            O => \N__23516\,
            I => \N__23502\
        );

    \I__5585\ : Span4Mux_v
    port map (
            O => \N__23511\,
            I => \N__23493\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__23508\,
            I => \N__23493\
        );

    \I__5583\ : ClkMux
    port map (
            O => \N__23507\,
            I => \N__23490\
        );

    \I__5582\ : ClkMux
    port map (
            O => \N__23506\,
            I => \N__23487\
        );

    \I__5581\ : ClkMux
    port map (
            O => \N__23505\,
            I => \N__23479\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__23502\,
            I => \N__23476\
        );

    \I__5579\ : ClkMux
    port map (
            O => \N__23501\,
            I => \N__23473\
        );

    \I__5578\ : ClkMux
    port map (
            O => \N__23500\,
            I => \N__23469\
        );

    \I__5577\ : ClkMux
    port map (
            O => \N__23499\,
            I => \N__23465\
        );

    \I__5576\ : ClkMux
    port map (
            O => \N__23498\,
            I => \N__23460\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__23493\,
            I => \N__23450\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__23490\,
            I => \N__23450\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__23487\,
            I => \N__23447\
        );

    \I__5572\ : ClkMux
    port map (
            O => \N__23486\,
            I => \N__23444\
        );

    \I__5571\ : ClkMux
    port map (
            O => \N__23485\,
            I => \N__23441\
        );

    \I__5570\ : ClkMux
    port map (
            O => \N__23484\,
            I => \N__23437\
        );

    \I__5569\ : ClkMux
    port map (
            O => \N__23483\,
            I => \N__23430\
        );

    \I__5568\ : ClkMux
    port map (
            O => \N__23482\,
            I => \N__23423\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23419\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__23476\,
            I => \N__23414\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__23473\,
            I => \N__23414\
        );

    \I__5564\ : ClkMux
    port map (
            O => \N__23472\,
            I => \N__23411\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__23469\,
            I => \N__23408\
        );

    \I__5562\ : ClkMux
    port map (
            O => \N__23468\,
            I => \N__23405\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__23465\,
            I => \N__23401\
        );

    \I__5560\ : ClkMux
    port map (
            O => \N__23464\,
            I => \N__23398\
        );

    \I__5559\ : ClkMux
    port map (
            O => \N__23463\,
            I => \N__23394\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23386\
        );

    \I__5557\ : ClkMux
    port map (
            O => \N__23459\,
            I => \N__23383\
        );

    \I__5556\ : ClkMux
    port map (
            O => \N__23458\,
            I => \N__23380\
        );

    \I__5555\ : ClkMux
    port map (
            O => \N__23457\,
            I => \N__23373\
        );

    \I__5554\ : ClkMux
    port map (
            O => \N__23456\,
            I => \N__23368\
        );

    \I__5553\ : ClkMux
    port map (
            O => \N__23455\,
            I => \N__23365\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__23450\,
            I => \N__23361\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__23447\,
            I => \N__23354\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23354\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__23441\,
            I => \N__23354\
        );

    \I__5548\ : ClkMux
    port map (
            O => \N__23440\,
            I => \N__23351\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__23437\,
            I => \N__23348\
        );

    \I__5546\ : ClkMux
    port map (
            O => \N__23436\,
            I => \N__23345\
        );

    \I__5545\ : ClkMux
    port map (
            O => \N__23435\,
            I => \N__23342\
        );

    \I__5544\ : ClkMux
    port map (
            O => \N__23434\,
            I => \N__23339\
        );

    \I__5543\ : ClkMux
    port map (
            O => \N__23433\,
            I => \N__23336\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__23430\,
            I => \N__23332\
        );

    \I__5541\ : ClkMux
    port map (
            O => \N__23429\,
            I => \N__23329\
        );

    \I__5540\ : ClkMux
    port map (
            O => \N__23428\,
            I => \N__23325\
        );

    \I__5539\ : ClkMux
    port map (
            O => \N__23427\,
            I => \N__23322\
        );

    \I__5538\ : ClkMux
    port map (
            O => \N__23426\,
            I => \N__23313\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__23423\,
            I => \N__23309\
        );

    \I__5536\ : ClkMux
    port map (
            O => \N__23422\,
            I => \N__23306\
        );

    \I__5535\ : Span4Mux_h
    port map (
            O => \N__23419\,
            I => \N__23295\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__23414\,
            I => \N__23295\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__23411\,
            I => \N__23295\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__23408\,
            I => \N__23290\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__23405\,
            I => \N__23290\
        );

    \I__5530\ : ClkMux
    port map (
            O => \N__23404\,
            I => \N__23287\
        );

    \I__5529\ : Span4Mux_h
    port map (
            O => \N__23401\,
            I => \N__23282\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__23398\,
            I => \N__23282\
        );

    \I__5527\ : ClkMux
    port map (
            O => \N__23397\,
            I => \N__23279\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23276\
        );

    \I__5525\ : ClkMux
    port map (
            O => \N__23393\,
            I => \N__23273\
        );

    \I__5524\ : ClkMux
    port map (
            O => \N__23392\,
            I => \N__23270\
        );

    \I__5523\ : ClkMux
    port map (
            O => \N__23391\,
            I => \N__23267\
        );

    \I__5522\ : ClkMux
    port map (
            O => \N__23390\,
            I => \N__23264\
        );

    \I__5521\ : ClkMux
    port map (
            O => \N__23389\,
            I => \N__23259\
        );

    \I__5520\ : Span4Mux_h
    port map (
            O => \N__23386\,
            I => \N__23254\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__23383\,
            I => \N__23254\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__23380\,
            I => \N__23251\
        );

    \I__5517\ : ClkMux
    port map (
            O => \N__23379\,
            I => \N__23248\
        );

    \I__5516\ : ClkMux
    port map (
            O => \N__23378\,
            I => \N__23245\
        );

    \I__5515\ : ClkMux
    port map (
            O => \N__23377\,
            I => \N__23242\
        );

    \I__5514\ : ClkMux
    port map (
            O => \N__23376\,
            I => \N__23239\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__23373\,
            I => \N__23236\
        );

    \I__5512\ : ClkMux
    port map (
            O => \N__23372\,
            I => \N__23233\
        );

    \I__5511\ : ClkMux
    port map (
            O => \N__23371\,
            I => \N__23230\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__23368\,
            I => \N__23222\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__23365\,
            I => \N__23222\
        );

    \I__5508\ : ClkMux
    port map (
            O => \N__23364\,
            I => \N__23219\
        );

    \I__5507\ : Span4Mux_v
    port map (
            O => \N__23361\,
            I => \N__23213\
        );

    \I__5506\ : Span4Mux_h
    port map (
            O => \N__23354\,
            I => \N__23213\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__23351\,
            I => \N__23206\
        );

    \I__5504\ : Span4Mux_v
    port map (
            O => \N__23348\,
            I => \N__23206\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23206\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23201\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23201\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__23336\,
            I => \N__23198\
        );

    \I__5499\ : ClkMux
    port map (
            O => \N__23335\,
            I => \N__23195\
        );

    \I__5498\ : Span4Mux_h
    port map (
            O => \N__23332\,
            I => \N__23191\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__23329\,
            I => \N__23188\
        );

    \I__5496\ : ClkMux
    port map (
            O => \N__23328\,
            I => \N__23185\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__23325\,
            I => \N__23179\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__23322\,
            I => \N__23176\
        );

    \I__5493\ : ClkMux
    port map (
            O => \N__23321\,
            I => \N__23173\
        );

    \I__5492\ : ClkMux
    port map (
            O => \N__23320\,
            I => \N__23170\
        );

    \I__5491\ : ClkMux
    port map (
            O => \N__23319\,
            I => \N__23166\
        );

    \I__5490\ : ClkMux
    port map (
            O => \N__23318\,
            I => \N__23162\
        );

    \I__5489\ : ClkMux
    port map (
            O => \N__23317\,
            I => \N__23158\
        );

    \I__5488\ : ClkMux
    port map (
            O => \N__23316\,
            I => \N__23155\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__23313\,
            I => \N__23151\
        );

    \I__5486\ : ClkMux
    port map (
            O => \N__23312\,
            I => \N__23148\
        );

    \I__5485\ : Span4Mux_h
    port map (
            O => \N__23309\,
            I => \N__23142\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__23306\,
            I => \N__23142\
        );

    \I__5483\ : ClkMux
    port map (
            O => \N__23305\,
            I => \N__23139\
        );

    \I__5482\ : ClkMux
    port map (
            O => \N__23304\,
            I => \N__23136\
        );

    \I__5481\ : ClkMux
    port map (
            O => \N__23303\,
            I => \N__23133\
        );

    \I__5480\ : ClkMux
    port map (
            O => \N__23302\,
            I => \N__23126\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__23295\,
            I => \N__23112\
        );

    \I__5478\ : Span4Mux_h
    port map (
            O => \N__23290\,
            I => \N__23112\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__23287\,
            I => \N__23112\
        );

    \I__5476\ : Span4Mux_h
    port map (
            O => \N__23282\,
            I => \N__23112\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23112\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__23276\,
            I => \N__23105\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__23273\,
            I => \N__23105\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__23270\,
            I => \N__23105\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__23267\,
            I => \N__23102\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__23264\,
            I => \N__23099\
        );

    \I__5469\ : ClkMux
    port map (
            O => \N__23263\,
            I => \N__23096\
        );

    \I__5468\ : ClkMux
    port map (
            O => \N__23262\,
            I => \N__23093\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__23259\,
            I => \N__23088\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__23254\,
            I => \N__23081\
        );

    \I__5465\ : Span4Mux_h
    port map (
            O => \N__23251\,
            I => \N__23081\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__23248\,
            I => \N__23081\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23078\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__23242\,
            I => \N__23075\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__23239\,
            I => \N__23072\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__23236\,
            I => \N__23065\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__23233\,
            I => \N__23065\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__23230\,
            I => \N__23065\
        );

    \I__5457\ : ClkMux
    port map (
            O => \N__23229\,
            I => \N__23062\
        );

    \I__5456\ : ClkMux
    port map (
            O => \N__23228\,
            I => \N__23058\
        );

    \I__5455\ : ClkMux
    port map (
            O => \N__23227\,
            I => \N__23054\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__23222\,
            I => \N__23049\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23049\
        );

    \I__5452\ : ClkMux
    port map (
            O => \N__23218\,
            I => \N__23046\
        );

    \I__5451\ : Span4Mux_v
    port map (
            O => \N__23213\,
            I => \N__23035\
        );

    \I__5450\ : Span4Mux_h
    port map (
            O => \N__23206\,
            I => \N__23035\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__23201\,
            I => \N__23035\
        );

    \I__5448\ : Span4Mux_h
    port map (
            O => \N__23198\,
            I => \N__23035\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__23195\,
            I => \N__23035\
        );

    \I__5446\ : ClkMux
    port map (
            O => \N__23194\,
            I => \N__23032\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__23191\,
            I => \N__23026\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__23188\,
            I => \N__23026\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23023\
        );

    \I__5442\ : ClkMux
    port map (
            O => \N__23184\,
            I => \N__23020\
        );

    \I__5441\ : ClkMux
    port map (
            O => \N__23183\,
            I => \N__23016\
        );

    \I__5440\ : ClkMux
    port map (
            O => \N__23182\,
            I => \N__23012\
        );

    \I__5439\ : Span4Mux_s2_v
    port map (
            O => \N__23179\,
            I => \N__23004\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__23176\,
            I => \N__23004\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__23173\,
            I => \N__23004\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__23170\,
            I => \N__23001\
        );

    \I__5435\ : ClkMux
    port map (
            O => \N__23169\,
            I => \N__22998\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__23166\,
            I => \N__22994\
        );

    \I__5433\ : ClkMux
    port map (
            O => \N__23165\,
            I => \N__22991\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__23162\,
            I => \N__22988\
        );

    \I__5431\ : ClkMux
    port map (
            O => \N__23161\,
            I => \N__22985\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__23158\,
            I => \N__22980\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__23155\,
            I => \N__22980\
        );

    \I__5428\ : ClkMux
    port map (
            O => \N__23154\,
            I => \N__22977\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__23151\,
            I => \N__22973\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__23148\,
            I => \N__22970\
        );

    \I__5425\ : ClkMux
    port map (
            O => \N__23147\,
            I => \N__22966\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__23142\,
            I => \N__22961\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__23139\,
            I => \N__22961\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__23136\,
            I => \N__22956\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__23133\,
            I => \N__22956\
        );

    \I__5420\ : ClkMux
    port map (
            O => \N__23132\,
            I => \N__22953\
        );

    \I__5419\ : ClkMux
    port map (
            O => \N__23131\,
            I => \N__22950\
        );

    \I__5418\ : ClkMux
    port map (
            O => \N__23130\,
            I => \N__22947\
        );

    \I__5417\ : ClkMux
    port map (
            O => \N__23129\,
            I => \N__22944\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__23126\,
            I => \N__22941\
        );

    \I__5415\ : ClkMux
    port map (
            O => \N__23125\,
            I => \N__22938\
        );

    \I__5414\ : ClkMux
    port map (
            O => \N__23124\,
            I => \N__22933\
        );

    \I__5413\ : ClkMux
    port map (
            O => \N__23123\,
            I => \N__22929\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__23112\,
            I => \N__22922\
        );

    \I__5411\ : Span4Mux_v
    port map (
            O => \N__23105\,
            I => \N__22922\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__23102\,
            I => \N__22922\
        );

    \I__5409\ : Span4Mux_v
    port map (
            O => \N__23099\,
            I => \N__22915\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__23096\,
            I => \N__22915\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__23093\,
            I => \N__22915\
        );

    \I__5406\ : ClkMux
    port map (
            O => \N__23092\,
            I => \N__22912\
        );

    \I__5405\ : ClkMux
    port map (
            O => \N__23091\,
            I => \N__22907\
        );

    \I__5404\ : Span4Mux_h
    port map (
            O => \N__23088\,
            I => \N__22900\
        );

    \I__5403\ : Span4Mux_h
    port map (
            O => \N__23081\,
            I => \N__22900\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__23078\,
            I => \N__22900\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__23075\,
            I => \N__22891\
        );

    \I__5400\ : Span4Mux_h
    port map (
            O => \N__23072\,
            I => \N__22891\
        );

    \I__5399\ : Span4Mux_h
    port map (
            O => \N__23065\,
            I => \N__22891\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__23062\,
            I => \N__22891\
        );

    \I__5397\ : ClkMux
    port map (
            O => \N__23061\,
            I => \N__22888\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__22885\
        );

    \I__5395\ : ClkMux
    port map (
            O => \N__23057\,
            I => \N__22882\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__23054\,
            I => \N__22879\
        );

    \I__5393\ : Span4Mux_h
    port map (
            O => \N__23049\,
            I => \N__22870\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__23046\,
            I => \N__22870\
        );

    \I__5391\ : Span4Mux_h
    port map (
            O => \N__23035\,
            I => \N__22870\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__23032\,
            I => \N__22870\
        );

    \I__5389\ : ClkMux
    port map (
            O => \N__23031\,
            I => \N__22867\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__23026\,
            I => \N__22860\
        );

    \I__5387\ : Span4Mux_h
    port map (
            O => \N__23023\,
            I => \N__22860\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__23020\,
            I => \N__22860\
        );

    \I__5385\ : ClkMux
    port map (
            O => \N__23019\,
            I => \N__22857\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__23016\,
            I => \N__22854\
        );

    \I__5383\ : ClkMux
    port map (
            O => \N__23015\,
            I => \N__22851\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__23012\,
            I => \N__22848\
        );

    \I__5381\ : ClkMux
    port map (
            O => \N__23011\,
            I => \N__22845\
        );

    \I__5380\ : Span4Mux_v
    port map (
            O => \N__23004\,
            I => \N__22837\
        );

    \I__5379\ : Span4Mux_h
    port map (
            O => \N__23001\,
            I => \N__22837\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__22998\,
            I => \N__22837\
        );

    \I__5377\ : ClkMux
    port map (
            O => \N__22997\,
            I => \N__22834\
        );

    \I__5376\ : Span4Mux_v
    port map (
            O => \N__22994\,
            I => \N__22824\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22824\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__22988\,
            I => \N__22824\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__22985\,
            I => \N__22824\
        );

    \I__5372\ : Span4Mux_v
    port map (
            O => \N__22980\,
            I => \N__22819\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__22977\,
            I => \N__22819\
        );

    \I__5370\ : ClkMux
    port map (
            O => \N__22976\,
            I => \N__22816\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__22973\,
            I => \N__22811\
        );

    \I__5368\ : Span4Mux_h
    port map (
            O => \N__22970\,
            I => \N__22811\
        );

    \I__5367\ : ClkMux
    port map (
            O => \N__22969\,
            I => \N__22808\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22805\
        );

    \I__5365\ : Span4Mux_v
    port map (
            O => \N__22961\,
            I => \N__22796\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__22956\,
            I => \N__22796\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__22953\,
            I => \N__22796\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22796\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22793\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__22944\,
            I => \N__22786\
        );

    \I__5359\ : Span4Mux_v
    port map (
            O => \N__22941\,
            I => \N__22786\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__22938\,
            I => \N__22786\
        );

    \I__5357\ : ClkMux
    port map (
            O => \N__22937\,
            I => \N__22783\
        );

    \I__5356\ : ClkMux
    port map (
            O => \N__22936\,
            I => \N__22780\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__22933\,
            I => \N__22776\
        );

    \I__5354\ : ClkMux
    port map (
            O => \N__22932\,
            I => \N__22773\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__22929\,
            I => \N__22769\
        );

    \I__5352\ : Span4Mux_v
    port map (
            O => \N__22922\,
            I => \N__22764\
        );

    \I__5351\ : Span4Mux_h
    port map (
            O => \N__22915\,
            I => \N__22764\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__22912\,
            I => \N__22761\
        );

    \I__5349\ : ClkMux
    port map (
            O => \N__22911\,
            I => \N__22758\
        );

    \I__5348\ : IoInMux
    port map (
            O => \N__22910\,
            I => \N__22755\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__22907\,
            I => \N__22752\
        );

    \I__5346\ : Span4Mux_v
    port map (
            O => \N__22900\,
            I => \N__22748\
        );

    \I__5345\ : Span4Mux_h
    port map (
            O => \N__22891\,
            I => \N__22745\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__22888\,
            I => \N__22742\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__22885\,
            I => \N__22739\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__22882\,
            I => \N__22736\
        );

    \I__5341\ : Span4Mux_v
    port map (
            O => \N__22879\,
            I => \N__22729\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__22870\,
            I => \N__22729\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__22867\,
            I => \N__22729\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__22860\,
            I => \N__22724\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N__22724\
        );

    \I__5336\ : Span4Mux_v
    port map (
            O => \N__22854\,
            I => \N__22719\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__22851\,
            I => \N__22719\
        );

    \I__5334\ : Span4Mux_h
    port map (
            O => \N__22848\,
            I => \N__22714\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__22845\,
            I => \N__22714\
        );

    \I__5332\ : ClkMux
    port map (
            O => \N__22844\,
            I => \N__22711\
        );

    \I__5331\ : Span4Mux_v
    port map (
            O => \N__22837\,
            I => \N__22707\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__22834\,
            I => \N__22704\
        );

    \I__5329\ : ClkMux
    port map (
            O => \N__22833\,
            I => \N__22701\
        );

    \I__5328\ : Span4Mux_h
    port map (
            O => \N__22824\,
            I => \N__22693\
        );

    \I__5327\ : Span4Mux_h
    port map (
            O => \N__22819\,
            I => \N__22693\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__22816\,
            I => \N__22693\
        );

    \I__5325\ : Span4Mux_h
    port map (
            O => \N__22811\,
            I => \N__22688\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__22808\,
            I => \N__22688\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__22805\,
            I => \N__22675\
        );

    \I__5322\ : Span4Mux_h
    port map (
            O => \N__22796\,
            I => \N__22675\
        );

    \I__5321\ : Span4Mux_v
    port map (
            O => \N__22793\,
            I => \N__22675\
        );

    \I__5320\ : Span4Mux_h
    port map (
            O => \N__22786\,
            I => \N__22675\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__22783\,
            I => \N__22675\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22675\
        );

    \I__5317\ : ClkMux
    port map (
            O => \N__22779\,
            I => \N__22672\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__22776\,
            I => \N__22669\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__22773\,
            I => \N__22666\
        );

    \I__5314\ : ClkMux
    port map (
            O => \N__22772\,
            I => \N__22663\
        );

    \I__5313\ : Span4Mux_v
    port map (
            O => \N__22769\,
            I => \N__22654\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__22764\,
            I => \N__22654\
        );

    \I__5311\ : Span4Mux_h
    port map (
            O => \N__22761\,
            I => \N__22654\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__22758\,
            I => \N__22654\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__22755\,
            I => \N__22651\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__22752\,
            I => \N__22648\
        );

    \I__5307\ : ClkMux
    port map (
            O => \N__22751\,
            I => \N__22645\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__22748\,
            I => \N__22637\
        );

    \I__5305\ : Span4Mux_v
    port map (
            O => \N__22745\,
            I => \N__22637\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__22742\,
            I => \N__22637\
        );

    \I__5303\ : Span4Mux_v
    port map (
            O => \N__22739\,
            I => \N__22632\
        );

    \I__5302\ : Span4Mux_h
    port map (
            O => \N__22736\,
            I => \N__22632\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__22729\,
            I => \N__22625\
        );

    \I__5300\ : Span4Mux_h
    port map (
            O => \N__22724\,
            I => \N__22625\
        );

    \I__5299\ : Span4Mux_h
    port map (
            O => \N__22719\,
            I => \N__22625\
        );

    \I__5298\ : Span4Mux_v
    port map (
            O => \N__22714\,
            I => \N__22620\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__22711\,
            I => \N__22620\
        );

    \I__5296\ : ClkMux
    port map (
            O => \N__22710\,
            I => \N__22617\
        );

    \I__5295\ : Sp12to4
    port map (
            O => \N__22707\,
            I => \N__22612\
        );

    \I__5294\ : Sp12to4
    port map (
            O => \N__22704\,
            I => \N__22612\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__22701\,
            I => \N__22609\
        );

    \I__5292\ : ClkMux
    port map (
            O => \N__22700\,
            I => \N__22606\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__22693\,
            I => \N__22597\
        );

    \I__5290\ : Span4Mux_h
    port map (
            O => \N__22688\,
            I => \N__22597\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__22675\,
            I => \N__22597\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__22672\,
            I => \N__22597\
        );

    \I__5287\ : Span4Mux_h
    port map (
            O => \N__22669\,
            I => \N__22590\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__22666\,
            I => \N__22590\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__22663\,
            I => \N__22590\
        );

    \I__5284\ : Span4Mux_h
    port map (
            O => \N__22654\,
            I => \N__22587\
        );

    \I__5283\ : Span4Mux_s1_v
    port map (
            O => \N__22651\,
            I => \N__22584\
        );

    \I__5282\ : Span4Mux_v
    port map (
            O => \N__22648\,
            I => \N__22579\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__22645\,
            I => \N__22579\
        );

    \I__5280\ : ClkMux
    port map (
            O => \N__22644\,
            I => \N__22576\
        );

    \I__5279\ : Span4Mux_v
    port map (
            O => \N__22637\,
            I => \N__22573\
        );

    \I__5278\ : Span4Mux_h
    port map (
            O => \N__22632\,
            I => \N__22570\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__22625\,
            I => \N__22567\
        );

    \I__5276\ : Span4Mux_h
    port map (
            O => \N__22620\,
            I => \N__22564\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__22617\,
            I => \N__22561\
        );

    \I__5274\ : Span12Mux_h
    port map (
            O => \N__22612\,
            I => \N__22554\
        );

    \I__5273\ : Span12Mux_h
    port map (
            O => \N__22609\,
            I => \N__22554\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__22606\,
            I => \N__22554\
        );

    \I__5271\ : Span4Mux_v
    port map (
            O => \N__22597\,
            I => \N__22549\
        );

    \I__5270\ : Span4Mux_h
    port map (
            O => \N__22590\,
            I => \N__22549\
        );

    \I__5269\ : Span4Mux_v
    port map (
            O => \N__22587\,
            I => \N__22546\
        );

    \I__5268\ : Sp12to4
    port map (
            O => \N__22584\,
            I => \N__22541\
        );

    \I__5267\ : Sp12to4
    port map (
            O => \N__22579\,
            I => \N__22541\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__22576\,
            I => \N__22538\
        );

    \I__5265\ : Span4Mux_v
    port map (
            O => \N__22573\,
            I => \N__22535\
        );

    \I__5264\ : Span4Mux_h
    port map (
            O => \N__22570\,
            I => \N__22528\
        );

    \I__5263\ : Span4Mux_v
    port map (
            O => \N__22567\,
            I => \N__22528\
        );

    \I__5262\ : Span4Mux_h
    port map (
            O => \N__22564\,
            I => \N__22528\
        );

    \I__5261\ : Span12Mux_h
    port map (
            O => \N__22561\,
            I => \N__22521\
        );

    \I__5260\ : Span12Mux_v
    port map (
            O => \N__22554\,
            I => \N__22521\
        );

    \I__5259\ : Sp12to4
    port map (
            O => \N__22549\,
            I => \N__22521\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__22546\,
            I => \N__22518\
        );

    \I__5257\ : Span12Mux_h
    port map (
            O => \N__22541\,
            I => \N__22513\
        );

    \I__5256\ : Span12Mux_h
    port map (
            O => \N__22538\,
            I => \N__22513\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__22535\,
            I => \ADV_CLK_c\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__22528\,
            I => \ADV_CLK_c\
        );

    \I__5253\ : Odrv12
    port map (
            O => \N__22521\,
            I => \ADV_CLK_c\
        );

    \I__5252\ : Odrv4
    port map (
            O => \N__22518\,
            I => \ADV_CLK_c\
        );

    \I__5251\ : Odrv12
    port map (
            O => \N__22513\,
            I => \ADV_CLK_c\
        );

    \I__5250\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__22496\,
            I => \N__22493\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__22493\,
            I => \N__22490\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__22490\,
            I => \line_buffer.n517\
        );

    \I__5245\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22484\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22481\
        );

    \I__5243\ : Span12Mux_v
    port map (
            O => \N__22481\,
            I => \N__22478\
        );

    \I__5242\ : Span12Mux_v
    port map (
            O => \N__22478\,
            I => \N__22475\
        );

    \I__5241\ : Odrv12
    port map (
            O => \N__22475\,
            I => \line_buffer.n525\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__22472\,
            I => \line_buffer.n3603_cascade_\
        );

    \I__5239\ : InMux
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__22466\,
            I => \line_buffer.n3606\
        );

    \I__5237\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__22460\,
            I => \N__22457\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__22457\,
            I => \N__22454\
        );

    \I__5234\ : Span4Mux_h
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__22451\,
            I => \line_buffer.n462\
        );

    \I__5232\ : CascadeMux
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__5231\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22442\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__5229\ : Span12Mux_h
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__5228\ : Span12Mux_v
    port map (
            O => \N__22436\,
            I => \N__22433\
        );

    \I__5227\ : Odrv12
    port map (
            O => \N__22433\,
            I => \line_buffer.n454\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__22430\,
            I => \line_buffer.n3546_cascade_\
        );

    \I__5225\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__22424\,
            I => \line_buffer.n3576\
        );

    \I__5223\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22418\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__5221\ : Span12Mux_v
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__5220\ : Odrv12
    port map (
            O => \N__22412\,
            I => \line_buffer.n555\
        );

    \I__5219\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__5217\ : Odrv12
    port map (
            O => \N__22403\,
            I => \line_buffer.n547\
        );

    \I__5216\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__5213\ : Span4Mux_h
    port map (
            O => \N__22391\,
            I => \N__22388\
        );

    \I__5212\ : Odrv4
    port map (
            O => \N__22388\,
            I => \line_buffer.n461\
        );

    \I__5211\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22379\
        );

    \I__5209\ : Span12Mux_h
    port map (
            O => \N__22379\,
            I => \N__22376\
        );

    \I__5208\ : Span12Mux_v
    port map (
            O => \N__22376\,
            I => \N__22373\
        );

    \I__5207\ : Odrv12
    port map (
            O => \N__22373\,
            I => \line_buffer.n453\
        );

    \I__5206\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__5204\ : Span12Mux_h
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__5203\ : Odrv12
    port map (
            O => \N__22361\,
            I => \line_buffer.n588\
        );

    \I__5202\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__5200\ : Span12Mux_h
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__5199\ : Span12Mux_v
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__5198\ : Odrv12
    port map (
            O => \N__22346\,
            I => \line_buffer.n580\
        );

    \I__5197\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__5195\ : Odrv4
    port map (
            O => \N__22337\,
            I => \line_buffer.n3522\
        );

    \I__5194\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22328\
        );

    \I__5192\ : Span4Mux_h
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__5191\ : Span4Mux_h
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__22322\,
            I => \line_buffer.n458\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__5188\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__5186\ : Span4Mux_v
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__5183\ : Span4Mux_v
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__22298\,
            I => \line_buffer.n450\
        );

    \I__5181\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__22289\,
            I => \line_buffer.n3579\
        );

    \I__5178\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__22283\,
            I => \line_buffer.n3582\
        );

    \I__5176\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__5174\ : Span4Mux_v
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__22271\,
            I => \TX_DATA_2\
        );

    \I__5172\ : IoInMux
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__22265\,
            I => \N__22262\
        );

    \I__5170\ : IoSpan4Mux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__5169\ : IoSpan4Mux
    port map (
            O => \N__22259\,
            I => \N__22255\
        );

    \I__5168\ : IoInMux
    port map (
            O => \N__22258\,
            I => \N__22252\
        );

    \I__5167\ : IoSpan4Mux
    port map (
            O => \N__22255\,
            I => \N__22247\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__22252\,
            I => \N__22247\
        );

    \I__5165\ : IoSpan4Mux
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__5164\ : Span4Mux_s0_h
    port map (
            O => \N__22244\,
            I => \N__22240\
        );

    \I__5163\ : IoInMux
    port map (
            O => \N__22243\,
            I => \N__22237\
        );

    \I__5162\ : Sp12to4
    port map (
            O => \N__22240\,
            I => \N__22234\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22231\
        );

    \I__5160\ : Span12Mux_s11_h
    port map (
            O => \N__22234\,
            I => \N__22228\
        );

    \I__5159\ : Span12Mux_s11_v
    port map (
            O => \N__22231\,
            I => \N__22225\
        );

    \I__5158\ : Odrv12
    port map (
            O => \N__22228\,
            I => n1812
        );

    \I__5157\ : Odrv12
    port map (
            O => \N__22225\,
            I => n1812
        );

    \I__5156\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__5154\ : Span4Mux_v
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__22211\,
            I => \TX_DATA_7\
        );

    \I__5152\ : IoInMux
    port map (
            O => \N__22208\,
            I => \N__22204\
        );

    \I__5151\ : IoInMux
    port map (
            O => \N__22207\,
            I => \N__22201\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__22204\,
            I => \N__22198\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__22201\,
            I => \N__22194\
        );

    \I__5148\ : IoSpan4Mux
    port map (
            O => \N__22198\,
            I => \N__22191\
        );

    \I__5147\ : IoInMux
    port map (
            O => \N__22197\,
            I => \N__22188\
        );

    \I__5146\ : Span4Mux_s3_v
    port map (
            O => \N__22194\,
            I => \N__22185\
        );

    \I__5145\ : Sp12to4
    port map (
            O => \N__22191\,
            I => \N__22182\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__22188\,
            I => \N__22179\
        );

    \I__5143\ : Span4Mux_h
    port map (
            O => \N__22185\,
            I => \N__22176\
        );

    \I__5142\ : Span12Mux_s6_h
    port map (
            O => \N__22182\,
            I => \N__22173\
        );

    \I__5141\ : Span12Mux_s4_v
    port map (
            O => \N__22179\,
            I => \N__22170\
        );

    \I__5140\ : Span4Mux_h
    port map (
            O => \N__22176\,
            I => \N__22167\
        );

    \I__5139\ : Span12Mux_h
    port map (
            O => \N__22173\,
            I => \N__22162\
        );

    \I__5138\ : Span12Mux_h
    port map (
            O => \N__22170\,
            I => \N__22162\
        );

    \I__5137\ : Span4Mux_v
    port map (
            O => \N__22167\,
            I => \N__22159\
        );

    \I__5136\ : Odrv12
    port map (
            O => \N__22162\,
            I => \ADV_B_c\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__22159\,
            I => \ADV_B_c\
        );

    \I__5134\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22151\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__22151\,
            I => \N__22145\
        );

    \I__5132\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22142\
        );

    \I__5131\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22139\
        );

    \I__5130\ : InMux
    port map (
            O => \N__22148\,
            I => \N__22136\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__22145\,
            I => \N__22129\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__22142\,
            I => \N__22122\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__22139\,
            I => \N__22122\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__22136\,
            I => \N__22122\
        );

    \I__5125\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22119\
        );

    \I__5124\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22116\
        );

    \I__5123\ : InMux
    port map (
            O => \N__22133\,
            I => \N__22113\
        );

    \I__5122\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22110\
        );

    \I__5121\ : Sp12to4
    port map (
            O => \N__22129\,
            I => \N__22107\
        );

    \I__5120\ : Span12Mux_s11_v
    port map (
            O => \N__22122\,
            I => \N__22100\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__22119\,
            I => \N__22100\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__22116\,
            I => \N__22100\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__22113\,
            I => \N__22095\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__22110\,
            I => \N__22095\
        );

    \I__5115\ : Span12Mux_h
    port map (
            O => \N__22107\,
            I => \N__22092\
        );

    \I__5114\ : Span12Mux_v
    port map (
            O => \N__22100\,
            I => \N__22089\
        );

    \I__5113\ : Span4Mux_s2_v
    port map (
            O => \N__22095\,
            I => \N__22086\
        );

    \I__5112\ : Span12Mux_v
    port map (
            O => \N__22092\,
            I => \N__22081\
        );

    \I__5111\ : Span12Mux_h
    port map (
            O => \N__22089\,
            I => \N__22081\
        );

    \I__5110\ : Span4Mux_h
    port map (
            O => \N__22086\,
            I => \N__22078\
        );

    \I__5109\ : Odrv12
    port map (
            O => \N__22081\,
            I => \RX_DATA_7\
        );

    \I__5108\ : Odrv4
    port map (
            O => \N__22078\,
            I => \RX_DATA_7\
        );

    \I__5107\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__5105\ : Span4Mux_v
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__5104\ : Span4Mux_v
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__5103\ : Span4Mux_h
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__22058\,
            I => \line_buffer.n465\
        );

    \I__5101\ : CascadeMux
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__5100\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__5098\ : Sp12to4
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__5097\ : Span12Mux_v
    port map (
            O => \N__22043\,
            I => \N__22040\
        );

    \I__5096\ : Odrv12
    port map (
            O => \N__22040\,
            I => \line_buffer.n457\
        );

    \I__5095\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22034\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__22034\,
            I => \line_buffer.n3588\
        );

    \I__5093\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22028\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__5091\ : Span12Mux_v
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__5090\ : Odrv12
    port map (
            O => \N__22022\,
            I => \line_buffer.n557\
        );

    \I__5089\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22016\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__22016\,
            I => \N__22013\
        );

    \I__5087\ : Span4Mux_h
    port map (
            O => \N__22013\,
            I => \N__22010\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__22007\,
            I => \line_buffer.n549\
        );

    \I__5084\ : InMux
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__5082\ : Span4Mux_v
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__21992\,
            I => \line_buffer.n460\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__5078\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21983\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__5075\ : Span4Mux_v
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__5074\ : Sp12to4
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__5073\ : Span12Mux_h
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__5072\ : Odrv12
    port map (
            O => \N__21968\,
            I => \line_buffer.n452\
        );

    \I__5071\ : InMux
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__5069\ : Odrv4
    port map (
            O => \N__21959\,
            I => \line_buffer.n3549\
        );

    \I__5068\ : CascadeMux
    port map (
            O => \N__21956\,
            I => \line_buffer.n3552_cascade_\
        );

    \I__5067\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__5065\ : Span12Mux_v
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__5064\ : Span12Mux_h
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__5063\ : Odrv12
    port map (
            O => \N__21941\,
            I => \line_buffer.n527\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__5061\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21932\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__5059\ : Span4Mux_v
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__5058\ : Span4Mux_h
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__5057\ : Span4Mux_v
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__5056\ : Odrv4
    port map (
            O => \N__21920\,
            I => \line_buffer.n519\
        );

    \I__5055\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21914\,
            I => \line_buffer.n3573\
        );

    \I__5053\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21908\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__5051\ : Span4Mux_v
    port map (
            O => \N__21905\,
            I => \N__21902\
        );

    \I__5050\ : Sp12to4
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__5049\ : Odrv12
    port map (
            O => \N__21899\,
            I => \line_buffer.n589\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__5046\ : Span4Mux_v
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__5045\ : Span4Mux_h
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__5044\ : Sp12to4
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__5043\ : Odrv12
    port map (
            O => \N__21881\,
            I => \line_buffer.n581\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__21872\,
            I => \TX_DATA_6\
        );

    \I__5039\ : IoInMux
    port map (
            O => \N__21869\,
            I => \N__21866\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__5037\ : Span4Mux_s1_h
    port map (
            O => \N__21863\,
            I => \N__21859\
        );

    \I__5036\ : IoInMux
    port map (
            O => \N__21862\,
            I => \N__21856\
        );

    \I__5035\ : Span4Mux_h
    port map (
            O => \N__21859\,
            I => \N__21852\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__21856\,
            I => \N__21849\
        );

    \I__5033\ : IoInMux
    port map (
            O => \N__21855\,
            I => \N__21846\
        );

    \I__5032\ : Span4Mux_h
    port map (
            O => \N__21852\,
            I => \N__21843\
        );

    \I__5031\ : IoSpan4Mux
    port map (
            O => \N__21849\,
            I => \N__21840\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__21846\,
            I => \N__21837\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__21843\,
            I => \N__21832\
        );

    \I__5028\ : Span4Mux_s2_v
    port map (
            O => \N__21840\,
            I => \N__21832\
        );

    \I__5027\ : Span12Mux_s11_v
    port map (
            O => \N__21837\,
            I => \N__21829\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__21832\,
            I => \N__21826\
        );

    \I__5025\ : Span12Mux_h
    port map (
            O => \N__21829\,
            I => \N__21823\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__21826\,
            I => \N__21820\
        );

    \I__5023\ : Odrv12
    port map (
            O => \N__21823\,
            I => n1808
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__21820\,
            I => n1808
        );

    \I__5021\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__5019\ : Sp12to4
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__5018\ : Span12Mux_v
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__5017\ : Odrv12
    port map (
            O => \N__21803\,
            I => \line_buffer.n528\
        );

    \I__5016\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__5014\ : Span4Mux_h
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__21788\,
            I => \line_buffer.n520\
        );

    \I__5011\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__5009\ : Odrv12
    port map (
            O => \N__21779\,
            I => \line_buffer.n3594\
        );

    \I__5008\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__5005\ : Sp12to4
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__5004\ : Odrv12
    port map (
            O => \N__21764\,
            I => \line_buffer.n592\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__5001\ : Span4Mux_v
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__5000\ : Span4Mux_v
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__21749\,
            I => \N__21746\
        );

    \I__4998\ : Span4Mux_h
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__21743\,
            I => \line_buffer.n584\
        );

    \I__4996\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__21737\,
            I => \line_buffer.n3489\
        );

    \I__4994\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__4992\ : Odrv12
    port map (
            O => \N__21728\,
            I => \line_buffer.n3488\
        );

    \I__4991\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__21722\,
            I => \line_buffer.n3561\
        );

    \I__4989\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__4987\ : Span4Mux_v
    port map (
            O => \N__21713\,
            I => \N__21710\
        );

    \I__4986\ : Sp12to4
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__4985\ : Odrv12
    port map (
            O => \N__21707\,
            I => \line_buffer.n591\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__4982\ : Span4Mux_v
    port map (
            O => \N__21698\,
            I => \N__21695\
        );

    \I__4981\ : Span4Mux_v
    port map (
            O => \N__21695\,
            I => \N__21692\
        );

    \I__4980\ : Span4Mux_v
    port map (
            O => \N__21692\,
            I => \N__21689\
        );

    \I__4979\ : Span4Mux_h
    port map (
            O => \N__21689\,
            I => \N__21686\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__21686\,
            I => \line_buffer.n583\
        );

    \I__4977\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21680\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__4975\ : Span4Mux_h
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__4973\ : Span4Mux_h
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__4972\ : Sp12to4
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__4971\ : Span12Mux_v
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__4970\ : Odrv12
    port map (
            O => \N__21662\,
            I => \line_buffer.n523\
        );

    \I__4969\ : CascadeMux
    port map (
            O => \N__21659\,
            I => \N__21656\
        );

    \I__4968\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__4966\ : Span4Mux_h
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__4965\ : Span4Mux_v
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__4964\ : Span4Mux_v
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__21641\,
            I => \line_buffer.n515\
        );

    \I__4962\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__21635\,
            I => \line_buffer.n3597\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__21632\,
            I => \line_buffer.n3600_cascade_\
        );

    \I__4959\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21626\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__21626\,
            I => \TX_DATA_0\
        );

    \I__4957\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21619\
        );

    \I__4956\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21615\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__21619\,
            I => \N__21608\
        );

    \I__4954\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21599\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__21615\,
            I => \N__21596\
        );

    \I__4952\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21593\
        );

    \I__4951\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21586\
        );

    \I__4950\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21586\
        );

    \I__4949\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21586\
        );

    \I__4948\ : Span4Mux_v
    port map (
            O => \N__21608\,
            I => \N__21582\
        );

    \I__4947\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21579\
        );

    \I__4946\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21572\
        );

    \I__4945\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21572\
        );

    \I__4944\ : InMux
    port map (
            O => \N__21604\,
            I => \N__21572\
        );

    \I__4943\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21569\
        );

    \I__4942\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21566\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21563\
        );

    \I__4940\ : Span4Mux_h
    port map (
            O => \N__21596\,
            I => \N__21558\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__21593\,
            I => \N__21558\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__21586\,
            I => \N__21555\
        );

    \I__4937\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21552\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__21582\,
            I => \N__21543\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__21579\,
            I => \N__21543\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__21572\,
            I => \N__21543\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21543\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__21566\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__4931\ : Odrv12
    port map (
            O => \N__21563\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__21558\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__21555\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__21552\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__4927\ : Odrv4
    port map (
            O => \N__21543\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__4926\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__4924\ : Odrv12
    port map (
            O => \N__21524\,
            I => \line_buffer.n3525\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__21521\,
            I => \line_buffer.n3524_cascade_\
        );

    \I__4922\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21515\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__21515\,
            I => \N__21512\
        );

    \I__4920\ : Odrv12
    port map (
            O => \N__21512\,
            I => \line_buffer.n3521\
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__21509\,
            I => \line_buffer.n3555_cascade_\
        );

    \I__4918\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21503\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__21503\,
            I => \line_buffer.n3519\
        );

    \I__4916\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__21497\,
            I => \N__21494\
        );

    \I__4914\ : Span4Mux_h
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__4913\ : Span4Mux_h
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__4912\ : Span4Mux_h
    port map (
            O => \N__21488\,
            I => \N__21485\
        );

    \I__4911\ : Odrv4
    port map (
            O => \N__21485\,
            I => \line_buffer.n561\
        );

    \I__4910\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__4908\ : Span4Mux_h
    port map (
            O => \N__21476\,
            I => \N__21473\
        );

    \I__4907\ : Span4Mux_h
    port map (
            O => \N__21473\,
            I => \N__21470\
        );

    \I__4906\ : Sp12to4
    port map (
            O => \N__21470\,
            I => \N__21467\
        );

    \I__4905\ : Span12Mux_v
    port map (
            O => \N__21467\,
            I => \N__21464\
        );

    \I__4904\ : Odrv12
    port map (
            O => \N__21464\,
            I => \line_buffer.n553\
        );

    \I__4903\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21458\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__21458\,
            I => \line_buffer.n3498\
        );

    \I__4901\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21452\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__21452\,
            I => \N__21449\
        );

    \I__4899\ : Odrv12
    port map (
            O => \N__21449\,
            I => \line_buffer.n587\
        );

    \I__4898\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21443\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__21443\,
            I => \N__21440\
        );

    \I__4896\ : Span12Mux_h
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__4895\ : Span12Mux_v
    port map (
            O => \N__21437\,
            I => \N__21434\
        );

    \I__4894\ : Odrv12
    port map (
            O => \N__21434\,
            I => \line_buffer.n579\
        );

    \I__4893\ : IoInMux
    port map (
            O => \N__21431\,
            I => \N__21427\
        );

    \I__4892\ : IoInMux
    port map (
            O => \N__21430\,
            I => \N__21424\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21420\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21417\
        );

    \I__4889\ : IoInMux
    port map (
            O => \N__21423\,
            I => \N__21414\
        );

    \I__4888\ : Span4Mux_s1_h
    port map (
            O => \N__21420\,
            I => \N__21411\
        );

    \I__4887\ : IoSpan4Mux
    port map (
            O => \N__21417\,
            I => \N__21408\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__21414\,
            I => \N__21403\
        );

    \I__4885\ : Sp12to4
    port map (
            O => \N__21411\,
            I => \N__21403\
        );

    \I__4884\ : Span4Mux_s3_v
    port map (
            O => \N__21408\,
            I => \N__21400\
        );

    \I__4883\ : Span12Mux_s11_v
    port map (
            O => \N__21403\,
            I => \N__21397\
        );

    \I__4882\ : Sp12to4
    port map (
            O => \N__21400\,
            I => \N__21394\
        );

    \I__4881\ : Span12Mux_h
    port map (
            O => \N__21397\,
            I => \N__21389\
        );

    \I__4880\ : Span12Mux_s11_v
    port map (
            O => \N__21394\,
            I => \N__21389\
        );

    \I__4879\ : Odrv12
    port map (
            O => \N__21389\,
            I => n1814
        );

    \I__4878\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21383\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__21380\,
            I => \TX_DATA_1\
        );

    \I__4875\ : IoInMux
    port map (
            O => \N__21377\,
            I => \N__21374\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__21374\,
            I => \N__21370\
        );

    \I__4873\ : IoInMux
    port map (
            O => \N__21373\,
            I => \N__21367\
        );

    \I__4872\ : Span4Mux_s1_v
    port map (
            O => \N__21370\,
            I => \N__21364\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__21367\,
            I => \N__21361\
        );

    \I__4870\ : Span4Mux_v
    port map (
            O => \N__21364\,
            I => \N__21356\
        );

    \I__4869\ : Span4Mux_s2_h
    port map (
            O => \N__21361\,
            I => \N__21356\
        );

    \I__4868\ : Span4Mux_h
    port map (
            O => \N__21356\,
            I => \N__21352\
        );

    \I__4867\ : IoInMux
    port map (
            O => \N__21355\,
            I => \N__21349\
        );

    \I__4866\ : Span4Mux_h
    port map (
            O => \N__21352\,
            I => \N__21346\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__21349\,
            I => \N__21343\
        );

    \I__4864\ : Sp12to4
    port map (
            O => \N__21346\,
            I => \N__21340\
        );

    \I__4863\ : Span4Mux_s3_v
    port map (
            O => \N__21343\,
            I => \N__21337\
        );

    \I__4862\ : Span12Mux_s10_v
    port map (
            O => \N__21340\,
            I => \N__21334\
        );

    \I__4861\ : Span4Mux_v
    port map (
            O => \N__21337\,
            I => \N__21331\
        );

    \I__4860\ : Odrv12
    port map (
            O => \N__21334\,
            I => n1813
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__21331\,
            I => n1813
        );

    \I__4858\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21323\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__21323\,
            I => \N__21320\
        );

    \I__4856\ : Odrv12
    port map (
            O => \N__21320\,
            I => \TX_DATA_5\
        );

    \I__4855\ : IoInMux
    port map (
            O => \N__21317\,
            I => \N__21314\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__21314\,
            I => \N__21311\
        );

    \I__4853\ : Span4Mux_s0_h
    port map (
            O => \N__21311\,
            I => \N__21307\
        );

    \I__4852\ : IoInMux
    port map (
            O => \N__21310\,
            I => \N__21304\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__21307\,
            I => \N__21300\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21297\
        );

    \I__4849\ : IoInMux
    port map (
            O => \N__21303\,
            I => \N__21294\
        );

    \I__4848\ : Span4Mux_v
    port map (
            O => \N__21300\,
            I => \N__21289\
        );

    \I__4847\ : Span4Mux_s3_v
    port map (
            O => \N__21297\,
            I => \N__21289\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__21294\,
            I => \N__21286\
        );

    \I__4845\ : Sp12to4
    port map (
            O => \N__21289\,
            I => \N__21283\
        );

    \I__4844\ : Span12Mux_s9_v
    port map (
            O => \N__21286\,
            I => \N__21280\
        );

    \I__4843\ : Span12Mux_h
    port map (
            O => \N__21283\,
            I => \N__21277\
        );

    \I__4842\ : Odrv12
    port map (
            O => \N__21280\,
            I => n1809
        );

    \I__4841\ : Odrv12
    port map (
            O => \N__21277\,
            I => n1809
        );

    \I__4840\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21269\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__21260\,
            I => \line_buffer.n464\
        );

    \I__4835\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__4833\ : Span4Mux_v
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__4832\ : Span4Mux_h
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__4831\ : Span4Mux_h
    port map (
            O => \N__21245\,
            I => \N__21242\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__21242\,
            I => \line_buffer.n456\
        );

    \I__4829\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21236\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__21236\,
            I => \line_buffer.n3497\
        );

    \I__4827\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21230\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__21230\,
            I => \N__21227\
        );

    \I__4825\ : Span4Mux_v
    port map (
            O => \N__21227\,
            I => \N__21224\
        );

    \I__4824\ : Span4Mux_v
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__4823\ : Sp12to4
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__21218\,
            I => \line_buffer.n524\
        );

    \I__4821\ : InMux
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__21212\,
            I => \N__21209\
        );

    \I__4819\ : Odrv12
    port map (
            O => \N__21209\,
            I => \line_buffer.n516\
        );

    \I__4818\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__4816\ : Span4Mux_v
    port map (
            O => \N__21200\,
            I => \N__21197\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__4814\ : Sp12to4
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__4813\ : Odrv12
    port map (
            O => \N__21191\,
            I => \line_buffer.n560\
        );

    \I__4812\ : InMux
    port map (
            O => \N__21188\,
            I => \N__21185\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__4810\ : Odrv12
    port map (
            O => \N__21182\,
            I => \line_buffer.n552\
        );

    \I__4809\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21176\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__21176\,
            I => \N__21173\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__4806\ : Odrv4
    port map (
            O => \N__21170\,
            I => \transmit_module.X_DELTA_PATTERN_1\
        );

    \I__4805\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__21164\,
            I => \transmit_module.X_DELTA_PATTERN_2\
        );

    \I__4803\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__21158\,
            I => \transmit_module.X_DELTA_PATTERN_3\
        );

    \I__4801\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__21152\,
            I => \transmit_module.X_DELTA_PATTERN_5\
        );

    \I__4799\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__21146\,
            I => \transmit_module.X_DELTA_PATTERN_4\
        );

    \I__4797\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__21140\,
            I => \transmit_module.X_DELTA_PATTERN_7\
        );

    \I__4795\ : InMux
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__21134\,
            I => \transmit_module.X_DELTA_PATTERN_6\
        );

    \I__4793\ : CEMux
    port map (
            O => \N__21131\,
            I => \N__21126\
        );

    \I__4792\ : CEMux
    port map (
            O => \N__21130\,
            I => \N__21123\
        );

    \I__4791\ : CEMux
    port map (
            O => \N__21129\,
            I => \N__21120\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__21126\,
            I => \N__21112\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__21123\,
            I => \N__21112\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__21120\,
            I => \N__21108\
        );

    \I__4787\ : CEMux
    port map (
            O => \N__21119\,
            I => \N__21105\
        );

    \I__4786\ : CEMux
    port map (
            O => \N__21118\,
            I => \N__21102\
        );

    \I__4785\ : CEMux
    port map (
            O => \N__21117\,
            I => \N__21099\
        );

    \I__4784\ : Span4Mux_v
    port map (
            O => \N__21112\,
            I => \N__21096\
        );

    \I__4783\ : CEMux
    port map (
            O => \N__21111\,
            I => \N__21093\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__21108\,
            I => \N__21086\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__21105\,
            I => \N__21086\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__21102\,
            I => \N__21086\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21083\
        );

    \I__4778\ : Span4Mux_h
    port map (
            O => \N__21096\,
            I => \N__21080\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__21093\,
            I => \N__21077\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__21086\,
            I => \N__21074\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__21083\,
            I => \transmit_module.n2115\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__21080\,
            I => \transmit_module.n2115\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__21077\,
            I => \transmit_module.n2115\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__21074\,
            I => \transmit_module.n2115\
        );

    \I__4771\ : SRMux
    port map (
            O => \N__21065\,
            I => \N__21058\
        );

    \I__4770\ : SRMux
    port map (
            O => \N__21064\,
            I => \N__21051\
        );

    \I__4769\ : SRMux
    port map (
            O => \N__21063\,
            I => \N__21048\
        );

    \I__4768\ : CEMux
    port map (
            O => \N__21062\,
            I => \N__21043\
        );

    \I__4767\ : CEMux
    port map (
            O => \N__21061\,
            I => \N__21040\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21037\
        );

    \I__4765\ : SRMux
    port map (
            O => \N__21057\,
            I => \N__21034\
        );

    \I__4764\ : CEMux
    port map (
            O => \N__21056\,
            I => \N__21029\
        );

    \I__4763\ : SRMux
    port map (
            O => \N__21055\,
            I => \N__21026\
        );

    \I__4762\ : SRMux
    port map (
            O => \N__21054\,
            I => \N__21023\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__21051\,
            I => \N__21019\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__21048\,
            I => \N__21016\
        );

    \I__4759\ : CEMux
    port map (
            O => \N__21047\,
            I => \N__21013\
        );

    \I__4758\ : CEMux
    port map (
            O => \N__21046\,
            I => \N__21010\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__21043\,
            I => \N__21006\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__21040\,
            I => \N__21003\
        );

    \I__4755\ : Span4Mux_h
    port map (
            O => \N__21037\,
            I => \N__21000\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__21034\,
            I => \N__20997\
        );

    \I__4753\ : CEMux
    port map (
            O => \N__21033\,
            I => \N__20994\
        );

    \I__4752\ : CEMux
    port map (
            O => \N__21032\,
            I => \N__20991\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__20987\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__20984\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__21023\,
            I => \N__20981\
        );

    \I__4748\ : CEMux
    port map (
            O => \N__21022\,
            I => \N__20978\
        );

    \I__4747\ : Span4Mux_h
    port map (
            O => \N__21019\,
            I => \N__20973\
        );

    \I__4746\ : Span4Mux_h
    port map (
            O => \N__21016\,
            I => \N__20973\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__21013\,
            I => \N__20968\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__21010\,
            I => \N__20968\
        );

    \I__4743\ : CEMux
    port map (
            O => \N__21009\,
            I => \N__20965\
        );

    \I__4742\ : Span4Mux_h
    port map (
            O => \N__21006\,
            I => \N__20956\
        );

    \I__4741\ : Span4Mux_v
    port map (
            O => \N__21003\,
            I => \N__20956\
        );

    \I__4740\ : Span4Mux_v
    port map (
            O => \N__21000\,
            I => \N__20956\
        );

    \I__4739\ : Span4Mux_h
    port map (
            O => \N__20997\,
            I => \N__20956\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__20994\,
            I => \N__20953\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__20991\,
            I => \N__20950\
        );

    \I__4736\ : CEMux
    port map (
            O => \N__20990\,
            I => \N__20947\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__20987\,
            I => \N__20940\
        );

    \I__4734\ : Span4Mux_h
    port map (
            O => \N__20984\,
            I => \N__20940\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__20981\,
            I => \N__20940\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20937\
        );

    \I__4731\ : Span4Mux_h
    port map (
            O => \N__20973\,
            I => \N__20934\
        );

    \I__4730\ : Span4Mux_h
    port map (
            O => \N__20968\,
            I => \N__20927\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__20965\,
            I => \N__20927\
        );

    \I__4728\ : Span4Mux_h
    port map (
            O => \N__20956\,
            I => \N__20927\
        );

    \I__4727\ : Span4Mux_v
    port map (
            O => \N__20953\,
            I => \N__20918\
        );

    \I__4726\ : Span4Mux_h
    port map (
            O => \N__20950\,
            I => \N__20918\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__20947\,
            I => \N__20918\
        );

    \I__4724\ : Span4Mux_h
    port map (
            O => \N__20940\,
            I => \N__20918\
        );

    \I__4723\ : Odrv12
    port map (
            O => \N__20937\,
            I => \transmit_module.n3635\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__20934\,
            I => \transmit_module.n3635\
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__20927\,
            I => \transmit_module.n3635\
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__20918\,
            I => \transmit_module.n3635\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__4717\ : Span4Mux_h
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__20897\,
            I => \line_buffer.n463\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__4712\ : Span12Mux_h
    port map (
            O => \N__20888\,
            I => \N__20885\
        );

    \I__4711\ : Span12Mux_v
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__4710\ : Odrv12
    port map (
            O => \N__20882\,
            I => \line_buffer.n455\
        );

    \I__4709\ : CascadeMux
    port map (
            O => \N__20879\,
            I => \N__20872\
        );

    \I__4708\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20865\
        );

    \I__4707\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20862\
        );

    \I__4706\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20859\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__20875\,
            I => \N__20856\
        );

    \I__4704\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20850\
        );

    \I__4703\ : InMux
    port map (
            O => \N__20871\,
            I => \N__20850\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20845\
        );

    \I__4701\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20845\
        );

    \I__4700\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20842\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20865\,
            I => \N__20836\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__20862\,
            I => \N__20833\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__20859\,
            I => \N__20830\
        );

    \I__4696\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20825\
        );

    \I__4695\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20825\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20812\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__20845\,
            I => \N__20812\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__20842\,
            I => \N__20809\
        );

    \I__4691\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20806\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20801\
        );

    \I__4689\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20801\
        );

    \I__4688\ : Span4Mux_s3_v
    port map (
            O => \N__20836\,
            I => \N__20798\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__20833\,
            I => \N__20793\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__20830\,
            I => \N__20793\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__20825\,
            I => \N__20790\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20787\
        );

    \I__4683\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20782\
        );

    \I__4682\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20782\
        );

    \I__4681\ : InMux
    port map (
            O => \N__20821\,
            I => \N__20773\
        );

    \I__4680\ : InMux
    port map (
            O => \N__20820\,
            I => \N__20773\
        );

    \I__4679\ : InMux
    port map (
            O => \N__20819\,
            I => \N__20773\
        );

    \I__4678\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20773\
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__20817\,
            I => \N__20766\
        );

    \I__4676\ : Span4Mux_h
    port map (
            O => \N__20812\,
            I => \N__20756\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__20809\,
            I => \N__20756\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__20806\,
            I => \N__20756\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__20801\,
            I => \N__20753\
        );

    \I__4672\ : Sp12to4
    port map (
            O => \N__20798\,
            I => \N__20748\
        );

    \I__4671\ : Sp12to4
    port map (
            O => \N__20793\,
            I => \N__20748\
        );

    \I__4670\ : Span4Mux_h
    port map (
            O => \N__20790\,
            I => \N__20743\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__20787\,
            I => \N__20743\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__20782\,
            I => \N__20738\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__20773\,
            I => \N__20738\
        );

    \I__4666\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20731\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20731\
        );

    \I__4664\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20731\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20728\
        );

    \I__4662\ : InMux
    port map (
            O => \N__20766\,
            I => \N__20725\
        );

    \I__4661\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20720\
        );

    \I__4660\ : InMux
    port map (
            O => \N__20764\,
            I => \N__20720\
        );

    \I__4659\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20717\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__20756\,
            I => \N__20712\
        );

    \I__4657\ : Span4Mux_v
    port map (
            O => \N__20753\,
            I => \N__20712\
        );

    \I__4656\ : Span12Mux_v
    port map (
            O => \N__20748\,
            I => \N__20709\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__20743\,
            I => \N__20704\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__20738\,
            I => \N__20704\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__20731\,
            I => \transmit_module.n3627\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__20728\,
            I => \transmit_module.n3627\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__20725\,
            I => \transmit_module.n3627\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__20720\,
            I => \transmit_module.n3627\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__20717\,
            I => \transmit_module.n3627\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__20712\,
            I => \transmit_module.n3627\
        );

    \I__4647\ : Odrv12
    port map (
            O => \N__20709\,
            I => \transmit_module.n3627\
        );

    \I__4646\ : Odrv4
    port map (
            O => \N__20704\,
            I => \transmit_module.n3627\
        );

    \I__4645\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20684\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__20684\,
            I => \N__20681\
        );

    \I__4643\ : Span4Mux_v
    port map (
            O => \N__20681\,
            I => \N__20678\
        );

    \I__4642\ : Span4Mux_h
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__20672\,
            I => \line_buffer.n556\
        );

    \I__4639\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20666\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__20666\,
            I => \N__20663\
        );

    \I__4637\ : Span12Mux_v
    port map (
            O => \N__20663\,
            I => \N__20660\
        );

    \I__4636\ : Odrv12
    port map (
            O => \N__20660\,
            I => \line_buffer.n548\
        );

    \I__4635\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20649\
        );

    \I__4634\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20646\
        );

    \I__4633\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20643\
        );

    \I__4632\ : InMux
    port map (
            O => \N__20654\,
            I => \N__20636\
        );

    \I__4631\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20636\
        );

    \I__4630\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20636\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__20649\,
            I => \N__20631\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__20646\,
            I => \N__20628\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20625\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__20636\,
            I => \N__20622\
        );

    \I__4625\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20617\
        );

    \I__4624\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20614\
        );

    \I__4623\ : Span12Mux_h
    port map (
            O => \N__20631\,
            I => \N__20607\
        );

    \I__4622\ : Span4Mux_h
    port map (
            O => \N__20628\,
            I => \N__20604\
        );

    \I__4621\ : Span12Mux_h
    port map (
            O => \N__20625\,
            I => \N__20601\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__20622\,
            I => \N__20598\
        );

    \I__4619\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20595\
        );

    \I__4618\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20592\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__20617\,
            I => \N__20587\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__20614\,
            I => \N__20587\
        );

    \I__4615\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20584\
        );

    \I__4614\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20577\
        );

    \I__4613\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20577\
        );

    \I__4612\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20577\
        );

    \I__4611\ : Odrv12
    port map (
            O => \N__20607\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__20604\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4609\ : Odrv12
    port map (
            O => \N__20601\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__20598\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__20595\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__20592\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4605\ : Odrv4
    port map (
            O => \N__20587\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__20584\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__20577\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4602\ : CascadeMux
    port map (
            O => \N__20558\,
            I => \N__20554\
        );

    \I__4601\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20551\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20548\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20545\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__20548\,
            I => \N__20542\
        );

    \I__4597\ : Span12Mux_h
    port map (
            O => \N__20545\,
            I => \N__20539\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__20542\,
            I => \N__20536\
        );

    \I__4595\ : Span12Mux_v
    port map (
            O => \N__20539\,
            I => \N__20533\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__20536\,
            I => \transmit_module.n112\
        );

    \I__4593\ : Odrv12
    port map (
            O => \N__20533\,
            I => \transmit_module.n112\
        );

    \I__4592\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20525\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__20525\,
            I => \N__20520\
        );

    \I__4590\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20517\
        );

    \I__4589\ : CascadeMux
    port map (
            O => \N__20523\,
            I => \N__20513\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__20520\,
            I => \N__20508\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__20517\,
            I => \N__20508\
        );

    \I__4586\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20505\
        );

    \I__4585\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20502\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__20508\,
            I => \N__20499\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20496\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__20502\,
            I => \N__20493\
        );

    \I__4581\ : Odrv4
    port map (
            O => \N__20499\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4580\ : Odrv12
    port map (
            O => \N__20496\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__20493\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4578\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20483\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__20483\,
            I => \transmit_module.ADDR_Y_COMPONENT_4\
        );

    \I__4576\ : CEMux
    port map (
            O => \N__20480\,
            I => \N__20476\
        );

    \I__4575\ : CEMux
    port map (
            O => \N__20479\,
            I => \N__20473\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__20476\,
            I => \N__20469\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__20473\,
            I => \N__20466\
        );

    \I__4572\ : CEMux
    port map (
            O => \N__20472\,
            I => \N__20463\
        );

    \I__4571\ : Span4Mux_h
    port map (
            O => \N__20469\,
            I => \N__20456\
        );

    \I__4570\ : Span4Mux_h
    port map (
            O => \N__20466\,
            I => \N__20456\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__20463\,
            I => \N__20456\
        );

    \I__4568\ : Span4Mux_v
    port map (
            O => \N__20456\,
            I => \N__20451\
        );

    \I__4567\ : CEMux
    port map (
            O => \N__20455\,
            I => \N__20448\
        );

    \I__4566\ : CEMux
    port map (
            O => \N__20454\,
            I => \N__20445\
        );

    \I__4565\ : Span4Mux_h
    port map (
            O => \N__20451\,
            I => \N__20439\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__20448\,
            I => \N__20439\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__20445\,
            I => \N__20436\
        );

    \I__4562\ : CEMux
    port map (
            O => \N__20444\,
            I => \N__20433\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__20439\,
            I => \N__20430\
        );

    \I__4560\ : Span12Mux_v
    port map (
            O => \N__20436\,
            I => \N__20425\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__20433\,
            I => \N__20425\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__20430\,
            I => \transmit_module.n2069\
        );

    \I__4557\ : Odrv12
    port map (
            O => \N__20425\,
            I => \transmit_module.n2069\
        );

    \I__4556\ : IoInMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__20417\,
            I => \N__20410\
        );

    \I__4554\ : SRMux
    port map (
            O => \N__20416\,
            I => \N__20404\
        );

    \I__4553\ : SRMux
    port map (
            O => \N__20415\,
            I => \N__20401\
        );

    \I__4552\ : SRMux
    port map (
            O => \N__20414\,
            I => \N__20398\
        );

    \I__4551\ : SRMux
    port map (
            O => \N__20413\,
            I => \N__20394\
        );

    \I__4550\ : Span4Mux_s1_h
    port map (
            O => \N__20410\,
            I => \N__20389\
        );

    \I__4549\ : SRMux
    port map (
            O => \N__20409\,
            I => \N__20386\
        );

    \I__4548\ : CascadeMux
    port map (
            O => \N__20408\,
            I => \N__20381\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__20407\,
            I => \N__20378\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__20404\,
            I => \N__20375\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__20401\,
            I => \N__20372\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__20398\,
            I => \N__20369\
        );

    \I__4543\ : SRMux
    port map (
            O => \N__20397\,
            I => \N__20366\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__20394\,
            I => \N__20363\
        );

    \I__4541\ : SRMux
    port map (
            O => \N__20393\,
            I => \N__20360\
        );

    \I__4540\ : SRMux
    port map (
            O => \N__20392\,
            I => \N__20357\
        );

    \I__4539\ : Span4Mux_h
    port map (
            O => \N__20389\,
            I => \N__20349\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__20386\,
            I => \N__20346\
        );

    \I__4537\ : SRMux
    port map (
            O => \N__20385\,
            I => \N__20343\
        );

    \I__4536\ : SRMux
    port map (
            O => \N__20384\,
            I => \N__20340\
        );

    \I__4535\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20332\
        );

    \I__4534\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20329\
        );

    \I__4533\ : Span4Mux_h
    port map (
            O => \N__20375\,
            I => \N__20321\
        );

    \I__4532\ : Span4Mux_v
    port map (
            O => \N__20372\,
            I => \N__20321\
        );

    \I__4531\ : Span4Mux_h
    port map (
            O => \N__20369\,
            I => \N__20316\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__20366\,
            I => \N__20316\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__20363\,
            I => \N__20309\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__20360\,
            I => \N__20309\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__20357\,
            I => \N__20309\
        );

    \I__4526\ : SRMux
    port map (
            O => \N__20356\,
            I => \N__20306\
        );

    \I__4525\ : CascadeMux
    port map (
            O => \N__20355\,
            I => \N__20302\
        );

    \I__4524\ : SRMux
    port map (
            O => \N__20354\,
            I => \N__20299\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__20353\,
            I => \N__20289\
        );

    \I__4522\ : SRMux
    port map (
            O => \N__20352\,
            I => \N__20281\
        );

    \I__4521\ : Span4Mux_v
    port map (
            O => \N__20349\,
            I => \N__20272\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__20346\,
            I => \N__20272\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__20343\,
            I => \N__20272\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__20340\,
            I => \N__20272\
        );

    \I__4517\ : SRMux
    port map (
            O => \N__20339\,
            I => \N__20269\
        );

    \I__4516\ : SRMux
    port map (
            O => \N__20338\,
            I => \N__20264\
        );

    \I__4515\ : SRMux
    port map (
            O => \N__20337\,
            I => \N__20261\
        );

    \I__4514\ : SRMux
    port map (
            O => \N__20336\,
            I => \N__20255\
        );

    \I__4513\ : SRMux
    port map (
            O => \N__20335\,
            I => \N__20252\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__20332\,
            I => \N__20247\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__20329\,
            I => \N__20244\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__20328\,
            I => \N__20241\
        );

    \I__4509\ : SRMux
    port map (
            O => \N__20327\,
            I => \N__20233\
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__20326\,
            I => \N__20230\
        );

    \I__4507\ : Span4Mux_v
    port map (
            O => \N__20321\,
            I => \N__20220\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__20316\,
            I => \N__20220\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__20309\,
            I => \N__20220\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__20306\,
            I => \N__20220\
        );

    \I__4503\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20217\
        );

    \I__4502\ : InMux
    port map (
            O => \N__20302\,
            I => \N__20214\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20211\
        );

    \I__4500\ : SRMux
    port map (
            O => \N__20298\,
            I => \N__20208\
        );

    \I__4499\ : SRMux
    port map (
            O => \N__20297\,
            I => \N__20205\
        );

    \I__4498\ : SRMux
    port map (
            O => \N__20296\,
            I => \N__20202\
        );

    \I__4497\ : SRMux
    port map (
            O => \N__20295\,
            I => \N__20199\
        );

    \I__4496\ : SRMux
    port map (
            O => \N__20294\,
            I => \N__20196\
        );

    \I__4495\ : SRMux
    port map (
            O => \N__20293\,
            I => \N__20193\
        );

    \I__4494\ : SRMux
    port map (
            O => \N__20292\,
            I => \N__20190\
        );

    \I__4493\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20183\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__20288\,
            I => \N__20180\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__20287\,
            I => \N__20176\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__20286\,
            I => \N__20173\
        );

    \I__4489\ : SRMux
    port map (
            O => \N__20285\,
            I => \N__20165\
        );

    \I__4488\ : SRMux
    port map (
            O => \N__20284\,
            I => \N__20160\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20157\
        );

    \I__4486\ : Span4Mux_h
    port map (
            O => \N__20272\,
            I => \N__20152\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__20269\,
            I => \N__20152\
        );

    \I__4484\ : SRMux
    port map (
            O => \N__20268\,
            I => \N__20149\
        );

    \I__4483\ : SRMux
    port map (
            O => \N__20267\,
            I => \N__20146\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__20264\,
            I => \N__20141\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__20261\,
            I => \N__20141\
        );

    \I__4480\ : SRMux
    port map (
            O => \N__20260\,
            I => \N__20138\
        );

    \I__4479\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20135\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__20258\,
            I => \N__20132\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__20255\,
            I => \N__20127\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__20252\,
            I => \N__20127\
        );

    \I__4475\ : SRMux
    port map (
            O => \N__20251\,
            I => \N__20124\
        );

    \I__4474\ : SRMux
    port map (
            O => \N__20250\,
            I => \N__20118\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__20247\,
            I => \N__20113\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__20244\,
            I => \N__20113\
        );

    \I__4471\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20110\
        );

    \I__4470\ : SRMux
    port map (
            O => \N__20240\,
            I => \N__20107\
        );

    \I__4469\ : SRMux
    port map (
            O => \N__20239\,
            I => \N__20104\
        );

    \I__4468\ : SRMux
    port map (
            O => \N__20238\,
            I => \N__20101\
        );

    \I__4467\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20096\
        );

    \I__4466\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20096\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__20233\,
            I => \N__20093\
        );

    \I__4464\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20090\
        );

    \I__4463\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20087\
        );

    \I__4462\ : Span4Mux_h
    port map (
            O => \N__20220\,
            I => \N__20080\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__20217\,
            I => \N__20080\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__20214\,
            I => \N__20080\
        );

    \I__4459\ : Span4Mux_v
    port map (
            O => \N__20211\,
            I => \N__20075\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__20208\,
            I => \N__20075\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__20205\,
            I => \N__20070\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__20202\,
            I => \N__20070\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__20199\,
            I => \N__20061\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__20196\,
            I => \N__20061\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20061\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__20190\,
            I => \N__20061\
        );

    \I__4451\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20058\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__20188\,
            I => \N__20055\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__20187\,
            I => \N__20052\
        );

    \I__4448\ : SRMux
    port map (
            O => \N__20186\,
            I => \N__20049\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__20183\,
            I => \N__20046\
        );

    \I__4446\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20043\
        );

    \I__4445\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20038\
        );

    \I__4444\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20038\
        );

    \I__4443\ : InMux
    port map (
            O => \N__20173\,
            I => \N__20029\
        );

    \I__4442\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20029\
        );

    \I__4441\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20029\
        );

    \I__4440\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20029\
        );

    \I__4439\ : SRMux
    port map (
            O => \N__20169\,
            I => \N__20026\
        );

    \I__4438\ : SRMux
    port map (
            O => \N__20168\,
            I => \N__20023\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__20165\,
            I => \N__20020\
        );

    \I__4436\ : SRMux
    port map (
            O => \N__20164\,
            I => \N__20017\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__20163\,
            I => \N__20012\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20007\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__20157\,
            I => \N__20007\
        );

    \I__4432\ : Span4Mux_h
    port map (
            O => \N__20152\,
            I => \N__20002\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__20149\,
            I => \N__20002\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__20146\,
            I => \N__19995\
        );

    \I__4429\ : Span4Mux_v
    port map (
            O => \N__20141\,
            I => \N__19995\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__20138\,
            I => \N__19995\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__20135\,
            I => \N__19992\
        );

    \I__4426\ : InMux
    port map (
            O => \N__20132\,
            I => \N__19989\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__20127\,
            I => \N__19984\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__20124\,
            I => \N__19984\
        );

    \I__4423\ : InMux
    port map (
            O => \N__20123\,
            I => \N__19981\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__20122\,
            I => \N__19978\
        );

    \I__4421\ : CascadeMux
    port map (
            O => \N__20121\,
            I => \N__19975\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__20118\,
            I => \N__19972\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__20113\,
            I => \N__19969\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__20110\,
            I => \N__19966\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__20107\,
            I => \N__19963\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__19956\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__20101\,
            I => \N__19956\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__20096\,
            I => \N__19956\
        );

    \I__4413\ : Span4Mux_v
    port map (
            O => \N__20093\,
            I => \N__19951\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__20090\,
            I => \N__19951\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__20087\,
            I => \N__19946\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__20080\,
            I => \N__19946\
        );

    \I__4409\ : Span4Mux_h
    port map (
            O => \N__20075\,
            I => \N__19939\
        );

    \I__4408\ : Span4Mux_v
    port map (
            O => \N__20070\,
            I => \N__19939\
        );

    \I__4407\ : Span4Mux_v
    port map (
            O => \N__20061\,
            I => \N__19939\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__20058\,
            I => \N__19936\
        );

    \I__4405\ : InMux
    port map (
            O => \N__20055\,
            I => \N__19931\
        );

    \I__4404\ : InMux
    port map (
            O => \N__20052\,
            I => \N__19931\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__20049\,
            I => \N__19920\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__20046\,
            I => \N__19920\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__19920\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__20038\,
            I => \N__19920\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__20029\,
            I => \N__19920\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__20026\,
            I => \N__19915\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__19915\
        );

    \I__4396\ : Span4Mux_h
    port map (
            O => \N__20020\,
            I => \N__19910\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__20017\,
            I => \N__19910\
        );

    \I__4394\ : InMux
    port map (
            O => \N__20016\,
            I => \N__19907\
        );

    \I__4393\ : InMux
    port map (
            O => \N__20015\,
            I => \N__19902\
        );

    \I__4392\ : InMux
    port map (
            O => \N__20012\,
            I => \N__19902\
        );

    \I__4391\ : Span4Mux_h
    port map (
            O => \N__20007\,
            I => \N__19895\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__20002\,
            I => \N__19895\
        );

    \I__4389\ : Span4Mux_h
    port map (
            O => \N__19995\,
            I => \N__19895\
        );

    \I__4388\ : Span4Mux_h
    port map (
            O => \N__19992\,
            I => \N__19890\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__19989\,
            I => \N__19890\
        );

    \I__4386\ : Span4Mux_h
    port map (
            O => \N__19984\,
            I => \N__19885\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19981\,
            I => \N__19885\
        );

    \I__4384\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19882\
        );

    \I__4383\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19879\
        );

    \I__4382\ : Span12Mux_h
    port map (
            O => \N__19972\,
            I => \N__19872\
        );

    \I__4381\ : Sp12to4
    port map (
            O => \N__19969\,
            I => \N__19872\
        );

    \I__4380\ : Span12Mux_s4_v
    port map (
            O => \N__19966\,
            I => \N__19872\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__19963\,
            I => \N__19863\
        );

    \I__4378\ : Span4Mux_v
    port map (
            O => \N__19956\,
            I => \N__19863\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__19951\,
            I => \N__19863\
        );

    \I__4376\ : Span4Mux_h
    port map (
            O => \N__19946\,
            I => \N__19863\
        );

    \I__4375\ : Span4Mux_h
    port map (
            O => \N__19939\,
            I => \N__19854\
        );

    \I__4374\ : Span4Mux_v
    port map (
            O => \N__19936\,
            I => \N__19854\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__19931\,
            I => \N__19854\
        );

    \I__4372\ : Span4Mux_v
    port map (
            O => \N__19920\,
            I => \N__19854\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__19915\,
            I => \N__19845\
        );

    \I__4370\ : Span4Mux_h
    port map (
            O => \N__19910\,
            I => \N__19845\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19845\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__19902\,
            I => \N__19845\
        );

    \I__4367\ : Odrv4
    port map (
            O => \N__19895\,
            I => \ADV_VSYNC_c\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__19890\,
            I => \ADV_VSYNC_c\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__19885\,
            I => \ADV_VSYNC_c\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19882\,
            I => \ADV_VSYNC_c\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19879\,
            I => \ADV_VSYNC_c\
        );

    \I__4362\ : Odrv12
    port map (
            O => \N__19872\,
            I => \ADV_VSYNC_c\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__19863\,
            I => \ADV_VSYNC_c\
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__19854\,
            I => \ADV_VSYNC_c\
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__19845\,
            I => \ADV_VSYNC_c\
        );

    \I__4358\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__4356\ : Span4Mux_v
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__4355\ : Sp12to4
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__4354\ : Odrv12
    port map (
            O => \N__19814\,
            I => \line_buffer.n529\
        );

    \I__4353\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__4351\ : Span12Mux_v
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__4350\ : Span12Mux_v
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__4349\ : Odrv12
    port map (
            O => \N__19799\,
            I => \line_buffer.n521\
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__19796\,
            I => \line_buffer.n3500_cascade_\
        );

    \I__4347\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__4345\ : Span4Mux_h
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__19784\,
            I => \line_buffer.n3501\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__19781\,
            I => \line_buffer.n3537_cascade_\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19774\
        );

    \I__4341\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19771\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__19774\,
            I => \N__19767\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19771\,
            I => \N__19762\
        );

    \I__4338\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19759\
        );

    \I__4337\ : Span4Mux_s1_v
    port map (
            O => \N__19767\,
            I => \N__19756\
        );

    \I__4336\ : InMux
    port map (
            O => \N__19766\,
            I => \N__19752\
        );

    \I__4335\ : InMux
    port map (
            O => \N__19765\,
            I => \N__19749\
        );

    \I__4334\ : Span4Mux_v
    port map (
            O => \N__19762\,
            I => \N__19743\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__19759\,
            I => \N__19743\
        );

    \I__4332\ : Span4Mux_h
    port map (
            O => \N__19756\,
            I => \N__19739\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19736\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__19752\,
            I => \N__19733\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__19749\,
            I => \N__19730\
        );

    \I__4328\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19727\
        );

    \I__4327\ : Span4Mux_v
    port map (
            O => \N__19743\,
            I => \N__19724\
        );

    \I__4326\ : InMux
    port map (
            O => \N__19742\,
            I => \N__19721\
        );

    \I__4325\ : Span4Mux_h
    port map (
            O => \N__19739\,
            I => \N__19718\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__19736\,
            I => \N__19715\
        );

    \I__4323\ : Span4Mux_v
    port map (
            O => \N__19733\,
            I => \N__19712\
        );

    \I__4322\ : Span4Mux_v
    port map (
            O => \N__19730\,
            I => \N__19707\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19727\,
            I => \N__19707\
        );

    \I__4320\ : Span4Mux_v
    port map (
            O => \N__19724\,
            I => \N__19702\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19721\,
            I => \N__19702\
        );

    \I__4318\ : Sp12to4
    port map (
            O => \N__19718\,
            I => \N__19697\
        );

    \I__4317\ : Span12Mux_h
    port map (
            O => \N__19715\,
            I => \N__19697\
        );

    \I__4316\ : Span4Mux_v
    port map (
            O => \N__19712\,
            I => \N__19692\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__19707\,
            I => \N__19692\
        );

    \I__4314\ : Span4Mux_h
    port map (
            O => \N__19702\,
            I => \N__19689\
        );

    \I__4313\ : Span12Mux_v
    port map (
            O => \N__19697\,
            I => \N__19686\
        );

    \I__4312\ : Sp12to4
    port map (
            O => \N__19692\,
            I => \N__19683\
        );

    \I__4311\ : Span4Mux_h
    port map (
            O => \N__19689\,
            I => \N__19680\
        );

    \I__4310\ : Odrv12
    port map (
            O => \N__19686\,
            I => \RX_DATA_2\
        );

    \I__4309\ : Odrv12
    port map (
            O => \N__19683\,
            I => \RX_DATA_2\
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__19680\,
            I => \RX_DATA_2\
        );

    \I__4307\ : CascadeMux
    port map (
            O => \N__19673\,
            I => \N__19669\
        );

    \I__4306\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19666\
        );

    \I__4305\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19663\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__19666\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__19663\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19655\,
            I => \transmit_module.X_DELTA_PATTERN_10\
        );

    \I__4300\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19649\,
            I => \transmit_module.X_DELTA_PATTERN_15\
        );

    \I__4298\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__19643\,
            I => \transmit_module.X_DELTA_PATTERN_14\
        );

    \I__4296\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__19637\,
            I => \transmit_module.X_DELTA_PATTERN_13\
        );

    \I__4294\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__19631\,
            I => \transmit_module.X_DELTA_PATTERN_12\
        );

    \I__4292\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__19625\,
            I => \transmit_module.X_DELTA_PATTERN_11\
        );

    \I__4290\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19619\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__19619\,
            I => \transmit_module.X_DELTA_PATTERN_9\
        );

    \I__4288\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__19613\,
            I => \transmit_module.X_DELTA_PATTERN_8\
        );

    \I__4286\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__4284\ : Odrv12
    port map (
            O => \N__19604\,
            I => \transmit_module.Y_DELTA_PATTERN_1\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__4282\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__4280\ : Span4Mux_h
    port map (
            O => \N__19592\,
            I => \N__19588\
        );

    \I__4279\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19585\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__19588\,
            I => \transmit_module.n108\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__19585\,
            I => \transmit_module.n108\
        );

    \I__4276\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__19577\,
            I => \N__19573\
        );

    \I__4274\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19570\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__19573\,
            I => \transmit_module.n139\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__19570\,
            I => \transmit_module.n139\
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__19565\,
            I => \N__19561\
        );

    \I__4270\ : CascadeMux
    port map (
            O => \N__19564\,
            I => \N__19558\
        );

    \I__4269\ : CascadeBuf
    port map (
            O => \N__19561\,
            I => \N__19555\
        );

    \I__4268\ : CascadeBuf
    port map (
            O => \N__19558\,
            I => \N__19552\
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__19555\,
            I => \N__19549\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__19552\,
            I => \N__19546\
        );

    \I__4265\ : CascadeBuf
    port map (
            O => \N__19549\,
            I => \N__19543\
        );

    \I__4264\ : CascadeBuf
    port map (
            O => \N__19546\,
            I => \N__19540\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__19543\,
            I => \N__19537\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__19540\,
            I => \N__19534\
        );

    \I__4261\ : CascadeBuf
    port map (
            O => \N__19537\,
            I => \N__19531\
        );

    \I__4260\ : CascadeBuf
    port map (
            O => \N__19534\,
            I => \N__19528\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__19531\,
            I => \N__19525\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__19528\,
            I => \N__19522\
        );

    \I__4257\ : CascadeBuf
    port map (
            O => \N__19525\,
            I => \N__19519\
        );

    \I__4256\ : CascadeBuf
    port map (
            O => \N__19522\,
            I => \N__19516\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__19519\,
            I => \N__19513\
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__19516\,
            I => \N__19510\
        );

    \I__4253\ : CascadeBuf
    port map (
            O => \N__19513\,
            I => \N__19507\
        );

    \I__4252\ : CascadeBuf
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__19507\,
            I => \N__19501\
        );

    \I__4250\ : CascadeMux
    port map (
            O => \N__19504\,
            I => \N__19498\
        );

    \I__4249\ : CascadeBuf
    port map (
            O => \N__19501\,
            I => \N__19495\
        );

    \I__4248\ : CascadeBuf
    port map (
            O => \N__19498\,
            I => \N__19492\
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__19495\,
            I => \N__19489\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__19492\,
            I => \N__19486\
        );

    \I__4245\ : CascadeBuf
    port map (
            O => \N__19489\,
            I => \N__19483\
        );

    \I__4244\ : CascadeBuf
    port map (
            O => \N__19486\,
            I => \N__19480\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__19483\,
            I => \N__19477\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__4241\ : CascadeBuf
    port map (
            O => \N__19477\,
            I => \N__19471\
        );

    \I__4240\ : CascadeBuf
    port map (
            O => \N__19474\,
            I => \N__19468\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__19471\,
            I => \N__19465\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__19468\,
            I => \N__19462\
        );

    \I__4237\ : CascadeBuf
    port map (
            O => \N__19465\,
            I => \N__19459\
        );

    \I__4236\ : CascadeBuf
    port map (
            O => \N__19462\,
            I => \N__19456\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__19459\,
            I => \N__19453\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__19456\,
            I => \N__19450\
        );

    \I__4233\ : CascadeBuf
    port map (
            O => \N__19453\,
            I => \N__19447\
        );

    \I__4232\ : CascadeBuf
    port map (
            O => \N__19450\,
            I => \N__19444\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__19447\,
            I => \N__19441\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__19444\,
            I => \N__19438\
        );

    \I__4229\ : CascadeBuf
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__4228\ : CascadeBuf
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__19432\,
            I => \N__19426\
        );

    \I__4225\ : CascadeBuf
    port map (
            O => \N__19429\,
            I => \N__19423\
        );

    \I__4224\ : CascadeBuf
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__19423\,
            I => \N__19417\
        );

    \I__4222\ : CascadeMux
    port map (
            O => \N__19420\,
            I => \N__19414\
        );

    \I__4221\ : CascadeBuf
    port map (
            O => \N__19417\,
            I => \N__19411\
        );

    \I__4220\ : CascadeBuf
    port map (
            O => \N__19414\,
            I => \N__19408\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__19411\,
            I => \N__19405\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__19408\,
            I => \N__19402\
        );

    \I__4217\ : CascadeBuf
    port map (
            O => \N__19405\,
            I => \N__19399\
        );

    \I__4216\ : CascadeBuf
    port map (
            O => \N__19402\,
            I => \N__19396\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__19399\,
            I => \N__19393\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__19396\,
            I => \N__19390\
        );

    \I__4213\ : CascadeBuf
    port map (
            O => \N__19393\,
            I => \N__19387\
        );

    \I__4212\ : CascadeBuf
    port map (
            O => \N__19390\,
            I => \N__19384\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__19387\,
            I => \N__19381\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__19384\,
            I => \N__19378\
        );

    \I__4209\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19375\
        );

    \I__4208\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19372\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__19375\,
            I => \N__19369\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__19372\,
            I => \N__19366\
        );

    \I__4205\ : Span4Mux_h
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__19366\,
            I => \N__19360\
        );

    \I__4203\ : Span4Mux_h
    port map (
            O => \N__19363\,
            I => \N__19357\
        );

    \I__4202\ : Sp12to4
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__4201\ : Sp12to4
    port map (
            O => \N__19357\,
            I => \N__19351\
        );

    \I__4200\ : Span12Mux_h
    port map (
            O => \N__19354\,
            I => \N__19346\
        );

    \I__4199\ : Span12Mux_s5_v
    port map (
            O => \N__19351\,
            I => \N__19346\
        );

    \I__4198\ : Odrv12
    port map (
            O => \N__19346\,
            I => n20
        );

    \I__4197\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__4195\ : Odrv4
    port map (
            O => \N__19337\,
            I => \transmit_module.ADDR_Y_COMPONENT_7\
        );

    \I__4194\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19329\
        );

    \I__4193\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19325\
        );

    \I__4192\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19322\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__19329\,
            I => \N__19319\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__19328\,
            I => \N__19316\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__19325\,
            I => \N__19311\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__19322\,
            I => \N__19311\
        );

    \I__4187\ : Span4Mux_v
    port map (
            O => \N__19319\,
            I => \N__19308\
        );

    \I__4186\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19305\
        );

    \I__4185\ : Odrv12
    port map (
            O => \N__19311\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__19308\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__19305\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__4182\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__19295\,
            I => \N__19291\
        );

    \I__4180\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19288\
        );

    \I__4179\ : Odrv12
    port map (
            O => \N__19291\,
            I => \transmit_module.n109\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__19288\,
            I => \transmit_module.n109\
        );

    \I__4177\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__19280\,
            I => \transmit_module.ADDR_Y_COMPONENT_6\
        );

    \I__4175\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__19274\,
            I => \N__19269\
        );

    \I__4173\ : InMux
    port map (
            O => \N__19273\,
            I => \N__19266\
        );

    \I__4172\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19263\
        );

    \I__4171\ : Span4Mux_v
    port map (
            O => \N__19269\,
            I => \N__19255\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__19266\,
            I => \N__19255\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__19263\,
            I => \N__19255\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__19262\,
            I => \N__19252\
        );

    \I__4167\ : Span4Mux_v
    port map (
            O => \N__19255\,
            I => \N__19249\
        );

    \I__4166\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19246\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__19249\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__19246\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__4163\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__19238\,
            I => \N__19234\
        );

    \I__4161\ : InMux
    port map (
            O => \N__19237\,
            I => \N__19231\
        );

    \I__4160\ : Odrv12
    port map (
            O => \N__19234\,
            I => \transmit_module.n110\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__19231\,
            I => \transmit_module.n110\
        );

    \I__4158\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__4156\ : Odrv4
    port map (
            O => \N__19220\,
            I => \transmit_module.ADDR_Y_COMPONENT_2\
        );

    \I__4155\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19212\
        );

    \I__4154\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19209\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__19215\,
            I => \N__19205\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__19212\,
            I => \N__19200\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__19209\,
            I => \N__19200\
        );

    \I__4150\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19197\
        );

    \I__4149\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19194\
        );

    \I__4148\ : Odrv12
    port map (
            O => \N__19200\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__19197\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__19194\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__4145\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__19181\,
            I => \transmit_module.ADDR_Y_COMPONENT_9\
        );

    \I__4142\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19174\
        );

    \I__4141\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19171\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__19174\,
            I => \N__19164\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__19171\,
            I => \N__19164\
        );

    \I__4138\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19161\
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__19169\,
            I => \N__19158\
        );

    \I__4136\ : Span4Mux_v
    port map (
            O => \N__19164\,
            I => \N__19155\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__19161\,
            I => \N__19152\
        );

    \I__4134\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19149\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__19155\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__4132\ : Odrv12
    port map (
            O => \N__19152\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__19149\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__4130\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__4127\ : Odrv4
    port map (
            O => \N__19133\,
            I => \transmit_module.n107\
        );

    \I__4126\ : CascadeMux
    port map (
            O => \N__19130\,
            I => \transmit_module.n107_cascade_\
        );

    \I__4125\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19120\
        );

    \I__4123\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19117\
        );

    \I__4122\ : Odrv12
    port map (
            O => \N__19120\,
            I => \transmit_module.n138\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__19117\,
            I => \transmit_module.n138\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__4119\ : CascadeBuf
    port map (
            O => \N__19109\,
            I => \N__19105\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__19108\,
            I => \N__19102\
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__19105\,
            I => \N__19099\
        );

    \I__4116\ : CascadeBuf
    port map (
            O => \N__19102\,
            I => \N__19096\
        );

    \I__4115\ : CascadeBuf
    port map (
            O => \N__19099\,
            I => \N__19093\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__19096\,
            I => \N__19090\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__19093\,
            I => \N__19087\
        );

    \I__4112\ : CascadeBuf
    port map (
            O => \N__19090\,
            I => \N__19084\
        );

    \I__4111\ : CascadeBuf
    port map (
            O => \N__19087\,
            I => \N__19081\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__19084\,
            I => \N__19078\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__19081\,
            I => \N__19075\
        );

    \I__4108\ : CascadeBuf
    port map (
            O => \N__19078\,
            I => \N__19072\
        );

    \I__4107\ : CascadeBuf
    port map (
            O => \N__19075\,
            I => \N__19069\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__19072\,
            I => \N__19066\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__19069\,
            I => \N__19063\
        );

    \I__4104\ : CascadeBuf
    port map (
            O => \N__19066\,
            I => \N__19060\
        );

    \I__4103\ : CascadeBuf
    port map (
            O => \N__19063\,
            I => \N__19057\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__19060\,
            I => \N__19054\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__19057\,
            I => \N__19051\
        );

    \I__4100\ : CascadeBuf
    port map (
            O => \N__19054\,
            I => \N__19048\
        );

    \I__4099\ : CascadeBuf
    port map (
            O => \N__19051\,
            I => \N__19045\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__19048\,
            I => \N__19042\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__19045\,
            I => \N__19039\
        );

    \I__4096\ : CascadeBuf
    port map (
            O => \N__19042\,
            I => \N__19036\
        );

    \I__4095\ : CascadeBuf
    port map (
            O => \N__19039\,
            I => \N__19033\
        );

    \I__4094\ : CascadeMux
    port map (
            O => \N__19036\,
            I => \N__19030\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__19033\,
            I => \N__19027\
        );

    \I__4092\ : CascadeBuf
    port map (
            O => \N__19030\,
            I => \N__19024\
        );

    \I__4091\ : CascadeBuf
    port map (
            O => \N__19027\,
            I => \N__19021\
        );

    \I__4090\ : CascadeMux
    port map (
            O => \N__19024\,
            I => \N__19018\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__19021\,
            I => \N__19015\
        );

    \I__4088\ : CascadeBuf
    port map (
            O => \N__19018\,
            I => \N__19012\
        );

    \I__4087\ : CascadeBuf
    port map (
            O => \N__19015\,
            I => \N__19009\
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__19012\,
            I => \N__19006\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__19009\,
            I => \N__19003\
        );

    \I__4084\ : CascadeBuf
    port map (
            O => \N__19006\,
            I => \N__19000\
        );

    \I__4083\ : CascadeBuf
    port map (
            O => \N__19003\,
            I => \N__18997\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__19000\,
            I => \N__18994\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__18997\,
            I => \N__18991\
        );

    \I__4080\ : CascadeBuf
    port map (
            O => \N__18994\,
            I => \N__18988\
        );

    \I__4079\ : CascadeBuf
    port map (
            O => \N__18991\,
            I => \N__18985\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__18988\,
            I => \N__18982\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__18985\,
            I => \N__18979\
        );

    \I__4076\ : CascadeBuf
    port map (
            O => \N__18982\,
            I => \N__18976\
        );

    \I__4075\ : CascadeBuf
    port map (
            O => \N__18979\,
            I => \N__18973\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__18976\,
            I => \N__18970\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__18973\,
            I => \N__18967\
        );

    \I__4072\ : CascadeBuf
    port map (
            O => \N__18970\,
            I => \N__18964\
        );

    \I__4071\ : CascadeBuf
    port map (
            O => \N__18967\,
            I => \N__18961\
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__18964\,
            I => \N__18958\
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__18961\,
            I => \N__18955\
        );

    \I__4068\ : CascadeBuf
    port map (
            O => \N__18958\,
            I => \N__18952\
        );

    \I__4067\ : CascadeBuf
    port map (
            O => \N__18955\,
            I => \N__18949\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__18952\,
            I => \N__18946\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__18949\,
            I => \N__18943\
        );

    \I__4064\ : CascadeBuf
    port map (
            O => \N__18946\,
            I => \N__18940\
        );

    \I__4063\ : CascadeBuf
    port map (
            O => \N__18943\,
            I => \N__18937\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__18940\,
            I => \N__18934\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__18937\,
            I => \N__18931\
        );

    \I__4060\ : CascadeBuf
    port map (
            O => \N__18934\,
            I => \N__18928\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18931\,
            I => \N__18925\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__18928\,
            I => \N__18922\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__18925\,
            I => \N__18919\
        );

    \I__4056\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18916\
        );

    \I__4055\ : Span4Mux_v
    port map (
            O => \N__18919\,
            I => \N__18913\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__18916\,
            I => \N__18910\
        );

    \I__4053\ : Span4Mux_v
    port map (
            O => \N__18913\,
            I => \N__18907\
        );

    \I__4052\ : Span12Mux_h
    port map (
            O => \N__18910\,
            I => \N__18904\
        );

    \I__4051\ : Span4Mux_v
    port map (
            O => \N__18907\,
            I => \N__18901\
        );

    \I__4050\ : Span12Mux_v
    port map (
            O => \N__18904\,
            I => \N__18898\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__18901\,
            I => \N__18895\
        );

    \I__4048\ : Odrv12
    port map (
            O => \N__18898\,
            I => n19
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__18895\,
            I => n19
        );

    \I__4046\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18886\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18889\,
            I => \N__18883\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__18886\,
            I => \N__18880\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18883\,
            I => \N__18877\
        );

    \I__4042\ : Span12Mux_s2_v
    port map (
            O => \N__18880\,
            I => \N__18874\
        );

    \I__4041\ : Odrv12
    port map (
            O => \N__18877\,
            I => \transmit_module.n114\
        );

    \I__4040\ : Odrv12
    port map (
            O => \N__18874\,
            I => \transmit_module.n114\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__4037\ : Span12Mux_s6_v
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__4036\ : Span12Mux_v
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__4035\ : Odrv12
    port map (
            O => \N__18857\,
            I => \transmit_module.n145\
        );

    \I__4034\ : CascadeMux
    port map (
            O => \N__18854\,
            I => \N__18850\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__18853\,
            I => \N__18847\
        );

    \I__4032\ : CascadeBuf
    port map (
            O => \N__18850\,
            I => \N__18844\
        );

    \I__4031\ : CascadeBuf
    port map (
            O => \N__18847\,
            I => \N__18841\
        );

    \I__4030\ : CascadeMux
    port map (
            O => \N__18844\,
            I => \N__18838\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__4028\ : CascadeBuf
    port map (
            O => \N__18838\,
            I => \N__18832\
        );

    \I__4027\ : CascadeBuf
    port map (
            O => \N__18835\,
            I => \N__18829\
        );

    \I__4026\ : CascadeMux
    port map (
            O => \N__18832\,
            I => \N__18826\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__18829\,
            I => \N__18823\
        );

    \I__4024\ : CascadeBuf
    port map (
            O => \N__18826\,
            I => \N__18820\
        );

    \I__4023\ : CascadeBuf
    port map (
            O => \N__18823\,
            I => \N__18817\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__18820\,
            I => \N__18814\
        );

    \I__4021\ : CascadeMux
    port map (
            O => \N__18817\,
            I => \N__18811\
        );

    \I__4020\ : CascadeBuf
    port map (
            O => \N__18814\,
            I => \N__18808\
        );

    \I__4019\ : CascadeBuf
    port map (
            O => \N__18811\,
            I => \N__18805\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__18808\,
            I => \N__18802\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__18805\,
            I => \N__18799\
        );

    \I__4016\ : CascadeBuf
    port map (
            O => \N__18802\,
            I => \N__18796\
        );

    \I__4015\ : CascadeBuf
    port map (
            O => \N__18799\,
            I => \N__18793\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__18796\,
            I => \N__18790\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__18793\,
            I => \N__18787\
        );

    \I__4012\ : CascadeBuf
    port map (
            O => \N__18790\,
            I => \N__18784\
        );

    \I__4011\ : CascadeBuf
    port map (
            O => \N__18787\,
            I => \N__18781\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__18784\,
            I => \N__18778\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__18781\,
            I => \N__18775\
        );

    \I__4008\ : CascadeBuf
    port map (
            O => \N__18778\,
            I => \N__18772\
        );

    \I__4007\ : CascadeBuf
    port map (
            O => \N__18775\,
            I => \N__18769\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__18772\,
            I => \N__18766\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__18769\,
            I => \N__18763\
        );

    \I__4004\ : CascadeBuf
    port map (
            O => \N__18766\,
            I => \N__18760\
        );

    \I__4003\ : CascadeBuf
    port map (
            O => \N__18763\,
            I => \N__18757\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__18760\,
            I => \N__18754\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__18757\,
            I => \N__18751\
        );

    \I__4000\ : CascadeBuf
    port map (
            O => \N__18754\,
            I => \N__18748\
        );

    \I__3999\ : CascadeBuf
    port map (
            O => \N__18751\,
            I => \N__18745\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__18748\,
            I => \N__18742\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__18745\,
            I => \N__18739\
        );

    \I__3996\ : CascadeBuf
    port map (
            O => \N__18742\,
            I => \N__18736\
        );

    \I__3995\ : CascadeBuf
    port map (
            O => \N__18739\,
            I => \N__18733\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__18736\,
            I => \N__18730\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__18733\,
            I => \N__18727\
        );

    \I__3992\ : CascadeBuf
    port map (
            O => \N__18730\,
            I => \N__18724\
        );

    \I__3991\ : CascadeBuf
    port map (
            O => \N__18727\,
            I => \N__18721\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__18724\,
            I => \N__18718\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__18721\,
            I => \N__18715\
        );

    \I__3988\ : CascadeBuf
    port map (
            O => \N__18718\,
            I => \N__18712\
        );

    \I__3987\ : CascadeBuf
    port map (
            O => \N__18715\,
            I => \N__18709\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__18712\,
            I => \N__18706\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__18709\,
            I => \N__18703\
        );

    \I__3984\ : CascadeBuf
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__3983\ : CascadeBuf
    port map (
            O => \N__18703\,
            I => \N__18697\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__18700\,
            I => \N__18694\
        );

    \I__3981\ : CascadeMux
    port map (
            O => \N__18697\,
            I => \N__18691\
        );

    \I__3980\ : CascadeBuf
    port map (
            O => \N__18694\,
            I => \N__18688\
        );

    \I__3979\ : CascadeBuf
    port map (
            O => \N__18691\,
            I => \N__18685\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__18688\,
            I => \N__18682\
        );

    \I__3977\ : CascadeMux
    port map (
            O => \N__18685\,
            I => \N__18679\
        );

    \I__3976\ : CascadeBuf
    port map (
            O => \N__18682\,
            I => \N__18676\
        );

    \I__3975\ : CascadeBuf
    port map (
            O => \N__18679\,
            I => \N__18673\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__18676\,
            I => \N__18670\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__18673\,
            I => \N__18667\
        );

    \I__3972\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18664\
        );

    \I__3971\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18661\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__18664\,
            I => \N__18658\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__18661\,
            I => \N__18655\
        );

    \I__3968\ : Span4Mux_h
    port map (
            O => \N__18658\,
            I => \N__18652\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__18655\,
            I => \N__18649\
        );

    \I__3966\ : Span4Mux_h
    port map (
            O => \N__18652\,
            I => \N__18644\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__18649\,
            I => \N__18644\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__18644\,
            I => n26
        );

    \I__3963\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18638\,
            I => \N__18635\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__3960\ : Span4Mux_v
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__18629\,
            I => \tvp_video_buffer.BUFFER_1_4\
        );

    \I__3958\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18623\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__18623\,
            I => \transmit_module.Y_DELTA_PATTERN_17\
        );

    \I__3956\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__3954\ : Span4Mux_h
    port map (
            O => \N__18614\,
            I => \N__18611\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__18611\,
            I => \N__18608\
        );

    \I__3952\ : Odrv4
    port map (
            O => \N__18608\,
            I => \transmit_module.Y_DELTA_PATTERN_20\
        );

    \I__3951\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18602\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__18602\,
            I => \transmit_module.Y_DELTA_PATTERN_19\
        );

    \I__3949\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__18596\,
            I => \transmit_module.Y_DELTA_PATTERN_18\
        );

    \I__3947\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__18587\,
            I => \transmit_module.ADDR_Y_COMPONENT_13\
        );

    \I__3944\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__18581\,
            I => \transmit_module.ADDR_Y_COMPONENT_12\
        );

    \I__3942\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__18572\,
            I => \transmit_module.ADDR_Y_COMPONENT_11\
        );

    \I__3939\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18565\
        );

    \I__3938\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18562\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__18565\,
            I => \N__18553\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__18562\,
            I => \N__18553\
        );

    \I__3935\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18550\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18547\
        );

    \I__3933\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18544\
        );

    \I__3932\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18541\
        );

    \I__3931\ : Span4Mux_v
    port map (
            O => \N__18553\,
            I => \N__18533\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18533\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18533\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__18544\,
            I => \N__18529\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__18541\,
            I => \N__18526\
        );

    \I__3926\ : InMux
    port map (
            O => \N__18540\,
            I => \N__18523\
        );

    \I__3925\ : Span4Mux_v
    port map (
            O => \N__18533\,
            I => \N__18520\
        );

    \I__3924\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18517\
        );

    \I__3923\ : Span4Mux_v
    port map (
            O => \N__18529\,
            I => \N__18514\
        );

    \I__3922\ : Span4Mux_s2_v
    port map (
            O => \N__18526\,
            I => \N__18509\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__18523\,
            I => \N__18509\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__18520\,
            I => \N__18504\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__18517\,
            I => \N__18504\
        );

    \I__3918\ : Span4Mux_v
    port map (
            O => \N__18514\,
            I => \N__18501\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__18509\,
            I => \N__18498\
        );

    \I__3916\ : Span4Mux_v
    port map (
            O => \N__18504\,
            I => \N__18495\
        );

    \I__3915\ : Sp12to4
    port map (
            O => \N__18501\,
            I => \N__18492\
        );

    \I__3914\ : Span4Mux_h
    port map (
            O => \N__18498\,
            I => \N__18489\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__18495\,
            I => \N__18486\
        );

    \I__3912\ : Span12Mux_h
    port map (
            O => \N__18492\,
            I => \N__18483\
        );

    \I__3911\ : Span4Mux_h
    port map (
            O => \N__18489\,
            I => \N__18480\
        );

    \I__3910\ : Span4Mux_h
    port map (
            O => \N__18486\,
            I => \N__18477\
        );

    \I__3909\ : Odrv12
    port map (
            O => \N__18483\,
            I => \RX_DATA_6\
        );

    \I__3908\ : Odrv4
    port map (
            O => \N__18480\,
            I => \RX_DATA_6\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__18477\,
            I => \RX_DATA_6\
        );

    \I__3906\ : IoInMux
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__3904\ : IoSpan4Mux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__3903\ : Span4Mux_s3_h
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__3902\ : Sp12to4
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__3901\ : Span12Mux_v
    port map (
            O => \N__18455\,
            I => \N__18451\
        );

    \I__3900\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18448\
        );

    \I__3899\ : Span12Mux_h
    port map (
            O => \N__18451\,
            I => \N__18445\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__18448\,
            I => \N__18442\
        );

    \I__3897\ : Odrv12
    port map (
            O => \N__18445\,
            I => \DEBUG_c_6_c\
        );

    \I__3896\ : Odrv12
    port map (
            O => \N__18442\,
            I => \DEBUG_c_6_c\
        );

    \I__3895\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__18434\,
            I => \tvp_video_buffer.BUFFER_0_8\
        );

    \I__3893\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__18428\,
            I => \tvp_video_buffer.BUFFER_1_8\
        );

    \I__3891\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__18419\,
            I => \N__18415\
        );

    \I__3888\ : InMux
    port map (
            O => \N__18418\,
            I => \N__18412\
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__18415\,
            I => \transmit_module.n141\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__18412\,
            I => \transmit_module.n141\
        );

    \I__3885\ : CEMux
    port map (
            O => \N__18407\,
            I => \N__18403\
        );

    \I__3884\ : CEMux
    port map (
            O => \N__18406\,
            I => \N__18399\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__18403\,
            I => \N__18396\
        );

    \I__3882\ : CEMux
    port map (
            O => \N__18402\,
            I => \N__18393\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__18399\,
            I => \N__18388\
        );

    \I__3880\ : Span4Mux_h
    port map (
            O => \N__18396\,
            I => \N__18383\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__18393\,
            I => \N__18383\
        );

    \I__3878\ : CEMux
    port map (
            O => \N__18392\,
            I => \N__18379\
        );

    \I__3877\ : CEMux
    port map (
            O => \N__18391\,
            I => \N__18376\
        );

    \I__3876\ : Span4Mux_h
    port map (
            O => \N__18388\,
            I => \N__18371\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__18383\,
            I => \N__18371\
        );

    \I__3874\ : SRMux
    port map (
            O => \N__18382\,
            I => \N__18368\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__18379\,
            I => \N__18365\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__18376\,
            I => \N__18362\
        );

    \I__3871\ : Span4Mux_h
    port map (
            O => \N__18371\,
            I => \N__18357\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__18368\,
            I => \N__18357\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__18365\,
            I => \N__18354\
        );

    \I__3868\ : Span4Mux_v
    port map (
            O => \N__18362\,
            I => \N__18349\
        );

    \I__3867\ : Span4Mux_h
    port map (
            O => \N__18357\,
            I => \N__18349\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__18354\,
            I => \N__18346\
        );

    \I__3865\ : Span4Mux_h
    port map (
            O => \N__18349\,
            I => \N__18343\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__18346\,
            I => \transmit_module.n2167\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__18343\,
            I => \transmit_module.n2167\
        );

    \I__3862\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18335\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__3860\ : Span4Mux_v
    port map (
            O => \N__18332\,
            I => \N__18328\
        );

    \I__3859\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18325\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__18328\,
            I => \transmit_module.n140\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__18325\,
            I => \transmit_module.n140\
        );

    \I__3856\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18317\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__18317\,
            I => \transmit_module.n130\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__18314\,
            I => \transmit_module.n145_cascade_\
        );

    \I__3853\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18308\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__3851\ : Span4Mux_h
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__18302\,
            I => \transmit_module.Y_DELTA_PATTERN_16\
        );

    \I__3849\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__18296\,
            I => \N__18292\
        );

    \I__3847\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18289\
        );

    \I__3846\ : Span4Mux_h
    port map (
            O => \N__18292\,
            I => \N__18283\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__18289\,
            I => \N__18283\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__18288\,
            I => \N__18279\
        );

    \I__3843\ : Span4Mux_v
    port map (
            O => \N__18283\,
            I => \N__18276\
        );

    \I__3842\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18273\
        );

    \I__3841\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18270\
        );

    \I__3840\ : Odrv4
    port map (
            O => \N__18276\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__18273\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__18270\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3837\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18260\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__18260\,
            I => \transmit_module.ADDR_Y_COMPONENT_1\
        );

    \I__3835\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__3833\ : Span12Mux_v
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__3832\ : Odrv12
    port map (
            O => \N__18248\,
            I => \transmit_module.n128\
        );

    \I__3831\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18239\
        );

    \I__3829\ : Span4Mux_v
    port map (
            O => \N__18239\,
            I => \N__18235\
        );

    \I__3828\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18232\
        );

    \I__3827\ : Span4Mux_v
    port map (
            O => \N__18235\,
            I => \N__18229\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__18232\,
            I => \N__18226\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__18229\,
            I => \N__18223\
        );

    \I__3824\ : Odrv12
    port map (
            O => \N__18226\,
            I => \transmit_module.n143\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__18223\,
            I => \transmit_module.n143\
        );

    \I__3822\ : SRMux
    port map (
            O => \N__18218\,
            I => \N__18214\
        );

    \I__3821\ : SRMux
    port map (
            O => \N__18217\,
            I => \N__18209\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__18214\,
            I => \N__18204\
        );

    \I__3819\ : SRMux
    port map (
            O => \N__18213\,
            I => \N__18201\
        );

    \I__3818\ : SRMux
    port map (
            O => \N__18212\,
            I => \N__18198\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18193\
        );

    \I__3816\ : SRMux
    port map (
            O => \N__18208\,
            I => \N__18190\
        );

    \I__3815\ : SRMux
    port map (
            O => \N__18207\,
            I => \N__18187\
        );

    \I__3814\ : Span4Mux_s1_v
    port map (
            O => \N__18204\,
            I => \N__18178\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__18201\,
            I => \N__18178\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__18198\,
            I => \N__18178\
        );

    \I__3811\ : SRMux
    port map (
            O => \N__18197\,
            I => \N__18175\
        );

    \I__3810\ : SRMux
    port map (
            O => \N__18196\,
            I => \N__18172\
        );

    \I__3809\ : Span4Mux_s1_v
    port map (
            O => \N__18193\,
            I => \N__18163\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__18190\,
            I => \N__18163\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__18187\,
            I => \N__18163\
        );

    \I__3806\ : SRMux
    port map (
            O => \N__18186\,
            I => \N__18160\
        );

    \I__3805\ : SRMux
    port map (
            O => \N__18185\,
            I => \N__18157\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__18178\,
            I => \N__18148\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__18175\,
            I => \N__18148\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__18172\,
            I => \N__18148\
        );

    \I__3801\ : SRMux
    port map (
            O => \N__18171\,
            I => \N__18145\
        );

    \I__3800\ : SRMux
    port map (
            O => \N__18170\,
            I => \N__18142\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__18163\,
            I => \N__18133\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__18160\,
            I => \N__18133\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__18157\,
            I => \N__18133\
        );

    \I__3796\ : SRMux
    port map (
            O => \N__18156\,
            I => \N__18130\
        );

    \I__3795\ : SRMux
    port map (
            O => \N__18155\,
            I => \N__18127\
        );

    \I__3794\ : Span4Mux_v
    port map (
            O => \N__18148\,
            I => \N__18117\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__18145\,
            I => \N__18117\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__18142\,
            I => \N__18117\
        );

    \I__3791\ : SRMux
    port map (
            O => \N__18141\,
            I => \N__18114\
        );

    \I__3790\ : SRMux
    port map (
            O => \N__18140\,
            I => \N__18111\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__18133\,
            I => \N__18102\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__18130\,
            I => \N__18102\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__18127\,
            I => \N__18102\
        );

    \I__3786\ : SRMux
    port map (
            O => \N__18126\,
            I => \N__18099\
        );

    \I__3785\ : SRMux
    port map (
            O => \N__18125\,
            I => \N__18096\
        );

    \I__3784\ : SRMux
    port map (
            O => \N__18124\,
            I => \N__18090\
        );

    \I__3783\ : Span4Mux_v
    port map (
            O => \N__18117\,
            I => \N__18085\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__18114\,
            I => \N__18080\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__18111\,
            I => \N__18080\
        );

    \I__3780\ : SRMux
    port map (
            O => \N__18110\,
            I => \N__18077\
        );

    \I__3779\ : SRMux
    port map (
            O => \N__18109\,
            I => \N__18074\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__18102\,
            I => \N__18063\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__18099\,
            I => \N__18063\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__18096\,
            I => \N__18063\
        );

    \I__3775\ : SRMux
    port map (
            O => \N__18095\,
            I => \N__18060\
        );

    \I__3774\ : SRMux
    port map (
            O => \N__18094\,
            I => \N__18057\
        );

    \I__3773\ : SRMux
    port map (
            O => \N__18093\,
            I => \N__18054\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__18090\,
            I => \N__18047\
        );

    \I__3771\ : SRMux
    port map (
            O => \N__18089\,
            I => \N__18044\
        );

    \I__3770\ : SRMux
    port map (
            O => \N__18088\,
            I => \N__18041\
        );

    \I__3769\ : Span4Mux_v
    port map (
            O => \N__18085\,
            I => \N__18038\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__18080\,
            I => \N__18031\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__18077\,
            I => \N__18031\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__18074\,
            I => \N__18031\
        );

    \I__3765\ : SRMux
    port map (
            O => \N__18073\,
            I => \N__18028\
        );

    \I__3764\ : SRMux
    port map (
            O => \N__18072\,
            I => \N__18025\
        );

    \I__3763\ : IoInMux
    port map (
            O => \N__18071\,
            I => \N__18022\
        );

    \I__3762\ : IoInMux
    port map (
            O => \N__18070\,
            I => \N__18019\
        );

    \I__3761\ : Span4Mux_v
    port map (
            O => \N__18063\,
            I => \N__18012\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__18060\,
            I => \N__18012\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__18057\,
            I => \N__18012\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__18054\,
            I => \N__18009\
        );

    \I__3757\ : SRMux
    port map (
            O => \N__18053\,
            I => \N__18006\
        );

    \I__3756\ : SRMux
    port map (
            O => \N__18052\,
            I => \N__18003\
        );

    \I__3755\ : SRMux
    port map (
            O => \N__18051\,
            I => \N__18000\
        );

    \I__3754\ : SRMux
    port map (
            O => \N__18050\,
            I => \N__17997\
        );

    \I__3753\ : Span4Mux_s2_v
    port map (
            O => \N__18047\,
            I => \N__17990\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__18044\,
            I => \N__17990\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__18041\,
            I => \N__17990\
        );

    \I__3750\ : Span4Mux_v
    port map (
            O => \N__18038\,
            I => \N__17981\
        );

    \I__3749\ : Span4Mux_v
    port map (
            O => \N__18031\,
            I => \N__17981\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__18028\,
            I => \N__17981\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__18025\,
            I => \N__17981\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__18022\,
            I => \N__17976\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__18019\,
            I => \N__17976\
        );

    \I__3744\ : Span4Mux_v
    port map (
            O => \N__18012\,
            I => \N__17973\
        );

    \I__3743\ : Span4Mux_s2_v
    port map (
            O => \N__18009\,
            I => \N__17966\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__18006\,
            I => \N__17966\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__18003\,
            I => \N__17966\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__18000\,
            I => \N__17961\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17997\,
            I => \N__17961\
        );

    \I__3738\ : Span4Mux_v
    port map (
            O => \N__17990\,
            I => \N__17956\
        );

    \I__3737\ : Span4Mux_v
    port map (
            O => \N__17981\,
            I => \N__17956\
        );

    \I__3736\ : IoSpan4Mux
    port map (
            O => \N__17976\,
            I => \N__17953\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__17973\,
            I => \N__17950\
        );

    \I__3734\ : Span4Mux_v
    port map (
            O => \N__17966\,
            I => \N__17945\
        );

    \I__3733\ : Span4Mux_v
    port map (
            O => \N__17961\,
            I => \N__17945\
        );

    \I__3732\ : Span4Mux_h
    port map (
            O => \N__17956\,
            I => \N__17942\
        );

    \I__3731\ : Span4Mux_s2_v
    port map (
            O => \N__17953\,
            I => \N__17939\
        );

    \I__3730\ : Span4Mux_v
    port map (
            O => \N__17950\,
            I => \N__17934\
        );

    \I__3729\ : Span4Mux_h
    port map (
            O => \N__17945\,
            I => \N__17934\
        );

    \I__3728\ : Span4Mux_h
    port map (
            O => \N__17942\,
            I => \N__17929\
        );

    \I__3727\ : Span4Mux_v
    port map (
            O => \N__17939\,
            I => \N__17929\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__17934\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__17929\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3724\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__17921\,
            I => \N__17917\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17914\
        );

    \I__3721\ : Span4Mux_s3_v
    port map (
            O => \N__17917\,
            I => \N__17908\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__17914\,
            I => \N__17905\
        );

    \I__3719\ : InMux
    port map (
            O => \N__17913\,
            I => \N__17902\
        );

    \I__3718\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17899\
        );

    \I__3717\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17896\
        );

    \I__3716\ : Span4Mux_h
    port map (
            O => \N__17908\,
            I => \N__17893\
        );

    \I__3715\ : Span4Mux_v
    port map (
            O => \N__17905\,
            I => \N__17887\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__17902\,
            I => \N__17887\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__17899\,
            I => \N__17883\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17896\,
            I => \N__17879\
        );

    \I__3711\ : Sp12to4
    port map (
            O => \N__17893\,
            I => \N__17876\
        );

    \I__3710\ : InMux
    port map (
            O => \N__17892\,
            I => \N__17873\
        );

    \I__3709\ : Span4Mux_v
    port map (
            O => \N__17887\,
            I => \N__17870\
        );

    \I__3708\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17867\
        );

    \I__3707\ : Span4Mux_v
    port map (
            O => \N__17883\,
            I => \N__17864\
        );

    \I__3706\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17861\
        );

    \I__3705\ : Span12Mux_s9_h
    port map (
            O => \N__17879\,
            I => \N__17858\
        );

    \I__3704\ : Span12Mux_h
    port map (
            O => \N__17876\,
            I => \N__17855\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17852\
        );

    \I__3702\ : Span4Mux_v
    port map (
            O => \N__17870\,
            I => \N__17847\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__17867\,
            I => \N__17847\
        );

    \I__3700\ : Span4Mux_v
    port map (
            O => \N__17864\,
            I => \N__17842\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17842\
        );

    \I__3698\ : Span12Mux_v
    port map (
            O => \N__17858\,
            I => \N__17839\
        );

    \I__3697\ : Span12Mux_v
    port map (
            O => \N__17855\,
            I => \N__17834\
        );

    \I__3696\ : Span12Mux_s10_h
    port map (
            O => \N__17852\,
            I => \N__17834\
        );

    \I__3695\ : Span4Mux_v
    port map (
            O => \N__17847\,
            I => \N__17831\
        );

    \I__3694\ : Span4Mux_h
    port map (
            O => \N__17842\,
            I => \N__17828\
        );

    \I__3693\ : Span12Mux_v
    port map (
            O => \N__17839\,
            I => \N__17821\
        );

    \I__3692\ : Span12Mux_v
    port map (
            O => \N__17834\,
            I => \N__17821\
        );

    \I__3691\ : Sp12to4
    port map (
            O => \N__17831\,
            I => \N__17821\
        );

    \I__3690\ : Span4Mux_h
    port map (
            O => \N__17828\,
            I => \N__17818\
        );

    \I__3689\ : Odrv12
    port map (
            O => \N__17821\,
            I => \RX_DATA_3\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__17818\,
            I => \RX_DATA_3\
        );

    \I__3687\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17810\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__17810\,
            I => \tvp_video_buffer.BUFFER_0_5\
        );

    \I__3685\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17804\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__17804\,
            I => \tvp_video_buffer.BUFFER_1_5\
        );

    \I__3683\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17798\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__17798\,
            I => \tvp_video_buffer.BUFFER_0_6\
        );

    \I__3681\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__17792\,
            I => \tvp_video_buffer.BUFFER_1_6\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17785\
        );

    \I__3678\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17782\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__17785\,
            I => \N__17779\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__17782\,
            I => \N__17776\
        );

    \I__3675\ : Span4Mux_h
    port map (
            O => \N__17779\,
            I => \N__17771\
        );

    \I__3674\ : Span4Mux_v
    port map (
            O => \N__17776\,
            I => \N__17766\
        );

    \I__3673\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17763\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17758\
        );

    \I__3671\ : Sp12to4
    port map (
            O => \N__17771\,
            I => \N__17755\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17752\
        );

    \I__3669\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17749\
        );

    \I__3668\ : Span4Mux_v
    port map (
            O => \N__17766\,
            I => \N__17744\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__17763\,
            I => \N__17744\
        );

    \I__3666\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17741\
        );

    \I__3665\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17738\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17735\
        );

    \I__3663\ : Span12Mux_v
    port map (
            O => \N__17755\,
            I => \N__17732\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__17752\,
            I => \N__17729\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__17749\,
            I => \N__17726\
        );

    \I__3660\ : Sp12to4
    port map (
            O => \N__17744\,
            I => \N__17719\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__17741\,
            I => \N__17719\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__17738\,
            I => \N__17719\
        );

    \I__3657\ : Span4Mux_h
    port map (
            O => \N__17735\,
            I => \N__17716\
        );

    \I__3656\ : Span12Mux_v
    port map (
            O => \N__17732\,
            I => \N__17713\
        );

    \I__3655\ : Span12Mux_h
    port map (
            O => \N__17729\,
            I => \N__17708\
        );

    \I__3654\ : Span12Mux_h
    port map (
            O => \N__17726\,
            I => \N__17708\
        );

    \I__3653\ : Span12Mux_v
    port map (
            O => \N__17719\,
            I => \N__17705\
        );

    \I__3652\ : Span4Mux_h
    port map (
            O => \N__17716\,
            I => \N__17702\
        );

    \I__3651\ : Odrv12
    port map (
            O => \N__17713\,
            I => \RX_DATA_4\
        );

    \I__3650\ : Odrv12
    port map (
            O => \N__17708\,
            I => \RX_DATA_4\
        );

    \I__3649\ : Odrv12
    port map (
            O => \N__17705\,
            I => \RX_DATA_4\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__17702\,
            I => \RX_DATA_4\
        );

    \I__3647\ : InMux
    port map (
            O => \N__17693\,
            I => \N__17690\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__17690\,
            I => \tvp_video_buffer.BUFFER_1_7\
        );

    \I__3645\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__3643\ : Span4Mux_v
    port map (
            O => \N__17681\,
            I => \N__17678\
        );

    \I__3642\ : Span4Mux_v
    port map (
            O => \N__17678\,
            I => \N__17674\
        );

    \I__3641\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17668\
        );

    \I__3640\ : Span4Mux_v
    port map (
            O => \N__17674\,
            I => \N__17665\
        );

    \I__3639\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17662\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17659\
        );

    \I__3637\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17655\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__17668\,
            I => \N__17651\
        );

    \I__3635\ : Span4Mux_v
    port map (
            O => \N__17665\,
            I => \N__17646\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__17662\,
            I => \N__17646\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__17659\,
            I => \N__17642\
        );

    \I__3632\ : InMux
    port map (
            O => \N__17658\,
            I => \N__17639\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__17655\,
            I => \N__17636\
        );

    \I__3630\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17633\
        );

    \I__3629\ : Span4Mux_s2_v
    port map (
            O => \N__17651\,
            I => \N__17630\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__17646\,
            I => \N__17627\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17624\
        );

    \I__3626\ : Sp12to4
    port map (
            O => \N__17642\,
            I => \N__17621\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__17639\,
            I => \N__17618\
        );

    \I__3624\ : Span4Mux_v
    port map (
            O => \N__17636\,
            I => \N__17615\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__17633\,
            I => \N__17612\
        );

    \I__3622\ : Span4Mux_v
    port map (
            O => \N__17630\,
            I => \N__17605\
        );

    \I__3621\ : Span4Mux_v
    port map (
            O => \N__17627\,
            I => \N__17605\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__17624\,
            I => \N__17605\
        );

    \I__3619\ : Span12Mux_v
    port map (
            O => \N__17621\,
            I => \N__17600\
        );

    \I__3618\ : Sp12to4
    port map (
            O => \N__17618\,
            I => \N__17600\
        );

    \I__3617\ : Span4Mux_v
    port map (
            O => \N__17615\,
            I => \N__17597\
        );

    \I__3616\ : Sp12to4
    port map (
            O => \N__17612\,
            I => \N__17594\
        );

    \I__3615\ : Span4Mux_h
    port map (
            O => \N__17605\,
            I => \N__17591\
        );

    \I__3614\ : Span12Mux_v
    port map (
            O => \N__17600\,
            I => \N__17584\
        );

    \I__3613\ : Sp12to4
    port map (
            O => \N__17597\,
            I => \N__17584\
        );

    \I__3612\ : Span12Mux_s7_v
    port map (
            O => \N__17594\,
            I => \N__17584\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__17591\,
            I => \N__17581\
        );

    \I__3610\ : Odrv12
    port map (
            O => \N__17584\,
            I => \RX_DATA_5\
        );

    \I__3609\ : Odrv4
    port map (
            O => \N__17581\,
            I => \RX_DATA_5\
        );

    \I__3608\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__17570\,
            I => \transmit_module.n121\
        );

    \I__3605\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__17561\,
            I => \transmit_module.n119\
        );

    \I__3602\ : CEMux
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__17555\,
            I => \N__17552\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__17552\,
            I => \transmit_module.n2057\
        );

    \I__3599\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__3597\ : Odrv12
    port map (
            O => \N__17543\,
            I => \transmit_module.n124\
        );

    \I__3596\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17534\
        );

    \I__3594\ : Odrv12
    port map (
            O => \N__17534\,
            I => \transmit_module.n126\
        );

    \I__3593\ : InMux
    port map (
            O => \N__17531\,
            I => \N__17528\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__3591\ : Odrv12
    port map (
            O => \N__17525\,
            I => \transmit_module.n123\
        );

    \I__3590\ : InMux
    port map (
            O => \N__17522\,
            I => \N__17519\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__17519\,
            I => \N__17516\
        );

    \I__3588\ : Odrv12
    port map (
            O => \N__17516\,
            I => \transmit_module.n125\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__17513\,
            I => \N__17510\
        );

    \I__3586\ : CascadeBuf
    port map (
            O => \N__17510\,
            I => \N__17506\
        );

    \I__3585\ : CascadeMux
    port map (
            O => \N__17509\,
            I => \N__17503\
        );

    \I__3584\ : CascadeMux
    port map (
            O => \N__17506\,
            I => \N__17500\
        );

    \I__3583\ : CascadeBuf
    port map (
            O => \N__17503\,
            I => \N__17497\
        );

    \I__3582\ : CascadeBuf
    port map (
            O => \N__17500\,
            I => \N__17494\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__17497\,
            I => \N__17491\
        );

    \I__3580\ : CascadeMux
    port map (
            O => \N__17494\,
            I => \N__17488\
        );

    \I__3579\ : CascadeBuf
    port map (
            O => \N__17491\,
            I => \N__17485\
        );

    \I__3578\ : CascadeBuf
    port map (
            O => \N__17488\,
            I => \N__17482\
        );

    \I__3577\ : CascadeMux
    port map (
            O => \N__17485\,
            I => \N__17479\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__17482\,
            I => \N__17476\
        );

    \I__3575\ : CascadeBuf
    port map (
            O => \N__17479\,
            I => \N__17473\
        );

    \I__3574\ : CascadeBuf
    port map (
            O => \N__17476\,
            I => \N__17470\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__17473\,
            I => \N__17467\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__17470\,
            I => \N__17464\
        );

    \I__3571\ : CascadeBuf
    port map (
            O => \N__17467\,
            I => \N__17461\
        );

    \I__3570\ : CascadeBuf
    port map (
            O => \N__17464\,
            I => \N__17458\
        );

    \I__3569\ : CascadeMux
    port map (
            O => \N__17461\,
            I => \N__17455\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__17458\,
            I => \N__17452\
        );

    \I__3567\ : CascadeBuf
    port map (
            O => \N__17455\,
            I => \N__17449\
        );

    \I__3566\ : CascadeBuf
    port map (
            O => \N__17452\,
            I => \N__17446\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__17449\,
            I => \N__17443\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__17446\,
            I => \N__17440\
        );

    \I__3563\ : CascadeBuf
    port map (
            O => \N__17443\,
            I => \N__17437\
        );

    \I__3562\ : CascadeBuf
    port map (
            O => \N__17440\,
            I => \N__17434\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__17437\,
            I => \N__17431\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__17434\,
            I => \N__17428\
        );

    \I__3559\ : CascadeBuf
    port map (
            O => \N__17431\,
            I => \N__17425\
        );

    \I__3558\ : CascadeBuf
    port map (
            O => \N__17428\,
            I => \N__17422\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__17425\,
            I => \N__17419\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__17422\,
            I => \N__17416\
        );

    \I__3555\ : CascadeBuf
    port map (
            O => \N__17419\,
            I => \N__17413\
        );

    \I__3554\ : CascadeBuf
    port map (
            O => \N__17416\,
            I => \N__17410\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__17413\,
            I => \N__17407\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__17410\,
            I => \N__17404\
        );

    \I__3551\ : CascadeBuf
    port map (
            O => \N__17407\,
            I => \N__17401\
        );

    \I__3550\ : CascadeBuf
    port map (
            O => \N__17404\,
            I => \N__17398\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__17401\,
            I => \N__17395\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__17398\,
            I => \N__17392\
        );

    \I__3547\ : CascadeBuf
    port map (
            O => \N__17395\,
            I => \N__17389\
        );

    \I__3546\ : CascadeBuf
    port map (
            O => \N__17392\,
            I => \N__17386\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__17389\,
            I => \N__17383\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__17386\,
            I => \N__17380\
        );

    \I__3543\ : CascadeBuf
    port map (
            O => \N__17383\,
            I => \N__17377\
        );

    \I__3542\ : CascadeBuf
    port map (
            O => \N__17380\,
            I => \N__17374\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__17377\,
            I => \N__17371\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__17374\,
            I => \N__17368\
        );

    \I__3539\ : CascadeBuf
    port map (
            O => \N__17371\,
            I => \N__17365\
        );

    \I__3538\ : CascadeBuf
    port map (
            O => \N__17368\,
            I => \N__17362\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__17365\,
            I => \N__17359\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__17362\,
            I => \N__17356\
        );

    \I__3535\ : CascadeBuf
    port map (
            O => \N__17359\,
            I => \N__17353\
        );

    \I__3534\ : CascadeBuf
    port map (
            O => \N__17356\,
            I => \N__17350\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__17353\,
            I => \N__17347\
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__17350\,
            I => \N__17344\
        );

    \I__3531\ : CascadeBuf
    port map (
            O => \N__17347\,
            I => \N__17341\
        );

    \I__3530\ : CascadeBuf
    port map (
            O => \N__17344\,
            I => \N__17338\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__17341\,
            I => \N__17335\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__17338\,
            I => \N__17332\
        );

    \I__3527\ : CascadeBuf
    port map (
            O => \N__17335\,
            I => \N__17329\
        );

    \I__3526\ : InMux
    port map (
            O => \N__17332\,
            I => \N__17326\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__17329\,
            I => \N__17323\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__17326\,
            I => \N__17320\
        );

    \I__3523\ : InMux
    port map (
            O => \N__17323\,
            I => \N__17317\
        );

    \I__3522\ : Span4Mux_v
    port map (
            O => \N__17320\,
            I => \N__17314\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__17317\,
            I => \N__17311\
        );

    \I__3520\ : Span4Mux_v
    port map (
            O => \N__17314\,
            I => \N__17308\
        );

    \I__3519\ : Span4Mux_v
    port map (
            O => \N__17311\,
            I => \N__17305\
        );

    \I__3518\ : Span4Mux_v
    port map (
            O => \N__17308\,
            I => \N__17302\
        );

    \I__3517\ : Span4Mux_v
    port map (
            O => \N__17305\,
            I => \N__17299\
        );

    \I__3516\ : Span4Mux_h
    port map (
            O => \N__17302\,
            I => \N__17296\
        );

    \I__3515\ : Span4Mux_v
    port map (
            O => \N__17299\,
            I => \N__17293\
        );

    \I__3514\ : Span4Mux_h
    port map (
            O => \N__17296\,
            I => \N__17288\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__17293\,
            I => \N__17288\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__17288\,
            I => n22
        );

    \I__3511\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17282\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__17282\,
            I => \N__17279\
        );

    \I__3509\ : Odrv12
    port map (
            O => \N__17279\,
            I => \transmit_module.ADDR_Y_COMPONENT_8\
        );

    \I__3508\ : InMux
    port map (
            O => \N__17276\,
            I => \N__17273\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__17273\,
            I => \N__17268\
        );

    \I__3506\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17265\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__17271\,
            I => \N__17261\
        );

    \I__3504\ : Span4Mux_v
    port map (
            O => \N__17268\,
            I => \N__17256\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__17265\,
            I => \N__17256\
        );

    \I__3502\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17251\
        );

    \I__3501\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17251\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__17256\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__17251\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__17246\,
            I => \N__17242\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__17245\,
            I => \N__17239\
        );

    \I__3496\ : CascadeBuf
    port map (
            O => \N__17242\,
            I => \N__17236\
        );

    \I__3495\ : CascadeBuf
    port map (
            O => \N__17239\,
            I => \N__17233\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__17236\,
            I => \N__17230\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__17233\,
            I => \N__17227\
        );

    \I__3492\ : CascadeBuf
    port map (
            O => \N__17230\,
            I => \N__17224\
        );

    \I__3491\ : CascadeBuf
    port map (
            O => \N__17227\,
            I => \N__17221\
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__17224\,
            I => \N__17218\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__17221\,
            I => \N__17215\
        );

    \I__3488\ : CascadeBuf
    port map (
            O => \N__17218\,
            I => \N__17212\
        );

    \I__3487\ : CascadeBuf
    port map (
            O => \N__17215\,
            I => \N__17209\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__17212\,
            I => \N__17206\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__17209\,
            I => \N__17203\
        );

    \I__3484\ : CascadeBuf
    port map (
            O => \N__17206\,
            I => \N__17200\
        );

    \I__3483\ : CascadeBuf
    port map (
            O => \N__17203\,
            I => \N__17197\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__17200\,
            I => \N__17194\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__17197\,
            I => \N__17191\
        );

    \I__3480\ : CascadeBuf
    port map (
            O => \N__17194\,
            I => \N__17188\
        );

    \I__3479\ : CascadeBuf
    port map (
            O => \N__17191\,
            I => \N__17185\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__17188\,
            I => \N__17182\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__17185\,
            I => \N__17179\
        );

    \I__3476\ : CascadeBuf
    port map (
            O => \N__17182\,
            I => \N__17176\
        );

    \I__3475\ : CascadeBuf
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__3473\ : CascadeMux
    port map (
            O => \N__17173\,
            I => \N__17167\
        );

    \I__3472\ : CascadeBuf
    port map (
            O => \N__17170\,
            I => \N__17164\
        );

    \I__3471\ : CascadeBuf
    port map (
            O => \N__17167\,
            I => \N__17161\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__17164\,
            I => \N__17158\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__17161\,
            I => \N__17155\
        );

    \I__3468\ : CascadeBuf
    port map (
            O => \N__17158\,
            I => \N__17152\
        );

    \I__3467\ : CascadeBuf
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__17152\,
            I => \N__17146\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__17149\,
            I => \N__17143\
        );

    \I__3464\ : CascadeBuf
    port map (
            O => \N__17146\,
            I => \N__17140\
        );

    \I__3463\ : CascadeBuf
    port map (
            O => \N__17143\,
            I => \N__17137\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__17140\,
            I => \N__17134\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__3460\ : CascadeBuf
    port map (
            O => \N__17134\,
            I => \N__17128\
        );

    \I__3459\ : CascadeBuf
    port map (
            O => \N__17131\,
            I => \N__17125\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__17128\,
            I => \N__17122\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__17125\,
            I => \N__17119\
        );

    \I__3456\ : CascadeBuf
    port map (
            O => \N__17122\,
            I => \N__17116\
        );

    \I__3455\ : CascadeBuf
    port map (
            O => \N__17119\,
            I => \N__17113\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__17116\,
            I => \N__17110\
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__17113\,
            I => \N__17107\
        );

    \I__3452\ : CascadeBuf
    port map (
            O => \N__17110\,
            I => \N__17104\
        );

    \I__3451\ : CascadeBuf
    port map (
            O => \N__17107\,
            I => \N__17101\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__17104\,
            I => \N__17098\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__17101\,
            I => \N__17095\
        );

    \I__3448\ : CascadeBuf
    port map (
            O => \N__17098\,
            I => \N__17092\
        );

    \I__3447\ : CascadeBuf
    port map (
            O => \N__17095\,
            I => \N__17089\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__17092\,
            I => \N__17086\
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__17089\,
            I => \N__17083\
        );

    \I__3444\ : CascadeBuf
    port map (
            O => \N__17086\,
            I => \N__17080\
        );

    \I__3443\ : CascadeBuf
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__17080\,
            I => \N__17074\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__17077\,
            I => \N__17071\
        );

    \I__3440\ : CascadeBuf
    port map (
            O => \N__17074\,
            I => \N__17068\
        );

    \I__3439\ : CascadeBuf
    port map (
            O => \N__17071\,
            I => \N__17065\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__17068\,
            I => \N__17062\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__17065\,
            I => \N__17059\
        );

    \I__3436\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17056\
        );

    \I__3435\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17053\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__17056\,
            I => \N__17050\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__17053\,
            I => \N__17047\
        );

    \I__3432\ : Sp12to4
    port map (
            O => \N__17050\,
            I => \N__17044\
        );

    \I__3431\ : Span4Mux_h
    port map (
            O => \N__17047\,
            I => \N__17041\
        );

    \I__3430\ : Span12Mux_h
    port map (
            O => \N__17044\,
            I => \N__17038\
        );

    \I__3429\ : Sp12to4
    port map (
            O => \N__17041\,
            I => \N__17035\
        );

    \I__3428\ : Span12Mux_v
    port map (
            O => \N__17038\,
            I => \N__17030\
        );

    \I__3427\ : Span12Mux_v
    port map (
            O => \N__17035\,
            I => \N__17030\
        );

    \I__3426\ : Odrv12
    port map (
            O => \N__17030\,
            I => n21
        );

    \I__3425\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17024\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__17024\,
            I => \transmit_module.ADDR_Y_COMPONENT_5\
        );

    \I__3423\ : InMux
    port map (
            O => \N__17021\,
            I => \N__17017\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__17020\,
            I => \N__17012\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__17017\,
            I => \N__17009\
        );

    \I__3420\ : InMux
    port map (
            O => \N__17016\,
            I => \N__17006\
        );

    \I__3419\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17003\
        );

    \I__3418\ : InMux
    port map (
            O => \N__17012\,
            I => \N__17000\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__17009\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__17006\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__17003\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__17000\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__3413\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16988\,
            I => \transmit_module.n111\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__16985\,
            I => \transmit_module.n111_cascade_\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__16979\,
            I => \transmit_module.n142\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__3407\ : CascadeBuf
    port map (
            O => \N__16973\,
            I => \N__16969\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__16972\,
            I => \N__16966\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__16969\,
            I => \N__16963\
        );

    \I__3404\ : CascadeBuf
    port map (
            O => \N__16966\,
            I => \N__16960\
        );

    \I__3403\ : CascadeBuf
    port map (
            O => \N__16963\,
            I => \N__16957\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__16960\,
            I => \N__16954\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__16957\,
            I => \N__16951\
        );

    \I__3400\ : CascadeBuf
    port map (
            O => \N__16954\,
            I => \N__16948\
        );

    \I__3399\ : CascadeBuf
    port map (
            O => \N__16951\,
            I => \N__16945\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__16948\,
            I => \N__16942\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__16945\,
            I => \N__16939\
        );

    \I__3396\ : CascadeBuf
    port map (
            O => \N__16942\,
            I => \N__16936\
        );

    \I__3395\ : CascadeBuf
    port map (
            O => \N__16939\,
            I => \N__16933\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__16936\,
            I => \N__16930\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__16933\,
            I => \N__16927\
        );

    \I__3392\ : CascadeBuf
    port map (
            O => \N__16930\,
            I => \N__16924\
        );

    \I__3391\ : CascadeBuf
    port map (
            O => \N__16927\,
            I => \N__16921\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__16924\,
            I => \N__16918\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__16921\,
            I => \N__16915\
        );

    \I__3388\ : CascadeBuf
    port map (
            O => \N__16918\,
            I => \N__16912\
        );

    \I__3387\ : CascadeBuf
    port map (
            O => \N__16915\,
            I => \N__16909\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__16912\,
            I => \N__16906\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__16909\,
            I => \N__16903\
        );

    \I__3384\ : CascadeBuf
    port map (
            O => \N__16906\,
            I => \N__16900\
        );

    \I__3383\ : CascadeBuf
    port map (
            O => \N__16903\,
            I => \N__16897\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__16900\,
            I => \N__16894\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__16897\,
            I => \N__16891\
        );

    \I__3380\ : CascadeBuf
    port map (
            O => \N__16894\,
            I => \N__16888\
        );

    \I__3379\ : CascadeBuf
    port map (
            O => \N__16891\,
            I => \N__16885\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__16888\,
            I => \N__16882\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__16885\,
            I => \N__16879\
        );

    \I__3376\ : CascadeBuf
    port map (
            O => \N__16882\,
            I => \N__16876\
        );

    \I__3375\ : CascadeBuf
    port map (
            O => \N__16879\,
            I => \N__16873\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__16876\,
            I => \N__16870\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__16873\,
            I => \N__16867\
        );

    \I__3372\ : CascadeBuf
    port map (
            O => \N__16870\,
            I => \N__16864\
        );

    \I__3371\ : CascadeBuf
    port map (
            O => \N__16867\,
            I => \N__16861\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__16864\,
            I => \N__16858\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__16861\,
            I => \N__16855\
        );

    \I__3368\ : CascadeBuf
    port map (
            O => \N__16858\,
            I => \N__16852\
        );

    \I__3367\ : CascadeBuf
    port map (
            O => \N__16855\,
            I => \N__16849\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__16852\,
            I => \N__16846\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__16849\,
            I => \N__16843\
        );

    \I__3364\ : CascadeBuf
    port map (
            O => \N__16846\,
            I => \N__16840\
        );

    \I__3363\ : CascadeBuf
    port map (
            O => \N__16843\,
            I => \N__16837\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__16840\,
            I => \N__16834\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__16837\,
            I => \N__16831\
        );

    \I__3360\ : CascadeBuf
    port map (
            O => \N__16834\,
            I => \N__16828\
        );

    \I__3359\ : CascadeBuf
    port map (
            O => \N__16831\,
            I => \N__16825\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__16828\,
            I => \N__16822\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__16825\,
            I => \N__16819\
        );

    \I__3356\ : CascadeBuf
    port map (
            O => \N__16822\,
            I => \N__16816\
        );

    \I__3355\ : CascadeBuf
    port map (
            O => \N__16819\,
            I => \N__16813\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__16816\,
            I => \N__16810\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__16813\,
            I => \N__16807\
        );

    \I__3352\ : CascadeBuf
    port map (
            O => \N__16810\,
            I => \N__16804\
        );

    \I__3351\ : CascadeBuf
    port map (
            O => \N__16807\,
            I => \N__16801\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__16804\,
            I => \N__16798\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__16801\,
            I => \N__16795\
        );

    \I__3348\ : CascadeBuf
    port map (
            O => \N__16798\,
            I => \N__16792\
        );

    \I__3347\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16789\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__16792\,
            I => \N__16786\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16789\,
            I => \N__16783\
        );

    \I__3344\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16780\
        );

    \I__3343\ : Span4Mux_v
    port map (
            O => \N__16783\,
            I => \N__16777\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__16780\,
            I => \N__16774\
        );

    \I__3341\ : Span4Mux_v
    port map (
            O => \N__16777\,
            I => \N__16771\
        );

    \I__3340\ : Span4Mux_v
    port map (
            O => \N__16774\,
            I => \N__16768\
        );

    \I__3339\ : Span4Mux_v
    port map (
            O => \N__16771\,
            I => \N__16765\
        );

    \I__3338\ : Span4Mux_v
    port map (
            O => \N__16768\,
            I => \N__16762\
        );

    \I__3337\ : Span4Mux_v
    port map (
            O => \N__16765\,
            I => \N__16759\
        );

    \I__3336\ : Span4Mux_v
    port map (
            O => \N__16762\,
            I => \N__16756\
        );

    \I__3335\ : Span4Mux_h
    port map (
            O => \N__16759\,
            I => \N__16753\
        );

    \I__3334\ : Span4Mux_v
    port map (
            O => \N__16756\,
            I => \N__16750\
        );

    \I__3333\ : Span4Mux_h
    port map (
            O => \N__16753\,
            I => \N__16745\
        );

    \I__3332\ : Span4Mux_h
    port map (
            O => \N__16750\,
            I => \N__16745\
        );

    \I__3331\ : Odrv4
    port map (
            O => \N__16745\,
            I => n23
        );

    \I__3330\ : InMux
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__16739\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_580\
        );

    \I__3328\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16732\
        );

    \I__3327\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16729\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__16732\,
            I => \N__16726\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__16729\,
            I => \transmit_module.video_signal_controller.n3333\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__16726\,
            I => \transmit_module.video_signal_controller.n3333\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__3322\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16713\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16708\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16705\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__16713\,
            I => \N__16702\
        );

    \I__3318\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16697\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16697\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__16708\,
            I => \N__16694\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__16705\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__16702\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__16697\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__16694\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16682\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__3309\ : Span4Mux_h
    port map (
            O => \N__16679\,
            I => \N__16676\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__16676\,
            I => \transmit_module.video_signal_controller.n7\
        );

    \I__3307\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__16670\,
            I => \transmit_module.ADDR_Y_COMPONENT_10\
        );

    \I__3305\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16661\
        );

    \I__3304\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16658\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16655\
        );

    \I__3302\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16652\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__16661\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__16658\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__16655\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__16652\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16639\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16636\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__16639\,
            I => \N__16633\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__16636\,
            I => \transmit_module.n106\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__16633\,
            I => \transmit_module.n106\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16625\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__16622\,
            I => \transmit_module.n120\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16619\,
            I => \transmit_module.n3110\
        );

    \I__3288\ : InMux
    port map (
            O => \N__16616\,
            I => \bfn_15_14_0_\
        );

    \I__3287\ : InMux
    port map (
            O => \N__16613\,
            I => \transmit_module.n3112\
        );

    \I__3286\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16607\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__16607\,
            I => \transmit_module.n122\
        );

    \I__3284\ : InMux
    port map (
            O => \N__16604\,
            I => \transmit_module.n3113\
        );

    \I__3283\ : InMux
    port map (
            O => \N__16601\,
            I => \transmit_module.n3114\
        );

    \I__3282\ : InMux
    port map (
            O => \N__16598\,
            I => \transmit_module.n3115\
        );

    \I__3281\ : InMux
    port map (
            O => \N__16595\,
            I => \transmit_module.n3116\
        );

    \I__3280\ : IoInMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__16589\,
            I => \N__16586\
        );

    \I__3278\ : IoSpan4Mux
    port map (
            O => \N__16586\,
            I => \N__16583\
        );

    \I__3277\ : Span4Mux_s2_h
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__3276\ : Sp12to4
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__3275\ : Span12Mux_v
    port map (
            O => \N__16577\,
            I => \N__16573\
        );

    \I__3274\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16570\
        );

    \I__3273\ : Span12Mux_h
    port map (
            O => \N__16573\,
            I => \N__16567\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__16570\,
            I => \N__16564\
        );

    \I__3271\ : Odrv12
    port map (
            O => \N__16567\,
            I => \DEBUG_c_5_c\
        );

    \I__3270\ : Odrv12
    port map (
            O => \N__16564\,
            I => \DEBUG_c_5_c\
        );

    \I__3269\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16556\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__16556\,
            I => \tvp_video_buffer.BUFFER_0_7\
        );

    \I__3267\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16548\
        );

    \I__3266\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16545\
        );

    \I__3265\ : InMux
    port map (
            O => \N__16551\,
            I => \N__16541\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16536\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__16545\,
            I => \N__16536\
        );

    \I__3262\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16533\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__16541\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3260\ : Odrv12
    port map (
            O => \N__16536\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__16533\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3258\ : InMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__16523\,
            I => \transmit_module.n132\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3255\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__16514\,
            I => \transmit_module.n131\
        );

    \I__3253\ : InMux
    port map (
            O => \N__16511\,
            I => \transmit_module.n3104\
        );

    \I__3252\ : InMux
    port map (
            O => \N__16508\,
            I => \transmit_module.n3105\
        );

    \I__3251\ : InMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__16502\,
            I => \N__16498\
        );

    \I__3249\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16495\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__16498\,
            I => \N__16488\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__16495\,
            I => \N__16488\
        );

    \I__3246\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16485\
        );

    \I__3245\ : CascadeMux
    port map (
            O => \N__16493\,
            I => \N__16482\
        );

    \I__3244\ : Sp12to4
    port map (
            O => \N__16488\,
            I => \N__16477\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__16485\,
            I => \N__16477\
        );

    \I__3242\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16474\
        );

    \I__3241\ : Odrv12
    port map (
            O => \N__16477\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__16474\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3239\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__16460\,
            I => \transmit_module.n129\
        );

    \I__3235\ : InMux
    port map (
            O => \N__16457\,
            I => \transmit_module.n3106\
        );

    \I__3234\ : InMux
    port map (
            O => \N__16454\,
            I => \transmit_module.n3107\
        );

    \I__3233\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__16448\,
            I => \transmit_module.n127\
        );

    \I__3231\ : InMux
    port map (
            O => \N__16445\,
            I => \transmit_module.n3108\
        );

    \I__3230\ : InMux
    port map (
            O => \N__16442\,
            I => \transmit_module.n3109\
        );

    \I__3229\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__16436\,
            I => \N__16433\
        );

    \I__3227\ : Span4Mux_v
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__16430\,
            I => \transmit_module.ADDR_Y_COMPONENT_0\
        );

    \I__3225\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16424\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__16424\,
            I => \N__16418\
        );

    \I__3223\ : InMux
    port map (
            O => \N__16423\,
            I => \N__16415\
        );

    \I__3222\ : InMux
    port map (
            O => \N__16422\,
            I => \N__16410\
        );

    \I__3221\ : InMux
    port map (
            O => \N__16421\,
            I => \N__16410\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__16418\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__16415\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__16410\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3217\ : InMux
    port map (
            O => \N__16403\,
            I => \N__16400\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__16400\,
            I => \N__16394\
        );

    \I__3215\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16391\
        );

    \I__3214\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16386\
        );

    \I__3213\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16386\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__16394\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__16391\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__16386\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__3209\ : IoInMux
    port map (
            O => \N__16379\,
            I => \N__16376\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__16376\,
            I => \N__16373\
        );

    \I__3207\ : Span4Mux_s3_h
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__3206\ : Sp12to4
    port map (
            O => \N__16370\,
            I => \N__16366\
        );

    \I__3205\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16363\
        );

    \I__3204\ : Span12Mux_v
    port map (
            O => \N__16366\,
            I => \N__16356\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__16363\,
            I => \N__16353\
        );

    \I__3202\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16348\
        );

    \I__3201\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16348\
        );

    \I__3200\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16343\
        );

    \I__3199\ : InMux
    port map (
            O => \N__16359\,
            I => \N__16343\
        );

    \I__3198\ : Odrv12
    port map (
            O => \N__16356\,
            I => \ADV_HSYNC_c\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__16353\,
            I => \ADV_HSYNC_c\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__16348\,
            I => \ADV_HSYNC_c\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__16343\,
            I => \ADV_HSYNC_c\
        );

    \I__3194\ : InMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__3192\ : Odrv12
    port map (
            O => \N__16328\,
            I => \transmit_module.n137\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__16325\,
            I => \N__16322\
        );

    \I__3190\ : CascadeBuf
    port map (
            O => \N__16322\,
            I => \N__16318\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__16321\,
            I => \N__16315\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__16318\,
            I => \N__16312\
        );

    \I__3187\ : CascadeBuf
    port map (
            O => \N__16315\,
            I => \N__16309\
        );

    \I__3186\ : CascadeBuf
    port map (
            O => \N__16312\,
            I => \N__16306\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__16309\,
            I => \N__16303\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__16306\,
            I => \N__16300\
        );

    \I__3183\ : CascadeBuf
    port map (
            O => \N__16303\,
            I => \N__16297\
        );

    \I__3182\ : CascadeBuf
    port map (
            O => \N__16300\,
            I => \N__16294\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__16297\,
            I => \N__16291\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__16294\,
            I => \N__16288\
        );

    \I__3179\ : CascadeBuf
    port map (
            O => \N__16291\,
            I => \N__16285\
        );

    \I__3178\ : CascadeBuf
    port map (
            O => \N__16288\,
            I => \N__16282\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__16285\,
            I => \N__16279\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__16282\,
            I => \N__16276\
        );

    \I__3175\ : CascadeBuf
    port map (
            O => \N__16279\,
            I => \N__16273\
        );

    \I__3174\ : CascadeBuf
    port map (
            O => \N__16276\,
            I => \N__16270\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__16273\,
            I => \N__16267\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__16270\,
            I => \N__16264\
        );

    \I__3171\ : CascadeBuf
    port map (
            O => \N__16267\,
            I => \N__16261\
        );

    \I__3170\ : CascadeBuf
    port map (
            O => \N__16264\,
            I => \N__16258\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__16261\,
            I => \N__16255\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__16258\,
            I => \N__16252\
        );

    \I__3167\ : CascadeBuf
    port map (
            O => \N__16255\,
            I => \N__16249\
        );

    \I__3166\ : CascadeBuf
    port map (
            O => \N__16252\,
            I => \N__16246\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__16249\,
            I => \N__16243\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__16246\,
            I => \N__16240\
        );

    \I__3163\ : CascadeBuf
    port map (
            O => \N__16243\,
            I => \N__16237\
        );

    \I__3162\ : CascadeBuf
    port map (
            O => \N__16240\,
            I => \N__16234\
        );

    \I__3161\ : CascadeMux
    port map (
            O => \N__16237\,
            I => \N__16231\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__16234\,
            I => \N__16228\
        );

    \I__3159\ : CascadeBuf
    port map (
            O => \N__16231\,
            I => \N__16225\
        );

    \I__3158\ : CascadeBuf
    port map (
            O => \N__16228\,
            I => \N__16222\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__16225\,
            I => \N__16219\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__16222\,
            I => \N__16216\
        );

    \I__3155\ : CascadeBuf
    port map (
            O => \N__16219\,
            I => \N__16213\
        );

    \I__3154\ : CascadeBuf
    port map (
            O => \N__16216\,
            I => \N__16210\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__16213\,
            I => \N__16207\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__16210\,
            I => \N__16204\
        );

    \I__3151\ : CascadeBuf
    port map (
            O => \N__16207\,
            I => \N__16201\
        );

    \I__3150\ : CascadeBuf
    port map (
            O => \N__16204\,
            I => \N__16198\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__16201\,
            I => \N__16195\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__16198\,
            I => \N__16192\
        );

    \I__3147\ : CascadeBuf
    port map (
            O => \N__16195\,
            I => \N__16189\
        );

    \I__3146\ : CascadeBuf
    port map (
            O => \N__16192\,
            I => \N__16186\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__16189\,
            I => \N__16183\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__16186\,
            I => \N__16180\
        );

    \I__3143\ : CascadeBuf
    port map (
            O => \N__16183\,
            I => \N__16177\
        );

    \I__3142\ : CascadeBuf
    port map (
            O => \N__16180\,
            I => \N__16174\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__16177\,
            I => \N__16171\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__16174\,
            I => \N__16168\
        );

    \I__3139\ : CascadeBuf
    port map (
            O => \N__16171\,
            I => \N__16165\
        );

    \I__3138\ : CascadeBuf
    port map (
            O => \N__16168\,
            I => \N__16162\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__16165\,
            I => \N__16159\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__16162\,
            I => \N__16156\
        );

    \I__3135\ : CascadeBuf
    port map (
            O => \N__16159\,
            I => \N__16153\
        );

    \I__3134\ : CascadeBuf
    port map (
            O => \N__16156\,
            I => \N__16150\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__16153\,
            I => \N__16147\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__16150\,
            I => \N__16144\
        );

    \I__3131\ : CascadeBuf
    port map (
            O => \N__16147\,
            I => \N__16141\
        );

    \I__3130\ : InMux
    port map (
            O => \N__16144\,
            I => \N__16138\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__16141\,
            I => \N__16135\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__16138\,
            I => \N__16132\
        );

    \I__3127\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16129\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__16132\,
            I => \N__16126\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__16129\,
            I => \N__16123\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__16126\,
            I => \N__16120\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__16123\,
            I => \N__16117\
        );

    \I__3122\ : Span4Mux_v
    port map (
            O => \N__16120\,
            I => \N__16114\
        );

    \I__3121\ : Span4Mux_v
    port map (
            O => \N__16117\,
            I => \N__16111\
        );

    \I__3120\ : Span4Mux_h
    port map (
            O => \N__16114\,
            I => \N__16108\
        );

    \I__3119\ : Span4Mux_v
    port map (
            O => \N__16111\,
            I => \N__16105\
        );

    \I__3118\ : Span4Mux_h
    port map (
            O => \N__16108\,
            I => \N__16100\
        );

    \I__3117\ : Span4Mux_h
    port map (
            O => \N__16105\,
            I => \N__16100\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__16100\,
            I => n18
        );

    \I__3115\ : InMux
    port map (
            O => \N__16097\,
            I => \N__16094\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__16094\,
            I => \N__16090\
        );

    \I__3113\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16087\
        );

    \I__3112\ : Odrv12
    port map (
            O => \N__16090\,
            I => \transmit_module.n116\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__16087\,
            I => \transmit_module.n116\
        );

    \I__3110\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16078\
        );

    \I__3109\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16075\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__16078\,
            I => \N__16072\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__16075\,
            I => \transmit_module.n147\
        );

    \I__3106\ : Odrv12
    port map (
            O => \N__16072\,
            I => \transmit_module.n147\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__16067\,
            I => \N__16063\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__16066\,
            I => \N__16060\
        );

    \I__3103\ : CascadeBuf
    port map (
            O => \N__16063\,
            I => \N__16057\
        );

    \I__3102\ : CascadeBuf
    port map (
            O => \N__16060\,
            I => \N__16054\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__16057\,
            I => \N__16051\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__16054\,
            I => \N__16048\
        );

    \I__3099\ : CascadeBuf
    port map (
            O => \N__16051\,
            I => \N__16045\
        );

    \I__3098\ : CascadeBuf
    port map (
            O => \N__16048\,
            I => \N__16042\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__16045\,
            I => \N__16039\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__16042\,
            I => \N__16036\
        );

    \I__3095\ : CascadeBuf
    port map (
            O => \N__16039\,
            I => \N__16033\
        );

    \I__3094\ : CascadeBuf
    port map (
            O => \N__16036\,
            I => \N__16030\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__16033\,
            I => \N__16027\
        );

    \I__3092\ : CascadeMux
    port map (
            O => \N__16030\,
            I => \N__16024\
        );

    \I__3091\ : CascadeBuf
    port map (
            O => \N__16027\,
            I => \N__16021\
        );

    \I__3090\ : CascadeBuf
    port map (
            O => \N__16024\,
            I => \N__16018\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__16021\,
            I => \N__16015\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__16018\,
            I => \N__16012\
        );

    \I__3087\ : CascadeBuf
    port map (
            O => \N__16015\,
            I => \N__16009\
        );

    \I__3086\ : CascadeBuf
    port map (
            O => \N__16012\,
            I => \N__16006\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__16009\,
            I => \N__16003\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__16006\,
            I => \N__16000\
        );

    \I__3083\ : CascadeBuf
    port map (
            O => \N__16003\,
            I => \N__15997\
        );

    \I__3082\ : CascadeBuf
    port map (
            O => \N__16000\,
            I => \N__15994\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__15997\,
            I => \N__15991\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__15994\,
            I => \N__15988\
        );

    \I__3079\ : CascadeBuf
    port map (
            O => \N__15991\,
            I => \N__15985\
        );

    \I__3078\ : CascadeBuf
    port map (
            O => \N__15988\,
            I => \N__15982\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__15985\,
            I => \N__15979\
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__15982\,
            I => \N__15976\
        );

    \I__3075\ : CascadeBuf
    port map (
            O => \N__15979\,
            I => \N__15973\
        );

    \I__3074\ : CascadeBuf
    port map (
            O => \N__15976\,
            I => \N__15970\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__15973\,
            I => \N__15967\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__15970\,
            I => \N__15964\
        );

    \I__3071\ : CascadeBuf
    port map (
            O => \N__15967\,
            I => \N__15961\
        );

    \I__3070\ : CascadeBuf
    port map (
            O => \N__15964\,
            I => \N__15958\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__15961\,
            I => \N__15955\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__15958\,
            I => \N__15952\
        );

    \I__3067\ : CascadeBuf
    port map (
            O => \N__15955\,
            I => \N__15949\
        );

    \I__3066\ : CascadeBuf
    port map (
            O => \N__15952\,
            I => \N__15946\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__15949\,
            I => \N__15943\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__15946\,
            I => \N__15940\
        );

    \I__3063\ : CascadeBuf
    port map (
            O => \N__15943\,
            I => \N__15937\
        );

    \I__3062\ : CascadeBuf
    port map (
            O => \N__15940\,
            I => \N__15934\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__15937\,
            I => \N__15931\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__15934\,
            I => \N__15928\
        );

    \I__3059\ : CascadeBuf
    port map (
            O => \N__15931\,
            I => \N__15925\
        );

    \I__3058\ : CascadeBuf
    port map (
            O => \N__15928\,
            I => \N__15922\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__15925\,
            I => \N__15919\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__15922\,
            I => \N__15916\
        );

    \I__3055\ : CascadeBuf
    port map (
            O => \N__15919\,
            I => \N__15913\
        );

    \I__3054\ : CascadeBuf
    port map (
            O => \N__15916\,
            I => \N__15910\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__15913\,
            I => \N__15907\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__15910\,
            I => \N__15904\
        );

    \I__3051\ : CascadeBuf
    port map (
            O => \N__15907\,
            I => \N__15901\
        );

    \I__3050\ : CascadeBuf
    port map (
            O => \N__15904\,
            I => \N__15898\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__15901\,
            I => \N__15895\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__15898\,
            I => \N__15892\
        );

    \I__3047\ : CascadeBuf
    port map (
            O => \N__15895\,
            I => \N__15889\
        );

    \I__3046\ : CascadeBuf
    port map (
            O => \N__15892\,
            I => \N__15886\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__15889\,
            I => \N__15883\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__15886\,
            I => \N__15880\
        );

    \I__3043\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15877\
        );

    \I__3042\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15874\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__15877\,
            I => \N__15871\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15874\,
            I => \N__15868\
        );

    \I__3039\ : Span4Mux_s2_v
    port map (
            O => \N__15871\,
            I => \N__15865\
        );

    \I__3038\ : Span12Mux_s11_h
    port map (
            O => \N__15868\,
            I => \N__15862\
        );

    \I__3037\ : Sp12to4
    port map (
            O => \N__15865\,
            I => \N__15859\
        );

    \I__3036\ : Span12Mux_v
    port map (
            O => \N__15862\,
            I => \N__15854\
        );

    \I__3035\ : Span12Mux_v
    port map (
            O => \N__15859\,
            I => \N__15854\
        );

    \I__3034\ : Odrv12
    port map (
            O => \N__15854\,
            I => n28
        );

    \I__3033\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15847\
        );

    \I__3032\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15844\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__15847\,
            I => \N__15841\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__15844\,
            I => \N__15838\
        );

    \I__3029\ : Span12Mux_v
    port map (
            O => \N__15841\,
            I => \N__15833\
        );

    \I__3028\ : Span12Mux_s5_v
    port map (
            O => \N__15838\,
            I => \N__15833\
        );

    \I__3027\ : Odrv12
    port map (
            O => \N__15833\,
            I => \transmit_module.n115\
        );

    \I__3026\ : InMux
    port map (
            O => \N__15830\,
            I => \N__15827\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__15827\,
            I => \N__15823\
        );

    \I__3024\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15820\
        );

    \I__3023\ : Span12Mux_s10_v
    port map (
            O => \N__15823\,
            I => \N__15817\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__15820\,
            I => \transmit_module.n146\
        );

    \I__3021\ : Odrv12
    port map (
            O => \N__15817\,
            I => \transmit_module.n146\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__15812\,
            I => \N__15808\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__15811\,
            I => \N__15805\
        );

    \I__3018\ : CascadeBuf
    port map (
            O => \N__15808\,
            I => \N__15802\
        );

    \I__3017\ : CascadeBuf
    port map (
            O => \N__15805\,
            I => \N__15799\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__15802\,
            I => \N__15796\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__15799\,
            I => \N__15793\
        );

    \I__3014\ : CascadeBuf
    port map (
            O => \N__15796\,
            I => \N__15790\
        );

    \I__3013\ : CascadeBuf
    port map (
            O => \N__15793\,
            I => \N__15787\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__15790\,
            I => \N__15784\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__15787\,
            I => \N__15781\
        );

    \I__3010\ : CascadeBuf
    port map (
            O => \N__15784\,
            I => \N__15778\
        );

    \I__3009\ : CascadeBuf
    port map (
            O => \N__15781\,
            I => \N__15775\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__15778\,
            I => \N__15772\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__15775\,
            I => \N__15769\
        );

    \I__3006\ : CascadeBuf
    port map (
            O => \N__15772\,
            I => \N__15766\
        );

    \I__3005\ : CascadeBuf
    port map (
            O => \N__15769\,
            I => \N__15763\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__15766\,
            I => \N__15760\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__15763\,
            I => \N__15757\
        );

    \I__3002\ : CascadeBuf
    port map (
            O => \N__15760\,
            I => \N__15754\
        );

    \I__3001\ : CascadeBuf
    port map (
            O => \N__15757\,
            I => \N__15751\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__15754\,
            I => \N__15748\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__15751\,
            I => \N__15745\
        );

    \I__2998\ : CascadeBuf
    port map (
            O => \N__15748\,
            I => \N__15742\
        );

    \I__2997\ : CascadeBuf
    port map (
            O => \N__15745\,
            I => \N__15739\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__15742\,
            I => \N__15736\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__15739\,
            I => \N__15733\
        );

    \I__2994\ : CascadeBuf
    port map (
            O => \N__15736\,
            I => \N__15730\
        );

    \I__2993\ : CascadeBuf
    port map (
            O => \N__15733\,
            I => \N__15727\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__15730\,
            I => \N__15724\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__15727\,
            I => \N__15721\
        );

    \I__2990\ : CascadeBuf
    port map (
            O => \N__15724\,
            I => \N__15718\
        );

    \I__2989\ : CascadeBuf
    port map (
            O => \N__15721\,
            I => \N__15715\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__15718\,
            I => \N__15712\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__15715\,
            I => \N__15709\
        );

    \I__2986\ : CascadeBuf
    port map (
            O => \N__15712\,
            I => \N__15706\
        );

    \I__2985\ : CascadeBuf
    port map (
            O => \N__15709\,
            I => \N__15703\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__15706\,
            I => \N__15700\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__15703\,
            I => \N__15697\
        );

    \I__2982\ : CascadeBuf
    port map (
            O => \N__15700\,
            I => \N__15694\
        );

    \I__2981\ : CascadeBuf
    port map (
            O => \N__15697\,
            I => \N__15691\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__15694\,
            I => \N__15688\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__15691\,
            I => \N__15685\
        );

    \I__2978\ : CascadeBuf
    port map (
            O => \N__15688\,
            I => \N__15682\
        );

    \I__2977\ : CascadeBuf
    port map (
            O => \N__15685\,
            I => \N__15679\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__15682\,
            I => \N__15676\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__15679\,
            I => \N__15673\
        );

    \I__2974\ : CascadeBuf
    port map (
            O => \N__15676\,
            I => \N__15670\
        );

    \I__2973\ : CascadeBuf
    port map (
            O => \N__15673\,
            I => \N__15667\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__15670\,
            I => \N__15664\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__15667\,
            I => \N__15661\
        );

    \I__2970\ : CascadeBuf
    port map (
            O => \N__15664\,
            I => \N__15658\
        );

    \I__2969\ : CascadeBuf
    port map (
            O => \N__15661\,
            I => \N__15655\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__15658\,
            I => \N__15652\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__15655\,
            I => \N__15649\
        );

    \I__2966\ : CascadeBuf
    port map (
            O => \N__15652\,
            I => \N__15646\
        );

    \I__2965\ : CascadeBuf
    port map (
            O => \N__15649\,
            I => \N__15643\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__15646\,
            I => \N__15640\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__15643\,
            I => \N__15637\
        );

    \I__2962\ : CascadeBuf
    port map (
            O => \N__15640\,
            I => \N__15634\
        );

    \I__2961\ : CascadeBuf
    port map (
            O => \N__15637\,
            I => \N__15631\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__15634\,
            I => \N__15628\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__15631\,
            I => \N__15625\
        );

    \I__2958\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15622\
        );

    \I__2957\ : InMux
    port map (
            O => \N__15625\,
            I => \N__15619\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N__15616\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__15619\,
            I => \N__15613\
        );

    \I__2954\ : Span12Mux_s9_h
    port map (
            O => \N__15616\,
            I => \N__15610\
        );

    \I__2953\ : Span4Mux_h
    port map (
            O => \N__15613\,
            I => \N__15607\
        );

    \I__2952\ : Odrv12
    port map (
            O => \N__15610\,
            I => n27
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__15607\,
            I => n27
        );

    \I__2950\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15598\
        );

    \I__2949\ : IoInMux
    port map (
            O => \N__15601\,
            I => \N__15595\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__15598\,
            I => \N__15592\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__15595\,
            I => \N__15589\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__15592\,
            I => \N__15586\
        );

    \I__2945\ : Span12Mux_s11_h
    port map (
            O => \N__15589\,
            I => \N__15583\
        );

    \I__2944\ : Span4Mux_v
    port map (
            O => \N__15586\,
            I => \N__15580\
        );

    \I__2943\ : Odrv12
    port map (
            O => \N__15583\,
            I => \DEBUG_c_3_c\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__15580\,
            I => \DEBUG_c_3_c\
        );

    \I__2941\ : IoInMux
    port map (
            O => \N__15575\,
            I => \N__15572\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__15572\,
            I => \N__15569\
        );

    \I__2939\ : IoSpan4Mux
    port map (
            O => \N__15569\,
            I => \N__15566\
        );

    \I__2938\ : Span4Mux_s0_h
    port map (
            O => \N__15566\,
            I => \N__15562\
        );

    \I__2937\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15559\
        );

    \I__2936\ : Sp12to4
    port map (
            O => \N__15562\,
            I => \N__15556\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__15559\,
            I => \N__15553\
        );

    \I__2934\ : Span12Mux_s11_h
    port map (
            O => \N__15556\,
            I => \N__15550\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__15553\,
            I => \N__15547\
        );

    \I__2932\ : Span12Mux_v
    port map (
            O => \N__15550\,
            I => \N__15544\
        );

    \I__2931\ : Span4Mux_v
    port map (
            O => \N__15547\,
            I => \N__15541\
        );

    \I__2930\ : Odrv12
    port map (
            O => \N__15544\,
            I => \DEBUG_c_4_c\
        );

    \I__2929\ : Odrv4
    port map (
            O => \N__15541\,
            I => \DEBUG_c_4_c\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__15536\,
            I => \N__15533\
        );

    \I__2927\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15529\
        );

    \I__2926\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15524\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__15529\,
            I => \N__15521\
        );

    \I__2924\ : InMux
    port map (
            O => \N__15528\,
            I => \N__15518\
        );

    \I__2923\ : InMux
    port map (
            O => \N__15527\,
            I => \N__15515\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__15524\,
            I => \N__15510\
        );

    \I__2921\ : Span4Mux_v
    port map (
            O => \N__15521\,
            I => \N__15510\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__15518\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__15515\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__15510\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__2917\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15500\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__15500\,
            I => \transmit_module.video_signal_controller.n3628\
        );

    \I__2915\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15493\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__15496\,
            I => \N__15489\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__15493\,
            I => \N__15485\
        );

    \I__2912\ : InMux
    port map (
            O => \N__15492\,
            I => \N__15482\
        );

    \I__2911\ : InMux
    port map (
            O => \N__15489\,
            I => \N__15479\
        );

    \I__2910\ : InMux
    port map (
            O => \N__15488\,
            I => \N__15476\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__15485\,
            I => \N__15469\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__15482\,
            I => \N__15469\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__15479\,
            I => \N__15469\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__15476\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__15469\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__2904\ : InMux
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__15461\,
            I => \N__15457\
        );

    \I__2902\ : InMux
    port map (
            O => \N__15460\,
            I => \N__15454\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__15457\,
            I => \transmit_module.video_signal_controller.n3331\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__15454\,
            I => \transmit_module.video_signal_controller.n3331\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__15449\,
            I => \transmit_module.video_signal_controller.n7_adj_618_cascade_\
        );

    \I__2898\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__15443\,
            I => \N__15440\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__15440\,
            I => \transmit_module.video_signal_controller.n3622\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__15437\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_580_cascade_\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__15431\,
            I => \N__15426\
        );

    \I__2892\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15423\
        );

    \I__2891\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15420\
        );

    \I__2890\ : Span4Mux_v
    port map (
            O => \N__15426\,
            I => \N__15415\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__15423\,
            I => \N__15415\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__15420\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__15415\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__2886\ : InMux
    port map (
            O => \N__15410\,
            I => \N__15407\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__15407\,
            I => \N__15404\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__15404\,
            I => \transmit_module.video_signal_controller.n3477\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__15401\,
            I => \N__15398\
        );

    \I__2882\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15395\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__15395\,
            I => \N__15392\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__15392\,
            I => \transmit_module.video_signal_controller.n16\
        );

    \I__2879\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15386\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__15386\,
            I => \N__15382\
        );

    \I__2877\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15378\
        );

    \I__2876\ : Span4Mux_v
    port map (
            O => \N__15382\,
            I => \N__15374\
        );

    \I__2875\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15371\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__15378\,
            I => \N__15368\
        );

    \I__2873\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15365\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__15374\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__15371\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__2870\ : Odrv12
    port map (
            O => \N__15368\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__15365\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__2868\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__15353\,
            I => \N__15347\
        );

    \I__2866\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15342\
        );

    \I__2865\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15342\
        );

    \I__2864\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15339\
        );

    \I__2863\ : Span4Mux_h
    port map (
            O => \N__15347\,
            I => \N__15334\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__15342\,
            I => \N__15334\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__15339\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__15334\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__2859\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__15326\,
            I => \N__15323\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__15323\,
            I => \transmit_module.video_signal_controller.n3471\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__15320\,
            I => \N__15317\
        );

    \I__2855\ : InMux
    port map (
            O => \N__15317\,
            I => \N__15314\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__15314\,
            I => \N__15311\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__15311\,
            I => \transmit_module.video_signal_controller.n4_adj_617\
        );

    \I__2852\ : InMux
    port map (
            O => \N__15308\,
            I => \N__15305\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__15305\,
            I => \N__15301\
        );

    \I__2850\ : InMux
    port map (
            O => \N__15304\,
            I => \N__15296\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__15301\,
            I => \N__15293\
        );

    \I__2848\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15290\
        );

    \I__2847\ : InMux
    port map (
            O => \N__15299\,
            I => \N__15287\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__15296\,
            I => \N__15284\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__15293\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__15290\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__15287\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__15284\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__2841\ : InMux
    port map (
            O => \N__15275\,
            I => \N__15272\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__15272\,
            I => \N__15269\
        );

    \I__2839\ : Span4Mux_h
    port map (
            O => \N__15269\,
            I => \N__15265\
        );

    \I__2838\ : InMux
    port map (
            O => \N__15268\,
            I => \N__15262\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__15265\,
            I => \transmit_module.n144\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__15262\,
            I => \transmit_module.n144\
        );

    \I__2835\ : CEMux
    port map (
            O => \N__15257\,
            I => \N__15245\
        );

    \I__2834\ : CEMux
    port map (
            O => \N__15256\,
            I => \N__15241\
        );

    \I__2833\ : CEMux
    port map (
            O => \N__15255\,
            I => \N__15237\
        );

    \I__2832\ : CEMux
    port map (
            O => \N__15254\,
            I => \N__15234\
        );

    \I__2831\ : CEMux
    port map (
            O => \N__15253\,
            I => \N__15231\
        );

    \I__2830\ : CEMux
    port map (
            O => \N__15252\,
            I => \N__15228\
        );

    \I__2829\ : CEMux
    port map (
            O => \N__15251\,
            I => \N__15225\
        );

    \I__2828\ : CEMux
    port map (
            O => \N__15250\,
            I => \N__15222\
        );

    \I__2827\ : CEMux
    port map (
            O => \N__15249\,
            I => \N__15216\
        );

    \I__2826\ : CEMux
    port map (
            O => \N__15248\,
            I => \N__15213\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__15245\,
            I => \N__15209\
        );

    \I__2824\ : CEMux
    port map (
            O => \N__15244\,
            I => \N__15206\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__15241\,
            I => \N__15203\
        );

    \I__2822\ : CEMux
    port map (
            O => \N__15240\,
            I => \N__15200\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__15237\,
            I => \N__15196\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__15234\,
            I => \N__15191\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__15231\,
            I => \N__15191\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__15228\,
            I => \N__15188\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__15225\,
            I => \N__15183\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__15222\,
            I => \N__15183\
        );

    \I__2815\ : CEMux
    port map (
            O => \N__15221\,
            I => \N__15180\
        );

    \I__2814\ : CEMux
    port map (
            O => \N__15220\,
            I => \N__15177\
        );

    \I__2813\ : CEMux
    port map (
            O => \N__15219\,
            I => \N__15174\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__15216\,
            I => \N__15171\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__15213\,
            I => \N__15168\
        );

    \I__2810\ : CEMux
    port map (
            O => \N__15212\,
            I => \N__15165\
        );

    \I__2809\ : Span4Mux_v
    port map (
            O => \N__15209\,
            I => \N__15161\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__15206\,
            I => \N__15158\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__15203\,
            I => \N__15153\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__15200\,
            I => \N__15153\
        );

    \I__2805\ : CEMux
    port map (
            O => \N__15199\,
            I => \N__15150\
        );

    \I__2804\ : Span4Mux_v
    port map (
            O => \N__15196\,
            I => \N__15147\
        );

    \I__2803\ : Span4Mux_v
    port map (
            O => \N__15191\,
            I => \N__15142\
        );

    \I__2802\ : Span4Mux_v
    port map (
            O => \N__15188\,
            I => \N__15142\
        );

    \I__2801\ : Span4Mux_v
    port map (
            O => \N__15183\,
            I => \N__15135\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__15180\,
            I => \N__15135\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__15177\,
            I => \N__15135\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__15174\,
            I => \N__15132\
        );

    \I__2797\ : Span4Mux_h
    port map (
            O => \N__15171\,
            I => \N__15129\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__15168\,
            I => \N__15124\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__15165\,
            I => \N__15124\
        );

    \I__2794\ : CEMux
    port map (
            O => \N__15164\,
            I => \N__15121\
        );

    \I__2793\ : Span4Mux_h
    port map (
            O => \N__15161\,
            I => \N__15112\
        );

    \I__2792\ : Span4Mux_v
    port map (
            O => \N__15158\,
            I => \N__15112\
        );

    \I__2791\ : Span4Mux_v
    port map (
            O => \N__15153\,
            I => \N__15112\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__15150\,
            I => \N__15112\
        );

    \I__2789\ : Span4Mux_h
    port map (
            O => \N__15147\,
            I => \N__15103\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__15142\,
            I => \N__15103\
        );

    \I__2787\ : Span4Mux_h
    port map (
            O => \N__15135\,
            I => \N__15103\
        );

    \I__2786\ : Span4Mux_v
    port map (
            O => \N__15132\,
            I => \N__15103\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__15129\,
            I => \N__15098\
        );

    \I__2784\ : Span4Mux_h
    port map (
            O => \N__15124\,
            I => \N__15098\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__15121\,
            I => \N__15095\
        );

    \I__2782\ : Span4Mux_h
    port map (
            O => \N__15112\,
            I => \N__15092\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__15103\,
            I => \transmit_module.n3636\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__15098\,
            I => \transmit_module.n3636\
        );

    \I__2779\ : Odrv12
    port map (
            O => \N__15095\,
            I => \transmit_module.n3636\
        );

    \I__2778\ : Odrv4
    port map (
            O => \N__15092\,
            I => \transmit_module.n3636\
        );

    \I__2777\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15080\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__15077\,
            I => \transmit_module.video_signal_controller.n3412\
        );

    \I__2774\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15069\
        );

    \I__2773\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15066\
        );

    \I__2772\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15063\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__15069\,
            I => \N__15060\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__15066\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__15063\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__15060\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__2767\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15049\
        );

    \I__2766\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15045\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__15049\,
            I => \N__15042\
        );

    \I__2764\ : InMux
    port map (
            O => \N__15048\,
            I => \N__15039\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__15045\,
            I => \N__15036\
        );

    \I__2762\ : Span4Mux_h
    port map (
            O => \N__15042\,
            I => \N__15033\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__15039\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__15036\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__15033\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__2758\ : InMux
    port map (
            O => \N__15026\,
            I => \N__15023\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__15020\,
            I => \transmit_module.video_signal_controller.n3626\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__15017\,
            I => \N__15013\
        );

    \I__2754\ : InMux
    port map (
            O => \N__15016\,
            I => \N__15009\
        );

    \I__2753\ : InMux
    port map (
            O => \N__15013\,
            I => \N__15006\
        );

    \I__2752\ : InMux
    port map (
            O => \N__15012\,
            I => \N__15002\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__15009\,
            I => \N__14997\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__15006\,
            I => \N__14997\
        );

    \I__2749\ : InMux
    port map (
            O => \N__15005\,
            I => \N__14994\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__15002\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__14997\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__14994\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__14987\,
            I => \transmit_module.video_signal_controller.n3626_cascade_\
        );

    \I__2744\ : InMux
    port map (
            O => \N__14984\,
            I => \N__14979\
        );

    \I__2743\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14976\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14982\,
            I => \N__14973\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__14979\,
            I => \N__14970\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__14976\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__14973\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__14970\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__14963\,
            I => \transmit_module.n137_cascade_\
        );

    \I__2736\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14956\
        );

    \I__2735\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14951\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__14956\,
            I => \N__14948\
        );

    \I__2733\ : InMux
    port map (
            O => \N__14955\,
            I => \N__14945\
        );

    \I__2732\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14942\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__14951\,
            I => \N__14937\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__14948\,
            I => \N__14937\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__14945\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__14942\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__14937\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14926\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14923\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__14926\,
            I => \N__14917\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14917\
        );

    \I__2722\ : InMux
    port map (
            O => \N__14922\,
            I => \N__14913\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__14917\,
            I => \N__14910\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14907\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__14913\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__14910\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__14907\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__2716\ : InMux
    port map (
            O => \N__14900\,
            I => \N__14897\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__14897\,
            I => \N__14893\
        );

    \I__2714\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14888\
        );

    \I__2713\ : Span4Mux_v
    port map (
            O => \N__14893\,
            I => \N__14885\
        );

    \I__2712\ : InMux
    port map (
            O => \N__14892\,
            I => \N__14880\
        );

    \I__2711\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14880\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__14888\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__14885\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__14880\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14869\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14866\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__14869\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__14866\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__2703\ : InMux
    port map (
            O => \N__14861\,
            I => \N__14858\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__14858\,
            I => \N__14854\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__14857\,
            I => \N__14851\
        );

    \I__2700\ : Span4Mux_v
    port map (
            O => \N__14854\,
            I => \N__14848\
        );

    \I__2699\ : InMux
    port map (
            O => \N__14851\,
            I => \N__14845\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__14848\,
            I => \transmit_module.n113\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__14845\,
            I => \transmit_module.n113\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__14840\,
            I => \transmit_module.n142_cascade_\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__14837\,
            I => \N__14834\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14834\,
            I => \N__14831\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__14831\,
            I => \N__14828\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__14828\,
            I => \transmit_module.video_signal_controller.n45\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14822\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__14822\,
            I => \RX_TX_SYNC\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14816\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__14816\,
            I => \sync_buffer.BUFFER_0_0\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14813\,
            I => \N__14807\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14804\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14800\
        );

    \I__2684\ : InMux
    port map (
            O => \N__14810\,
            I => \N__14796\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14807\,
            I => \N__14791\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__14804\,
            I => \N__14788\
        );

    \I__2681\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14785\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__14800\,
            I => \N__14782\
        );

    \I__2679\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14779\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__14796\,
            I => \N__14775\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14772\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14794\,
            I => \N__14769\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__14791\,
            I => \N__14764\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__14788\,
            I => \N__14764\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__14785\,
            I => \N__14757\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__14782\,
            I => \N__14757\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__14779\,
            I => \N__14757\
        );

    \I__2670\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14754\
        );

    \I__2669\ : Span4Mux_h
    port map (
            O => \N__14775\,
            I => \N__14747\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__14772\,
            I => \N__14747\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__14769\,
            I => \N__14747\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__14764\,
            I => \RX_ADDR_12\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__14757\,
            I => \RX_ADDR_12\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__14754\,
            I => \RX_ADDR_12\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__14747\,
            I => \RX_ADDR_12\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__14738\,
            I => \N__14735\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14726\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__14734\,
            I => \N__14723\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__14733\,
            I => \N__14719\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__14732\,
            I => \N__14715\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__14731\,
            I => \N__14711\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__14730\,
            I => \N__14708\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__14729\,
            I => \N__14705\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14702\
        );

    \I__2653\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14687\
        );

    \I__2652\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14687\
        );

    \I__2651\ : InMux
    port map (
            O => \N__14719\,
            I => \N__14687\
        );

    \I__2650\ : InMux
    port map (
            O => \N__14718\,
            I => \N__14687\
        );

    \I__2649\ : InMux
    port map (
            O => \N__14715\,
            I => \N__14687\
        );

    \I__2648\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14687\
        );

    \I__2647\ : InMux
    port map (
            O => \N__14711\,
            I => \N__14687\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14684\
        );

    \I__2645\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14681\
        );

    \I__2644\ : Span4Mux_v
    port map (
            O => \N__14702\,
            I => \N__14676\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__14687\,
            I => \N__14676\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14670\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__14681\,
            I => \N__14670\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__14676\,
            I => \N__14665\
        );

    \I__2639\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14662\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__14670\,
            I => \N__14659\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__14669\,
            I => \N__14656\
        );

    \I__2636\ : InMux
    port map (
            O => \N__14668\,
            I => \N__14650\
        );

    \I__2635\ : Span4Mux_v
    port map (
            O => \N__14665\,
            I => \N__14644\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__14662\,
            I => \N__14644\
        );

    \I__2633\ : Sp12to4
    port map (
            O => \N__14659\,
            I => \N__14640\
        );

    \I__2632\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14637\
        );

    \I__2631\ : InMux
    port map (
            O => \N__14655\,
            I => \N__14634\
        );

    \I__2630\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14631\
        );

    \I__2629\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14628\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__14650\,
            I => \N__14625\
        );

    \I__2627\ : InMux
    port map (
            O => \N__14649\,
            I => \N__14622\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__14644\,
            I => \N__14617\
        );

    \I__2625\ : InMux
    port map (
            O => \N__14643\,
            I => \N__14614\
        );

    \I__2624\ : Span12Mux_v
    port map (
            O => \N__14640\,
            I => \N__14603\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__14637\,
            I => \N__14603\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__14634\,
            I => \N__14603\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__14631\,
            I => \N__14603\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__14628\,
            I => \N__14603\
        );

    \I__2619\ : Span4Mux_h
    port map (
            O => \N__14625\,
            I => \N__14600\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__14622\,
            I => \N__14597\
        );

    \I__2617\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14594\
        );

    \I__2616\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14591\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__14617\,
            I => \RX_WE\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__14614\,
            I => \RX_WE\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__14603\,
            I => \RX_WE\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__14600\,
            I => \RX_WE\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__14597\,
            I => \RX_WE\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__14594\,
            I => \RX_WE\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__14591\,
            I => \RX_WE\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__14576\,
            I => \N__14570\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__14575\,
            I => \N__14567\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__14574\,
            I => \N__14562\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__14573\,
            I => \N__14557\
        );

    \I__2604\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14554\
        );

    \I__2603\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14551\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__14566\,
            I => \N__14548\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__14565\,
            I => \N__14545\
        );

    \I__2600\ : InMux
    port map (
            O => \N__14562\,
            I => \N__14542\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__14561\,
            I => \N__14539\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__14560\,
            I => \N__14536\
        );

    \I__2597\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14533\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__14554\,
            I => \N__14529\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__14551\,
            I => \N__14526\
        );

    \I__2594\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14523\
        );

    \I__2593\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14520\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__14542\,
            I => \N__14517\
        );

    \I__2591\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14514\
        );

    \I__2590\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14511\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__14533\,
            I => \N__14508\
        );

    \I__2588\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14505\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__14529\,
            I => \N__14500\
        );

    \I__2586\ : Span4Mux_v
    port map (
            O => \N__14526\,
            I => \N__14500\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__14523\,
            I => \N__14493\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__14520\,
            I => \N__14493\
        );

    \I__2583\ : Span4Mux_v
    port map (
            O => \N__14517\,
            I => \N__14493\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__14514\,
            I => \N__14490\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__14511\,
            I => \N__14485\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__14508\,
            I => \N__14485\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__14505\,
            I => \RX_ADDR_13\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__14500\,
            I => \RX_ADDR_13\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__14493\,
            I => \RX_ADDR_13\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__14490\,
            I => \RX_ADDR_13\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__14485\,
            I => \RX_ADDR_13\
        );

    \I__2574\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14468\
        );

    \I__2573\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14464\
        );

    \I__2572\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14461\
        );

    \I__2571\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14457\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__14468\,
            I => \N__14452\
        );

    \I__2569\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14449\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__14464\,
            I => \N__14446\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__14461\,
            I => \N__14443\
        );

    \I__2566\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14440\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__14457\,
            I => \N__14437\
        );

    \I__2564\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14434\
        );

    \I__2563\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14431\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__14452\,
            I => \N__14423\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__14449\,
            I => \N__14423\
        );

    \I__2560\ : Span4Mux_h
    port map (
            O => \N__14446\,
            I => \N__14423\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__14443\,
            I => \N__14414\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__14440\,
            I => \N__14414\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__14437\,
            I => \N__14414\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__14434\,
            I => \N__14414\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__14431\,
            I => \N__14411\
        );

    \I__2554\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14408\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__14423\,
            I => \RX_ADDR_11\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__14414\,
            I => \RX_ADDR_11\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__14411\,
            I => \RX_ADDR_11\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__14408\,
            I => \RX_ADDR_11\
        );

    \I__2549\ : SRMux
    port map (
            O => \N__14399\,
            I => \N__14396\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__14396\,
            I => \N__14390\
        );

    \I__2547\ : SRMux
    port map (
            O => \N__14395\,
            I => \N__14387\
        );

    \I__2546\ : SRMux
    port map (
            O => \N__14394\,
            I => \N__14384\
        );

    \I__2545\ : SRMux
    port map (
            O => \N__14393\,
            I => \N__14381\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__14390\,
            I => \N__14376\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__14387\,
            I => \N__14376\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__14384\,
            I => \N__14371\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__14381\,
            I => \N__14371\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__14376\,
            I => \N__14366\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__14371\,
            I => \N__14366\
        );

    \I__2538\ : Sp12to4
    port map (
            O => \N__14366\,
            I => \N__14363\
        );

    \I__2537\ : Odrv12
    port map (
            O => \N__14363\,
            I => \line_buffer.n532\
        );

    \I__2536\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14357\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14354\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__14354\,
            I => \N__14351\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__14351\,
            I => \tvp_video_buffer.BUFFER_1_3\
        );

    \I__2532\ : InMux
    port map (
            O => \N__14348\,
            I => \N__14343\
        );

    \I__2531\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14340\
        );

    \I__2530\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14336\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__14343\,
            I => \N__14331\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__14340\,
            I => \N__14328\
        );

    \I__2527\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14324\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__14336\,
            I => \N__14321\
        );

    \I__2525\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14318\
        );

    \I__2524\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14315\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__14331\,
            I => \N__14312\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__14328\,
            I => \N__14309\
        );

    \I__2521\ : InMux
    port map (
            O => \N__14327\,
            I => \N__14306\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__14324\,
            I => \N__14302\
        );

    \I__2519\ : Span12Mux_s9_v
    port map (
            O => \N__14321\,
            I => \N__14295\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__14318\,
            I => \N__14295\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__14315\,
            I => \N__14295\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__14312\,
            I => \N__14290\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__14309\,
            I => \N__14290\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__14306\,
            I => \N__14287\
        );

    \I__2513\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14284\
        );

    \I__2512\ : Span12Mux_s10_v
    port map (
            O => \N__14302\,
            I => \N__14279\
        );

    \I__2511\ : Span12Mux_v
    port map (
            O => \N__14295\,
            I => \N__14279\
        );

    \I__2510\ : Sp12to4
    port map (
            O => \N__14290\,
            I => \N__14272\
        );

    \I__2509\ : Span12Mux_h
    port map (
            O => \N__14287\,
            I => \N__14272\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14272\
        );

    \I__2507\ : Odrv12
    port map (
            O => \N__14279\,
            I => \RX_DATA_1\
        );

    \I__2506\ : Odrv12
    port map (
            O => \N__14272\,
            I => \RX_DATA_1\
        );

    \I__2505\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14264\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__14264\,
            I => \N__14261\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__14261\,
            I => \sync_buffer.BUFFER_1_0\
        );

    \I__2502\ : InMux
    port map (
            O => \N__14258\,
            I => \N__14255\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__14255\,
            I => \RX_TX_SYNC_BUFF\
        );

    \I__2500\ : SRMux
    port map (
            O => \N__14252\,
            I => \N__14249\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__14249\,
            I => \N__14243\
        );

    \I__2498\ : SRMux
    port map (
            O => \N__14248\,
            I => \N__14240\
        );

    \I__2497\ : CEMux
    port map (
            O => \N__14247\,
            I => \N__14236\
        );

    \I__2496\ : CEMux
    port map (
            O => \N__14246\,
            I => \N__14233\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__14243\,
            I => \N__14228\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__14240\,
            I => \N__14228\
        );

    \I__2493\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14225\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__14236\,
            I => \N__14222\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__14233\,
            I => \N__14217\
        );

    \I__2490\ : Span4Mux_h
    port map (
            O => \N__14228\,
            I => \N__14217\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__14225\,
            I => \N__14214\
        );

    \I__2488\ : Odrv12
    port map (
            O => \N__14222\,
            I => \transmit_module.video_signal_controller.n2036\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__14217\,
            I => \transmit_module.video_signal_controller.n2036\
        );

    \I__2486\ : Odrv4
    port map (
            O => \N__14214\,
            I => \transmit_module.video_signal_controller.n2036\
        );

    \I__2485\ : SRMux
    port map (
            O => \N__14207\,
            I => \N__14204\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__14204\,
            I => \N__14200\
        );

    \I__2483\ : SRMux
    port map (
            O => \N__14203\,
            I => \N__14197\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__14200\,
            I => \N__14194\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__14197\,
            I => \N__14191\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__14194\,
            I => \transmit_module.video_signal_controller.n2378\
        );

    \I__2479\ : Odrv12
    port map (
            O => \N__14191\,
            I => \transmit_module.video_signal_controller.n2378\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__14186\,
            I => \transmit_module.video_signal_controller.n49_cascade_\
        );

    \I__2477\ : SRMux
    port map (
            O => \N__14183\,
            I => \N__14179\
        );

    \I__2476\ : SRMux
    port map (
            O => \N__14182\,
            I => \N__14176\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__14179\,
            I => \N__14169\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__14176\,
            I => \N__14169\
        );

    \I__2473\ : SRMux
    port map (
            O => \N__14175\,
            I => \N__14166\
        );

    \I__2472\ : SRMux
    port map (
            O => \N__14174\,
            I => \N__14163\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__14169\,
            I => \N__14156\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__14166\,
            I => \N__14156\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__14163\,
            I => \N__14156\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__14156\,
            I => \N__14153\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__14153\,
            I => \N__14150\
        );

    \I__2466\ : Span4Mux_h
    port map (
            O => \N__14150\,
            I => \N__14147\
        );

    \I__2465\ : Span4Mux_h
    port map (
            O => \N__14147\,
            I => \N__14144\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__14144\,
            I => \line_buffer.n468\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__2462\ : CascadeBuf
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__14135\,
            I => \N__14132\
        );

    \I__2460\ : CascadeBuf
    port map (
            O => \N__14132\,
            I => \N__14128\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__14131\,
            I => \N__14125\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__14128\,
            I => \N__14122\
        );

    \I__2457\ : CascadeBuf
    port map (
            O => \N__14125\,
            I => \N__14119\
        );

    \I__2456\ : CascadeBuf
    port map (
            O => \N__14122\,
            I => \N__14116\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__14119\,
            I => \N__14113\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__14116\,
            I => \N__14110\
        );

    \I__2453\ : CascadeBuf
    port map (
            O => \N__14113\,
            I => \N__14107\
        );

    \I__2452\ : CascadeBuf
    port map (
            O => \N__14110\,
            I => \N__14104\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__14107\,
            I => \N__14101\
        );

    \I__2450\ : CascadeMux
    port map (
            O => \N__14104\,
            I => \N__14098\
        );

    \I__2449\ : CascadeBuf
    port map (
            O => \N__14101\,
            I => \N__14095\
        );

    \I__2448\ : CascadeBuf
    port map (
            O => \N__14098\,
            I => \N__14092\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__14095\,
            I => \N__14089\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__14092\,
            I => \N__14086\
        );

    \I__2445\ : CascadeBuf
    port map (
            O => \N__14089\,
            I => \N__14083\
        );

    \I__2444\ : CascadeBuf
    port map (
            O => \N__14086\,
            I => \N__14080\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__14083\,
            I => \N__14077\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__14080\,
            I => \N__14074\
        );

    \I__2441\ : CascadeBuf
    port map (
            O => \N__14077\,
            I => \N__14071\
        );

    \I__2440\ : CascadeBuf
    port map (
            O => \N__14074\,
            I => \N__14068\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__14071\,
            I => \N__14065\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__14068\,
            I => \N__14062\
        );

    \I__2437\ : CascadeBuf
    port map (
            O => \N__14065\,
            I => \N__14059\
        );

    \I__2436\ : CascadeBuf
    port map (
            O => \N__14062\,
            I => \N__14056\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__14059\,
            I => \N__14053\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__14056\,
            I => \N__14050\
        );

    \I__2433\ : CascadeBuf
    port map (
            O => \N__14053\,
            I => \N__14047\
        );

    \I__2432\ : CascadeBuf
    port map (
            O => \N__14050\,
            I => \N__14044\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__14047\,
            I => \N__14041\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__14044\,
            I => \N__14038\
        );

    \I__2429\ : CascadeBuf
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__2428\ : CascadeBuf
    port map (
            O => \N__14038\,
            I => \N__14032\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__14035\,
            I => \N__14029\
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__14032\,
            I => \N__14026\
        );

    \I__2425\ : CascadeBuf
    port map (
            O => \N__14029\,
            I => \N__14023\
        );

    \I__2424\ : CascadeBuf
    port map (
            O => \N__14026\,
            I => \N__14020\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__14023\,
            I => \N__14017\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__14020\,
            I => \N__14014\
        );

    \I__2421\ : CascadeBuf
    port map (
            O => \N__14017\,
            I => \N__14011\
        );

    \I__2420\ : CascadeBuf
    port map (
            O => \N__14014\,
            I => \N__14008\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__14011\,
            I => \N__14005\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__14008\,
            I => \N__14002\
        );

    \I__2417\ : CascadeBuf
    port map (
            O => \N__14005\,
            I => \N__13999\
        );

    \I__2416\ : CascadeBuf
    port map (
            O => \N__14002\,
            I => \N__13996\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__13999\,
            I => \N__13993\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__13996\,
            I => \N__13990\
        );

    \I__2413\ : CascadeBuf
    port map (
            O => \N__13993\,
            I => \N__13987\
        );

    \I__2412\ : CascadeBuf
    port map (
            O => \N__13990\,
            I => \N__13984\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__13987\,
            I => \N__13981\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__13984\,
            I => \N__13978\
        );

    \I__2409\ : CascadeBuf
    port map (
            O => \N__13981\,
            I => \N__13975\
        );

    \I__2408\ : CascadeBuf
    port map (
            O => \N__13978\,
            I => \N__13972\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__13975\,
            I => \N__13969\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__13972\,
            I => \N__13966\
        );

    \I__2405\ : CascadeBuf
    port map (
            O => \N__13969\,
            I => \N__13963\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13966\,
            I => \N__13960\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__13963\,
            I => \N__13957\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__13960\,
            I => \N__13954\
        );

    \I__2401\ : CascadeBuf
    port map (
            O => \N__13957\,
            I => \N__13951\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__13954\,
            I => \N__13948\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__13951\,
            I => \N__13945\
        );

    \I__2398\ : Span4Mux_v
    port map (
            O => \N__13948\,
            I => \N__13942\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13945\,
            I => \N__13939\
        );

    \I__2396\ : Span4Mux_h
    port map (
            O => \N__13942\,
            I => \N__13936\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__13939\,
            I => \N__13933\
        );

    \I__2394\ : Span4Mux_h
    port map (
            O => \N__13936\,
            I => \N__13930\
        );

    \I__2393\ : Span4Mux_v
    port map (
            O => \N__13933\,
            I => \N__13927\
        );

    \I__2392\ : Span4Mux_h
    port map (
            O => \N__13930\,
            I => \N__13922\
        );

    \I__2391\ : Span4Mux_h
    port map (
            O => \N__13927\,
            I => \N__13922\
        );

    \I__2390\ : Sp12to4
    port map (
            O => \N__13922\,
            I => \N__13919\
        );

    \I__2389\ : Odrv12
    port map (
            O => \N__13919\,
            I => n25
        );

    \I__2388\ : InMux
    port map (
            O => \N__13916\,
            I => \N__13913\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__13913\,
            I => \transmit_module.ADDR_Y_COMPONENT_3\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__13907\,
            I => \N__13904\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__13901\,
            I => \tvp_video_buffer.BUFFER_0_4\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13892\,
            I => \N__13886\
        );

    \I__2379\ : InMux
    port map (
            O => \N__13891\,
            I => \N__13883\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13890\,
            I => \N__13880\
        );

    \I__2377\ : InMux
    port map (
            O => \N__13889\,
            I => \N__13877\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__13886\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__13883\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__13880\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13877\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13864\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13859\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__13864\,
            I => \N__13856\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13853\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13850\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__13859\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__13856\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13853\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__13850\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__13841\,
            I => \N__13835\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13840\,
            I => \N__13832\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13829\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13838\,
            I => \N__13826\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13823\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13832\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__13829\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__13826\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__13823\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__2354\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13808\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13805\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13800\
        );

    \I__2351\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13800\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__13808\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__13805\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__13800\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__13793\,
            I => \N__13790\
        );

    \I__2346\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13784\
        );

    \I__2345\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13781\
        );

    \I__2344\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13776\
        );

    \I__2343\ : InMux
    port map (
            O => \N__13787\,
            I => \N__13776\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__13784\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13781\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__13776\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__13769\,
            I => \N__13765\
        );

    \I__2338\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13758\
        );

    \I__2337\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13758\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13755\
        );

    \I__2335\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13752\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__13758\,
            I => \N__13747\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__13755\,
            I => \N__13747\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13752\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__13747\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13742\,
            I => \N__13739\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13739\,
            I => \receive_module.rx_counter.n10_adj_610\
        );

    \I__2328\ : InMux
    port map (
            O => \N__13736\,
            I => \N__13728\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13735\,
            I => \N__13728\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13734\,
            I => \N__13725\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13722\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__13728\,
            I => \N__13719\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__13725\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13722\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__13719\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__13712\,
            I => \receive_module.rx_counter.n14_cascade_\
        );

    \I__2319\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13705\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13708\,
            I => \N__13702\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13705\,
            I => \receive_module.rx_counter.n3633\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__13702\,
            I => \receive_module.rx_counter.n3633\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__13697\,
            I => \transmit_module.video_signal_controller.n2947_cascade_\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__13694\,
            I => \N__13691\
        );

    \I__2313\ : InMux
    port map (
            O => \N__13691\,
            I => \N__13688\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__13688\,
            I => \N__13685\
        );

    \I__2311\ : Span12Mux_v
    port map (
            O => \N__13685\,
            I => \N__13682\
        );

    \I__2310\ : Span12Mux_h
    port map (
            O => \N__13682\,
            I => \N__13679\
        );

    \I__2309\ : Odrv12
    port map (
            O => \N__13679\,
            I => \line_buffer.n522\
        );

    \I__2308\ : InMux
    port map (
            O => \N__13676\,
            I => \N__13673\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__13673\,
            I => \N__13670\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__13670\,
            I => \N__13667\
        );

    \I__2305\ : Span4Mux_h
    port map (
            O => \N__13667\,
            I => \N__13664\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__13664\,
            I => \line_buffer.n530\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__13661\,
            I => \N__13658\
        );

    \I__2302\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13652\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13649\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13646\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13643\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__13652\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__13649\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__13646\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__13643\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13628\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13633\,
            I => \N__13625\
        );

    \I__2292\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13622\
        );

    \I__2291\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13619\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__13628\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__13625\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__13622\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__13619\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__2286\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13607\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__13607\,
            I => \transmit_module.video_signal_controller.n18\
        );

    \I__2284\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13599\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__13603\,
            I => \N__13596\
        );

    \I__2282\ : InMux
    port map (
            O => \N__13602\,
            I => \N__13592\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__13599\,
            I => \N__13589\
        );

    \I__2280\ : InMux
    port map (
            O => \N__13596\,
            I => \N__13584\
        );

    \I__2279\ : InMux
    port map (
            O => \N__13595\,
            I => \N__13584\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__13592\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__13589\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__13584\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__2275\ : InMux
    port map (
            O => \N__13577\,
            I => \N__13574\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__13574\,
            I => \N__13569\
        );

    \I__2273\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13565\
        );

    \I__2272\ : InMux
    port map (
            O => \N__13572\,
            I => \N__13562\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__13569\,
            I => \N__13559\
        );

    \I__2270\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13556\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__13565\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__13562\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__13559\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__13556\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__2265\ : InMux
    port map (
            O => \N__13547\,
            I => \N__13544\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__13544\,
            I => \transmit_module.video_signal_controller.n4\
        );

    \I__2263\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13535\
        );

    \I__2262\ : InMux
    port map (
            O => \N__13540\,
            I => \N__13532\
        );

    \I__2261\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13529\
        );

    \I__2260\ : InMux
    port map (
            O => \N__13538\,
            I => \N__13526\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__13535\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__13532\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__13529\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__13526\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__13517\,
            I => \transmit_module.video_signal_controller.n3625_cascade_\
        );

    \I__2254\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13508\
        );

    \I__2253\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13503\
        );

    \I__2252\ : InMux
    port map (
            O => \N__13512\,
            I => \N__13503\
        );

    \I__2251\ : InMux
    port map (
            O => \N__13511\,
            I => \N__13500\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__13508\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__13503\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__13500\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__2247\ : SRMux
    port map (
            O => \N__13493\,
            I => \N__13490\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__13487\,
            I => \N__13481\
        );

    \I__2244\ : SRMux
    port map (
            O => \N__13486\,
            I => \N__13478\
        );

    \I__2243\ : SRMux
    port map (
            O => \N__13485\,
            I => \N__13475\
        );

    \I__2242\ : SRMux
    port map (
            O => \N__13484\,
            I => \N__13472\
        );

    \I__2241\ : Span4Mux_v
    port map (
            O => \N__13481\,
            I => \N__13467\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__13478\,
            I => \N__13467\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__13475\,
            I => \N__13464\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__13472\,
            I => \N__13461\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__13467\,
            I => \N__13456\
        );

    \I__2236\ : Span4Mux_h
    port map (
            O => \N__13464\,
            I => \N__13456\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__13461\,
            I => \N__13453\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__13456\,
            I => \N__13448\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__13453\,
            I => \N__13448\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__13448\,
            I => \line_buffer.n597\
        );

    \I__2231\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__13442\,
            I => \N__13439\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2228\ : Span4Mux_v
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2227\ : Span4Mux_h
    port map (
            O => \N__13433\,
            I => \N__13430\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__13430\,
            I => \line_buffer.n594\
        );

    \I__2225\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13424\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__13424\,
            I => \N__13421\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__13421\,
            I => \N__13418\
        );

    \I__2222\ : Span4Mux_h
    port map (
            O => \N__13418\,
            I => \N__13415\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__13415\,
            I => \line_buffer.n586\
        );

    \I__2220\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13409\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__13409\,
            I => \line_buffer.n3591\
        );

    \I__2218\ : InMux
    port map (
            O => \N__13406\,
            I => \transmit_module.video_signal_controller.n3145\
        );

    \I__2217\ : InMux
    port map (
            O => \N__13403\,
            I => \transmit_module.video_signal_controller.n3146\
        );

    \I__2216\ : SRMux
    port map (
            O => \N__13400\,
            I => \N__13396\
        );

    \I__2215\ : SRMux
    port map (
            O => \N__13399\,
            I => \N__13393\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__13396\,
            I => \N__13389\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__13393\,
            I => \N__13386\
        );

    \I__2212\ : SRMux
    port map (
            O => \N__13392\,
            I => \N__13383\
        );

    \I__2211\ : Span4Mux_v
    port map (
            O => \N__13389\,
            I => \N__13380\
        );

    \I__2210\ : Span4Mux_h
    port map (
            O => \N__13386\,
            I => \N__13375\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__13383\,
            I => \N__13375\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__13380\,
            I => \N__13371\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__13375\,
            I => \N__13368\
        );

    \I__2206\ : SRMux
    port map (
            O => \N__13374\,
            I => \N__13365\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__13371\,
            I => \N__13358\
        );

    \I__2204\ : Span4Mux_h
    port map (
            O => \N__13368\,
            I => \N__13358\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__13365\,
            I => \N__13358\
        );

    \I__2202\ : Span4Mux_h
    port map (
            O => \N__13358\,
            I => \N__13355\
        );

    \I__2201\ : Sp12to4
    port map (
            O => \N__13355\,
            I => \N__13352\
        );

    \I__2200\ : Odrv12
    port map (
            O => \N__13352\,
            I => \line_buffer.n564\
        );

    \I__2199\ : InMux
    port map (
            O => \N__13349\,
            I => \N__13346\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__13346\,
            I => \transmit_module.video_signal_controller.n3624\
        );

    \I__2197\ : InMux
    port map (
            O => \N__13343\,
            I => \N__13337\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__13342\,
            I => \N__13334\
        );

    \I__2195\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13331\
        );

    \I__2194\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13328\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__13337\,
            I => \N__13325\
        );

    \I__2192\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13322\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__13331\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__13328\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__13325\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__13322\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__2187\ : InMux
    port map (
            O => \N__13313\,
            I => \N__13307\
        );

    \I__2186\ : InMux
    port map (
            O => \N__13312\,
            I => \N__13304\
        );

    \I__2185\ : InMux
    port map (
            O => \N__13311\,
            I => \N__13299\
        );

    \I__2184\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13299\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__13307\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__13304\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__13299\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__2180\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13287\
        );

    \I__2179\ : InMux
    port map (
            O => \N__13291\,
            I => \N__13284\
        );

    \I__2178\ : InMux
    port map (
            O => \N__13290\,
            I => \N__13281\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__13287\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__13284\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__13281\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__13274\,
            I => \N__13271\
        );

    \I__2173\ : InMux
    port map (
            O => \N__13271\,
            I => \N__13265\
        );

    \I__2172\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13265\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__13265\,
            I => \N__13262\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__13262\,
            I => \transmit_module.video_signal_controller.n2001\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__13259\,
            I => \transmit_module.video_signal_controller.n2917_cascade_\
        );

    \I__2168\ : InMux
    port map (
            O => \N__13256\,
            I => \N__13250\
        );

    \I__2167\ : InMux
    port map (
            O => \N__13255\,
            I => \N__13250\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__13250\,
            I => \transmit_module.video_signal_controller.n3313\
        );

    \I__2165\ : InMux
    port map (
            O => \N__13247\,
            I => \transmit_module.video_signal_controller.n3136\
        );

    \I__2164\ : InMux
    port map (
            O => \N__13244\,
            I => \transmit_module.video_signal_controller.n3137\
        );

    \I__2163\ : InMux
    port map (
            O => \N__13241\,
            I => \transmit_module.video_signal_controller.n3138\
        );

    \I__2162\ : InMux
    port map (
            O => \N__13238\,
            I => \transmit_module.video_signal_controller.n3139\
        );

    \I__2161\ : InMux
    port map (
            O => \N__13235\,
            I => \transmit_module.video_signal_controller.n3140\
        );

    \I__2160\ : InMux
    port map (
            O => \N__13232\,
            I => \transmit_module.video_signal_controller.n3141\
        );

    \I__2159\ : InMux
    port map (
            O => \N__13229\,
            I => \transmit_module.video_signal_controller.n3142\
        );

    \I__2158\ : InMux
    port map (
            O => \N__13226\,
            I => \bfn_13_13_0_\
        );

    \I__2157\ : InMux
    port map (
            O => \N__13223\,
            I => \transmit_module.video_signal_controller.n3144\
        );

    \I__2156\ : InMux
    port map (
            O => \N__13220\,
            I => \receive_module.rx_counter.n3118\
        );

    \I__2155\ : InMux
    port map (
            O => \N__13217\,
            I => \receive_module.rx_counter.n3119\
        );

    \I__2154\ : InMux
    port map (
            O => \N__13214\,
            I => \receive_module.rx_counter.n3120\
        );

    \I__2153\ : InMux
    port map (
            O => \N__13211\,
            I => \N__13206\
        );

    \I__2152\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13201\
        );

    \I__2151\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13201\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__13206\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__13201\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__2148\ : InMux
    port map (
            O => \N__13196\,
            I => \receive_module.rx_counter.n3121\
        );

    \I__2147\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13188\
        );

    \I__2146\ : InMux
    port map (
            O => \N__13192\,
            I => \N__13185\
        );

    \I__2145\ : InMux
    port map (
            O => \N__13191\,
            I => \N__13182\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__13188\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__13185\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__13182\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__2141\ : InMux
    port map (
            O => \N__13175\,
            I => \receive_module.rx_counter.n3122\
        );

    \I__2140\ : InMux
    port map (
            O => \N__13172\,
            I => \receive_module.rx_counter.n3123\
        );

    \I__2139\ : InMux
    port map (
            O => \N__13169\,
            I => \bfn_13_10_0_\
        );

    \I__2138\ : CEMux
    port map (
            O => \N__13166\,
            I => \N__13162\
        );

    \I__2137\ : CEMux
    port map (
            O => \N__13165\,
            I => \N__13159\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__13162\,
            I => \N__13156\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__13159\,
            I => \N__13153\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__13156\,
            I => \receive_module.rx_counter.n2063\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__13153\,
            I => \receive_module.rx_counter.n2063\
        );

    \I__2132\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13145\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__13145\,
            I => \receive_module.n134\
        );

    \I__2130\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13138\
        );

    \I__2129\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13135\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__13138\,
            I => \N__13130\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__13135\,
            I => \N__13130\
        );

    \I__2126\ : Span4Mux_v
    port map (
            O => \N__13130\,
            I => \N__13126\
        );

    \I__2125\ : InMux
    port map (
            O => \N__13129\,
            I => \N__13123\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__13126\,
            I => \N__13111\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__13123\,
            I => \N__13111\
        );

    \I__2122\ : InMux
    port map (
            O => \N__13122\,
            I => \N__13096\
        );

    \I__2121\ : InMux
    port map (
            O => \N__13121\,
            I => \N__13096\
        );

    \I__2120\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13096\
        );

    \I__2119\ : InMux
    port map (
            O => \N__13119\,
            I => \N__13096\
        );

    \I__2118\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13096\
        );

    \I__2117\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13096\
        );

    \I__2116\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13096\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__13111\,
            I => \N__13090\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__13096\,
            I => \N__13090\
        );

    \I__2113\ : InMux
    port map (
            O => \N__13095\,
            I => \N__13083\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__13090\,
            I => \N__13080\
        );

    \I__2111\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13077\
        );

    \I__2110\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13074\
        );

    \I__2109\ : InMux
    port map (
            O => \N__13087\,
            I => \N__13069\
        );

    \I__2108\ : InMux
    port map (
            O => \N__13086\,
            I => \N__13069\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__13083\,
            I => \N__13064\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__13080\,
            I => \N__13059\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__13077\,
            I => \N__13059\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__13074\,
            I => \N__13054\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__13069\,
            I => \N__13054\
        );

    \I__2102\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13049\
        );

    \I__2101\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13049\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__13064\,
            I => \TVP_VSYNC_buff\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__13059\,
            I => \TVP_VSYNC_buff\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__13054\,
            I => \TVP_VSYNC_buff\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__13049\,
            I => \TVP_VSYNC_buff\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__13040\,
            I => \N__13037\
        );

    \I__2095\ : CascadeBuf
    port map (
            O => \N__13037\,
            I => \N__13033\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__13036\,
            I => \N__13030\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__13033\,
            I => \N__13027\
        );

    \I__2092\ : CascadeBuf
    port map (
            O => \N__13030\,
            I => \N__13024\
        );

    \I__2091\ : CascadeBuf
    port map (
            O => \N__13027\,
            I => \N__13021\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__13024\,
            I => \N__13018\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__13021\,
            I => \N__13015\
        );

    \I__2088\ : CascadeBuf
    port map (
            O => \N__13018\,
            I => \N__13012\
        );

    \I__2087\ : CascadeBuf
    port map (
            O => \N__13015\,
            I => \N__13009\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__13012\,
            I => \N__13006\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__13009\,
            I => \N__13003\
        );

    \I__2084\ : CascadeBuf
    port map (
            O => \N__13006\,
            I => \N__13000\
        );

    \I__2083\ : CascadeBuf
    port map (
            O => \N__13003\,
            I => \N__12997\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__13000\,
            I => \N__12994\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__12997\,
            I => \N__12991\
        );

    \I__2080\ : CascadeBuf
    port map (
            O => \N__12994\,
            I => \N__12988\
        );

    \I__2079\ : CascadeBuf
    port map (
            O => \N__12991\,
            I => \N__12985\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__12988\,
            I => \N__12982\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__12985\,
            I => \N__12979\
        );

    \I__2076\ : CascadeBuf
    port map (
            O => \N__12982\,
            I => \N__12976\
        );

    \I__2075\ : CascadeBuf
    port map (
            O => \N__12979\,
            I => \N__12973\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__12976\,
            I => \N__12970\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__12973\,
            I => \N__12967\
        );

    \I__2072\ : CascadeBuf
    port map (
            O => \N__12970\,
            I => \N__12964\
        );

    \I__2071\ : CascadeBuf
    port map (
            O => \N__12967\,
            I => \N__12961\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__12964\,
            I => \N__12958\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__12961\,
            I => \N__12955\
        );

    \I__2068\ : CascadeBuf
    port map (
            O => \N__12958\,
            I => \N__12952\
        );

    \I__2067\ : CascadeBuf
    port map (
            O => \N__12955\,
            I => \N__12949\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__12952\,
            I => \N__12946\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__12949\,
            I => \N__12943\
        );

    \I__2064\ : CascadeBuf
    port map (
            O => \N__12946\,
            I => \N__12940\
        );

    \I__2063\ : CascadeBuf
    port map (
            O => \N__12943\,
            I => \N__12937\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__12940\,
            I => \N__12934\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__12937\,
            I => \N__12931\
        );

    \I__2060\ : CascadeBuf
    port map (
            O => \N__12934\,
            I => \N__12928\
        );

    \I__2059\ : CascadeBuf
    port map (
            O => \N__12931\,
            I => \N__12925\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__12928\,
            I => \N__12922\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__12925\,
            I => \N__12919\
        );

    \I__2056\ : CascadeBuf
    port map (
            O => \N__12922\,
            I => \N__12916\
        );

    \I__2055\ : CascadeBuf
    port map (
            O => \N__12919\,
            I => \N__12913\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__12916\,
            I => \N__12910\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__12913\,
            I => \N__12907\
        );

    \I__2052\ : CascadeBuf
    port map (
            O => \N__12910\,
            I => \N__12904\
        );

    \I__2051\ : CascadeBuf
    port map (
            O => \N__12907\,
            I => \N__12901\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__12904\,
            I => \N__12898\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__12901\,
            I => \N__12895\
        );

    \I__2048\ : CascadeBuf
    port map (
            O => \N__12898\,
            I => \N__12892\
        );

    \I__2047\ : CascadeBuf
    port map (
            O => \N__12895\,
            I => \N__12889\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__12892\,
            I => \N__12886\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__12889\,
            I => \N__12883\
        );

    \I__2044\ : CascadeBuf
    port map (
            O => \N__12886\,
            I => \N__12880\
        );

    \I__2043\ : CascadeBuf
    port map (
            O => \N__12883\,
            I => \N__12877\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__12880\,
            I => \N__12874\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__12877\,
            I => \N__12871\
        );

    \I__2040\ : CascadeBuf
    port map (
            O => \N__12874\,
            I => \N__12868\
        );

    \I__2039\ : CascadeBuf
    port map (
            O => \N__12871\,
            I => \N__12865\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__12868\,
            I => \N__12862\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__12865\,
            I => \N__12859\
        );

    \I__2036\ : CascadeBuf
    port map (
            O => \N__12862\,
            I => \N__12856\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12859\,
            I => \N__12853\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__12856\,
            I => \N__12850\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__12853\,
            I => \N__12847\
        );

    \I__2032\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12844\
        );

    \I__2031\ : Span4Mux_s1_v
    port map (
            O => \N__12847\,
            I => \N__12841\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__12844\,
            I => \N__12838\
        );

    \I__2029\ : Span4Mux_h
    port map (
            O => \N__12841\,
            I => \N__12835\
        );

    \I__2028\ : Span12Mux_s1_v
    port map (
            O => \N__12838\,
            I => \N__12832\
        );

    \I__2027\ : Sp12to4
    port map (
            O => \N__12835\,
            I => \N__12825\
        );

    \I__2026\ : Span12Mux_h
    port map (
            O => \N__12832\,
            I => \N__12825\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12831\,
            I => \N__12822\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12830\,
            I => \N__12819\
        );

    \I__2023\ : Span12Mux_v
    port map (
            O => \N__12825\,
            I => \N__12816\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__12822\,
            I => \RX_ADDR_2\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__12819\,
            I => \RX_ADDR_2\
        );

    \I__2020\ : Odrv12
    port map (
            O => \N__12816\,
            I => \RX_ADDR_2\
        );

    \I__2019\ : SRMux
    port map (
            O => \N__12809\,
            I => \N__12805\
        );

    \I__2018\ : SRMux
    port map (
            O => \N__12808\,
            I => \N__12802\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__12805\,
            I => \N__12799\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12802\,
            I => \N__12796\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__12799\,
            I => \N__12790\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__12796\,
            I => \N__12790\
        );

    \I__2013\ : SRMux
    port map (
            O => \N__12795\,
            I => \N__12787\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__12790\,
            I => \N__12781\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__12787\,
            I => \N__12781\
        );

    \I__2010\ : SRMux
    port map (
            O => \N__12786\,
            I => \N__12778\
        );

    \I__2009\ : Span4Mux_v
    port map (
            O => \N__12781\,
            I => \N__12773\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__12778\,
            I => \N__12773\
        );

    \I__2007\ : Span4Mux_v
    port map (
            O => \N__12773\,
            I => \N__12768\
        );

    \I__2006\ : SRMux
    port map (
            O => \N__12772\,
            I => \N__12765\
        );

    \I__2005\ : SRMux
    port map (
            O => \N__12771\,
            I => \N__12762\
        );

    \I__2004\ : Span4Mux_v
    port map (
            O => \N__12768\,
            I => \N__12755\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__12765\,
            I => \N__12755\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12762\,
            I => \N__12752\
        );

    \I__2001\ : SRMux
    port map (
            O => \N__12761\,
            I => \N__12749\
        );

    \I__2000\ : SRMux
    port map (
            O => \N__12760\,
            I => \N__12746\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__12755\,
            I => \N__12743\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__12752\,
            I => \N__12736\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12749\,
            I => \N__12736\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__12746\,
            I => \N__12736\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__12743\,
            I => \receive_module.n3631\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__12736\,
            I => \receive_module.n3631\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12731\,
            I => \bfn_13_12_0_\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12725\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__12725\,
            I => \receive_module.rx_counter.n4_adj_605\
        );

    \I__1990\ : CascadeMux
    port map (
            O => \N__12722\,
            I => \receive_module.rx_counter.n3422_cascade_\
        );

    \I__1989\ : InMux
    port map (
            O => \N__12719\,
            I => \N__12716\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__12716\,
            I => \receive_module.rx_counter.n55_adj_606\
        );

    \I__1987\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12710\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__12710\,
            I => \receive_module.rx_counter.n3394\
        );

    \I__1985\ : InMux
    port map (
            O => \N__12707\,
            I => \N__12704\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__12704\,
            I => \receive_module.rx_counter.n5\
        );

    \I__1983\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12698\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__12698\,
            I => \receive_module.rx_counter.n3413\
        );

    \I__1981\ : SRMux
    port map (
            O => \N__12695\,
            I => \N__12692\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__12692\,
            I => \N__12687\
        );

    \I__1979\ : SRMux
    port map (
            O => \N__12691\,
            I => \N__12684\
        );

    \I__1978\ : SRMux
    port map (
            O => \N__12690\,
            I => \N__12681\
        );

    \I__1977\ : Span4Mux_s2_v
    port map (
            O => \N__12687\,
            I => \N__12673\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__12684\,
            I => \N__12673\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__12681\,
            I => \N__12673\
        );

    \I__1974\ : SRMux
    port map (
            O => \N__12680\,
            I => \N__12670\
        );

    \I__1973\ : Span4Mux_v
    port map (
            O => \N__12673\,
            I => \N__12667\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__12670\,
            I => \N__12664\
        );

    \I__1971\ : Sp12to4
    port map (
            O => \N__12667\,
            I => \N__12661\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__12664\,
            I => \N__12658\
        );

    \I__1969\ : Span12Mux_v
    port map (
            O => \N__12661\,
            I => \N__12655\
        );

    \I__1968\ : Span4Mux_v
    port map (
            O => \N__12658\,
            I => \N__12652\
        );

    \I__1967\ : Span12Mux_h
    port map (
            O => \N__12655\,
            I => \N__12649\
        );

    \I__1966\ : Span4Mux_h
    port map (
            O => \N__12652\,
            I => \N__12646\
        );

    \I__1965\ : Odrv12
    port map (
            O => \N__12649\,
            I => \line_buffer.n596\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__12646\,
            I => \line_buffer.n596\
        );

    \I__1963\ : InMux
    port map (
            O => \N__12641\,
            I => \N__12638\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__12638\,
            I => \receive_module.rx_counter.n4_adj_604\
        );

    \I__1961\ : InMux
    port map (
            O => \N__12635\,
            I => \bfn_13_9_0_\
        );

    \I__1960\ : InMux
    port map (
            O => \N__12632\,
            I => \receive_module.rx_counter.n3117\
        );

    \I__1959\ : InMux
    port map (
            O => \N__12629\,
            I => \receive_module.rx_counter.n3159\
        );

    \I__1958\ : InMux
    port map (
            O => \N__12626\,
            I => \receive_module.rx_counter.n3160\
        );

    \I__1957\ : CEMux
    port map (
            O => \N__12623\,
            I => \N__12619\
        );

    \I__1956\ : CEMux
    port map (
            O => \N__12622\,
            I => \N__12616\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__12619\,
            I => \receive_module.rx_counter.n3623\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__12616\,
            I => \receive_module.rx_counter.n3623\
        );

    \I__1953\ : InMux
    port map (
            O => \N__12611\,
            I => \N__12607\
        );

    \I__1952\ : InMux
    port map (
            O => \N__12610\,
            I => \N__12604\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__12607\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__12604\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__1949\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12595\
        );

    \I__1948\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12592\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__12595\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__12592\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__1945\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12583\
        );

    \I__1944\ : InMux
    port map (
            O => \N__12586\,
            I => \N__12580\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__12583\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__12580\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__1941\ : InMux
    port map (
            O => \N__12575\,
            I => \N__12571\
        );

    \I__1940\ : InMux
    port map (
            O => \N__12574\,
            I => \N__12568\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__12571\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__12568\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__1937\ : InMux
    port map (
            O => \N__12563\,
            I => \N__12559\
        );

    \I__1936\ : InMux
    port map (
            O => \N__12562\,
            I => \N__12556\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__12559\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__12556\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__1933\ : InMux
    port map (
            O => \N__12551\,
            I => \N__12547\
        );

    \I__1932\ : InMux
    port map (
            O => \N__12550\,
            I => \N__12544\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__12547\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__12544\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__12539\,
            I => \receive_module.rx_counter.n3473_cascade_\
        );

    \I__1928\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12533\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__12533\,
            I => \receive_module.rx_counter.n7\
        );

    \I__1926\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12527\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__12527\,
            I => \N__12524\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__12524\,
            I => \receive_module.rx_counter.n11\
        );

    \I__1923\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12517\
        );

    \I__1922\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12514\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__12517\,
            I => \receive_module.rx_counter.old_VS\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__12514\,
            I => \receive_module.rx_counter.old_VS\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__12509\,
            I => \receive_module.rx_counter.n11_cascade_\
        );

    \I__1918\ : SRMux
    port map (
            O => \N__12506\,
            I => \N__12503\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__12503\,
            I => \N__12500\
        );

    \I__1916\ : Span4Mux_h
    port map (
            O => \N__12500\,
            I => \N__12497\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__12497\,
            I => \receive_module.rx_counter.n2529\
        );

    \I__1914\ : InMux
    port map (
            O => \N__12494\,
            I => \N__12491\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__12491\,
            I => \N__12488\
        );

    \I__1912\ : Span12Mux_s10_v
    port map (
            O => \N__12488\,
            I => \N__12485\
        );

    \I__1911\ : Odrv12
    port map (
            O => \N__12485\,
            I => \receive_module.n126\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__12482\,
            I => \N__12479\
        );

    \I__1909\ : CascadeBuf
    port map (
            O => \N__12479\,
            I => \N__12476\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__12476\,
            I => \N__12473\
        );

    \I__1907\ : CascadeBuf
    port map (
            O => \N__12473\,
            I => \N__12469\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__12472\,
            I => \N__12466\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__12469\,
            I => \N__12463\
        );

    \I__1904\ : CascadeBuf
    port map (
            O => \N__12466\,
            I => \N__12460\
        );

    \I__1903\ : CascadeBuf
    port map (
            O => \N__12463\,
            I => \N__12457\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__12460\,
            I => \N__12454\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__12457\,
            I => \N__12451\
        );

    \I__1900\ : CascadeBuf
    port map (
            O => \N__12454\,
            I => \N__12448\
        );

    \I__1899\ : CascadeBuf
    port map (
            O => \N__12451\,
            I => \N__12445\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__12448\,
            I => \N__12442\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__12445\,
            I => \N__12439\
        );

    \I__1896\ : CascadeBuf
    port map (
            O => \N__12442\,
            I => \N__12436\
        );

    \I__1895\ : CascadeBuf
    port map (
            O => \N__12439\,
            I => \N__12433\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__12436\,
            I => \N__12430\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__12433\,
            I => \N__12427\
        );

    \I__1892\ : CascadeBuf
    port map (
            O => \N__12430\,
            I => \N__12424\
        );

    \I__1891\ : CascadeBuf
    port map (
            O => \N__12427\,
            I => \N__12421\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__12424\,
            I => \N__12418\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__12421\,
            I => \N__12415\
        );

    \I__1888\ : CascadeBuf
    port map (
            O => \N__12418\,
            I => \N__12412\
        );

    \I__1887\ : CascadeBuf
    port map (
            O => \N__12415\,
            I => \N__12409\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__12412\,
            I => \N__12406\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__12409\,
            I => \N__12403\
        );

    \I__1884\ : CascadeBuf
    port map (
            O => \N__12406\,
            I => \N__12400\
        );

    \I__1883\ : CascadeBuf
    port map (
            O => \N__12403\,
            I => \N__12397\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__12400\,
            I => \N__12394\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__12397\,
            I => \N__12391\
        );

    \I__1880\ : CascadeBuf
    port map (
            O => \N__12394\,
            I => \N__12388\
        );

    \I__1879\ : CascadeBuf
    port map (
            O => \N__12391\,
            I => \N__12385\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__12388\,
            I => \N__12382\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__12385\,
            I => \N__12379\
        );

    \I__1876\ : CascadeBuf
    port map (
            O => \N__12382\,
            I => \N__12376\
        );

    \I__1875\ : CascadeBuf
    port map (
            O => \N__12379\,
            I => \N__12373\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__12376\,
            I => \N__12370\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__12373\,
            I => \N__12367\
        );

    \I__1872\ : CascadeBuf
    port map (
            O => \N__12370\,
            I => \N__12364\
        );

    \I__1871\ : CascadeBuf
    port map (
            O => \N__12367\,
            I => \N__12361\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__12364\,
            I => \N__12358\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__12361\,
            I => \N__12355\
        );

    \I__1868\ : CascadeBuf
    port map (
            O => \N__12358\,
            I => \N__12352\
        );

    \I__1867\ : CascadeBuf
    port map (
            O => \N__12355\,
            I => \N__12349\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__12352\,
            I => \N__12346\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__12349\,
            I => \N__12343\
        );

    \I__1864\ : CascadeBuf
    port map (
            O => \N__12346\,
            I => \N__12340\
        );

    \I__1863\ : CascadeBuf
    port map (
            O => \N__12343\,
            I => \N__12337\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__12340\,
            I => \N__12334\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__12337\,
            I => \N__12331\
        );

    \I__1860\ : CascadeBuf
    port map (
            O => \N__12334\,
            I => \N__12328\
        );

    \I__1859\ : CascadeBuf
    port map (
            O => \N__12331\,
            I => \N__12325\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__12328\,
            I => \N__12322\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__12325\,
            I => \N__12319\
        );

    \I__1856\ : CascadeBuf
    port map (
            O => \N__12322\,
            I => \N__12316\
        );

    \I__1855\ : CascadeBuf
    port map (
            O => \N__12319\,
            I => \N__12313\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__12316\,
            I => \N__12310\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__12313\,
            I => \N__12307\
        );

    \I__1852\ : CascadeBuf
    port map (
            O => \N__12310\,
            I => \N__12304\
        );

    \I__1851\ : InMux
    port map (
            O => \N__12307\,
            I => \N__12301\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__12304\,
            I => \N__12298\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__12301\,
            I => \N__12295\
        );

    \I__1848\ : CascadeBuf
    port map (
            O => \N__12298\,
            I => \N__12291\
        );

    \I__1847\ : Span4Mux_s3_v
    port map (
            O => \N__12295\,
            I => \N__12288\
        );

    \I__1846\ : InMux
    port map (
            O => \N__12294\,
            I => \N__12285\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__12291\,
            I => \N__12282\
        );

    \I__1844\ : Span4Mux_h
    port map (
            O => \N__12288\,
            I => \N__12279\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__12285\,
            I => \N__12276\
        );

    \I__1842\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12273\
        );

    \I__1841\ : Span4Mux_h
    port map (
            O => \N__12279\,
            I => \N__12270\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__12276\,
            I => \N__12266\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__12273\,
            I => \N__12263\
        );

    \I__1838\ : Span4Mux_h
    port map (
            O => \N__12270\,
            I => \N__12260\
        );

    \I__1837\ : InMux
    port map (
            O => \N__12269\,
            I => \N__12257\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__12266\,
            I => \N__12254\
        );

    \I__1835\ : Span12Mux_s9_v
    port map (
            O => \N__12263\,
            I => \N__12251\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__12260\,
            I => \N__12248\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__12257\,
            I => \RX_ADDR_10\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__12254\,
            I => \RX_ADDR_10\
        );

    \I__1831\ : Odrv12
    port map (
            O => \N__12251\,
            I => \RX_ADDR_10\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__12248\,
            I => \RX_ADDR_10\
        );

    \I__1829\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12236\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__12236\,
            I => \N__12233\
        );

    \I__1827\ : Span12Mux_s10_v
    port map (
            O => \N__12233\,
            I => \N__12230\
        );

    \I__1826\ : Odrv12
    port map (
            O => \N__12230\,
            I => \receive_module.n133\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__12227\,
            I => \N__12224\
        );

    \I__1824\ : CascadeBuf
    port map (
            O => \N__12224\,
            I => \N__12221\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__12221\,
            I => \N__12217\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__12220\,
            I => \N__12214\
        );

    \I__1821\ : CascadeBuf
    port map (
            O => \N__12217\,
            I => \N__12211\
        );

    \I__1820\ : CascadeBuf
    port map (
            O => \N__12214\,
            I => \N__12208\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__12211\,
            I => \N__12205\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__12208\,
            I => \N__12202\
        );

    \I__1817\ : CascadeBuf
    port map (
            O => \N__12205\,
            I => \N__12199\
        );

    \I__1816\ : CascadeBuf
    port map (
            O => \N__12202\,
            I => \N__12196\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__12199\,
            I => \N__12193\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__12196\,
            I => \N__12190\
        );

    \I__1813\ : CascadeBuf
    port map (
            O => \N__12193\,
            I => \N__12187\
        );

    \I__1812\ : CascadeBuf
    port map (
            O => \N__12190\,
            I => \N__12184\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__12187\,
            I => \N__12181\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__12184\,
            I => \N__12178\
        );

    \I__1809\ : CascadeBuf
    port map (
            O => \N__12181\,
            I => \N__12175\
        );

    \I__1808\ : CascadeBuf
    port map (
            O => \N__12178\,
            I => \N__12172\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__12175\,
            I => \N__12169\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__12172\,
            I => \N__12166\
        );

    \I__1805\ : CascadeBuf
    port map (
            O => \N__12169\,
            I => \N__12163\
        );

    \I__1804\ : CascadeBuf
    port map (
            O => \N__12166\,
            I => \N__12160\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__12163\,
            I => \N__12157\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__12160\,
            I => \N__12154\
        );

    \I__1801\ : CascadeBuf
    port map (
            O => \N__12157\,
            I => \N__12151\
        );

    \I__1800\ : CascadeBuf
    port map (
            O => \N__12154\,
            I => \N__12148\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__12151\,
            I => \N__12145\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__12148\,
            I => \N__12142\
        );

    \I__1797\ : CascadeBuf
    port map (
            O => \N__12145\,
            I => \N__12139\
        );

    \I__1796\ : CascadeBuf
    port map (
            O => \N__12142\,
            I => \N__12136\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__12139\,
            I => \N__12133\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__12136\,
            I => \N__12130\
        );

    \I__1793\ : CascadeBuf
    port map (
            O => \N__12133\,
            I => \N__12127\
        );

    \I__1792\ : CascadeBuf
    port map (
            O => \N__12130\,
            I => \N__12124\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__12127\,
            I => \N__12121\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__12124\,
            I => \N__12118\
        );

    \I__1789\ : CascadeBuf
    port map (
            O => \N__12121\,
            I => \N__12115\
        );

    \I__1788\ : CascadeBuf
    port map (
            O => \N__12118\,
            I => \N__12112\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__12115\,
            I => \N__12109\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__12112\,
            I => \N__12106\
        );

    \I__1785\ : CascadeBuf
    port map (
            O => \N__12109\,
            I => \N__12103\
        );

    \I__1784\ : CascadeBuf
    port map (
            O => \N__12106\,
            I => \N__12100\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__12103\,
            I => \N__12097\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__12100\,
            I => \N__12094\
        );

    \I__1781\ : CascadeBuf
    port map (
            O => \N__12097\,
            I => \N__12091\
        );

    \I__1780\ : CascadeBuf
    port map (
            O => \N__12094\,
            I => \N__12088\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__12091\,
            I => \N__12085\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__12088\,
            I => \N__12082\
        );

    \I__1777\ : CascadeBuf
    port map (
            O => \N__12085\,
            I => \N__12079\
        );

    \I__1776\ : CascadeBuf
    port map (
            O => \N__12082\,
            I => \N__12076\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__12079\,
            I => \N__12073\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__12076\,
            I => \N__12070\
        );

    \I__1773\ : CascadeBuf
    port map (
            O => \N__12073\,
            I => \N__12067\
        );

    \I__1772\ : CascadeBuf
    port map (
            O => \N__12070\,
            I => \N__12064\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__12067\,
            I => \N__12061\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__12064\,
            I => \N__12058\
        );

    \I__1769\ : CascadeBuf
    port map (
            O => \N__12061\,
            I => \N__12055\
        );

    \I__1768\ : CascadeBuf
    port map (
            O => \N__12058\,
            I => \N__12052\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__12055\,
            I => \N__12049\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__12052\,
            I => \N__12046\
        );

    \I__1765\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12042\
        );

    \I__1764\ : CascadeBuf
    port map (
            O => \N__12046\,
            I => \N__12039\
        );

    \I__1763\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12036\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__12042\,
            I => \N__12033\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__12039\,
            I => \N__12030\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__12036\,
            I => \N__12027\
        );

    \I__1759\ : Span4Mux_s3_v
    port map (
            O => \N__12033\,
            I => \N__12024\
        );

    \I__1758\ : InMux
    port map (
            O => \N__12030\,
            I => \N__12021\
        );

    \I__1757\ : Sp12to4
    port map (
            O => \N__12027\,
            I => \N__12018\
        );

    \I__1756\ : Span4Mux_h
    port map (
            O => \N__12024\,
            I => \N__12014\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__12021\,
            I => \N__12011\
        );

    \I__1754\ : Span12Mux_v
    port map (
            O => \N__12018\,
            I => \N__12008\
        );

    \I__1753\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12005\
        );

    \I__1752\ : Sp12to4
    port map (
            O => \N__12014\,
            I => \N__12002\
        );

    \I__1751\ : Span4Mux_h
    port map (
            O => \N__12011\,
            I => \N__11999\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__12008\,
            I => \RX_ADDR_3\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__12005\,
            I => \RX_ADDR_3\
        );

    \I__1748\ : Odrv12
    port map (
            O => \N__12002\,
            I => \RX_ADDR_3\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__11999\,
            I => \RX_ADDR_3\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11990\,
            I => \N__11987\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__11987\,
            I => \N__11984\
        );

    \I__1744\ : Span4Mux_v
    port map (
            O => \N__11984\,
            I => \N__11981\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__11981\,
            I => \N__11978\
        );

    \I__1742\ : Span4Mux_v
    port map (
            O => \N__11978\,
            I => \N__11975\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__11975\,
            I => \N__11972\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__11972\,
            I => \receive_module.n132\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__11969\,
            I => \N__11966\
        );

    \I__1738\ : CascadeBuf
    port map (
            O => \N__11966\,
            I => \N__11963\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__11963\,
            I => \N__11959\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__11962\,
            I => \N__11956\
        );

    \I__1735\ : CascadeBuf
    port map (
            O => \N__11959\,
            I => \N__11953\
        );

    \I__1734\ : CascadeBuf
    port map (
            O => \N__11956\,
            I => \N__11950\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__11953\,
            I => \N__11947\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__11950\,
            I => \N__11944\
        );

    \I__1731\ : CascadeBuf
    port map (
            O => \N__11947\,
            I => \N__11941\
        );

    \I__1730\ : CascadeBuf
    port map (
            O => \N__11944\,
            I => \N__11938\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__11941\,
            I => \N__11935\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__11938\,
            I => \N__11932\
        );

    \I__1727\ : CascadeBuf
    port map (
            O => \N__11935\,
            I => \N__11929\
        );

    \I__1726\ : CascadeBuf
    port map (
            O => \N__11932\,
            I => \N__11926\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__11929\,
            I => \N__11923\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__11926\,
            I => \N__11920\
        );

    \I__1723\ : CascadeBuf
    port map (
            O => \N__11923\,
            I => \N__11917\
        );

    \I__1722\ : CascadeBuf
    port map (
            O => \N__11920\,
            I => \N__11914\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__11917\,
            I => \N__11911\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__11914\,
            I => \N__11908\
        );

    \I__1719\ : CascadeBuf
    port map (
            O => \N__11911\,
            I => \N__11905\
        );

    \I__1718\ : CascadeBuf
    port map (
            O => \N__11908\,
            I => \N__11902\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__11905\,
            I => \N__11899\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__11902\,
            I => \N__11896\
        );

    \I__1715\ : CascadeBuf
    port map (
            O => \N__11899\,
            I => \N__11893\
        );

    \I__1714\ : CascadeBuf
    port map (
            O => \N__11896\,
            I => \N__11890\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__11893\,
            I => \N__11887\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__11890\,
            I => \N__11884\
        );

    \I__1711\ : CascadeBuf
    port map (
            O => \N__11887\,
            I => \N__11881\
        );

    \I__1710\ : CascadeBuf
    port map (
            O => \N__11884\,
            I => \N__11878\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__11881\,
            I => \N__11875\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__11878\,
            I => \N__11872\
        );

    \I__1707\ : CascadeBuf
    port map (
            O => \N__11875\,
            I => \N__11869\
        );

    \I__1706\ : CascadeBuf
    port map (
            O => \N__11872\,
            I => \N__11866\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__11869\,
            I => \N__11863\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__11866\,
            I => \N__11860\
        );

    \I__1703\ : CascadeBuf
    port map (
            O => \N__11863\,
            I => \N__11857\
        );

    \I__1702\ : CascadeBuf
    port map (
            O => \N__11860\,
            I => \N__11854\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__11857\,
            I => \N__11851\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__11854\,
            I => \N__11848\
        );

    \I__1699\ : CascadeBuf
    port map (
            O => \N__11851\,
            I => \N__11845\
        );

    \I__1698\ : CascadeBuf
    port map (
            O => \N__11848\,
            I => \N__11842\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__11845\,
            I => \N__11839\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__11842\,
            I => \N__11836\
        );

    \I__1695\ : CascadeBuf
    port map (
            O => \N__11839\,
            I => \N__11833\
        );

    \I__1694\ : CascadeBuf
    port map (
            O => \N__11836\,
            I => \N__11830\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__11833\,
            I => \N__11827\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__11830\,
            I => \N__11824\
        );

    \I__1691\ : CascadeBuf
    port map (
            O => \N__11827\,
            I => \N__11821\
        );

    \I__1690\ : CascadeBuf
    port map (
            O => \N__11824\,
            I => \N__11818\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__11821\,
            I => \N__11815\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__11818\,
            I => \N__11812\
        );

    \I__1687\ : CascadeBuf
    port map (
            O => \N__11815\,
            I => \N__11809\
        );

    \I__1686\ : CascadeBuf
    port map (
            O => \N__11812\,
            I => \N__11806\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__11809\,
            I => \N__11803\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__11806\,
            I => \N__11800\
        );

    \I__1683\ : CascadeBuf
    port map (
            O => \N__11803\,
            I => \N__11797\
        );

    \I__1682\ : CascadeBuf
    port map (
            O => \N__11800\,
            I => \N__11794\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__11797\,
            I => \N__11791\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__11794\,
            I => \N__11788\
        );

    \I__1679\ : InMux
    port map (
            O => \N__11791\,
            I => \N__11784\
        );

    \I__1678\ : CascadeBuf
    port map (
            O => \N__11788\,
            I => \N__11781\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11787\,
            I => \N__11778\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__11784\,
            I => \N__11775\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__11781\,
            I => \N__11772\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__11778\,
            I => \N__11769\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__11775\,
            I => \N__11766\
        );

    \I__1672\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11763\
        );

    \I__1671\ : Sp12to4
    port map (
            O => \N__11769\,
            I => \N__11760\
        );

    \I__1670\ : Sp12to4
    port map (
            O => \N__11766\,
            I => \N__11756\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__11763\,
            I => \N__11753\
        );

    \I__1668\ : Span12Mux_v
    port map (
            O => \N__11760\,
            I => \N__11750\
        );

    \I__1667\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11747\
        );

    \I__1666\ : Span12Mux_s2_v
    port map (
            O => \N__11756\,
            I => \N__11744\
        );

    \I__1665\ : Span4Mux_s2_v
    port map (
            O => \N__11753\,
            I => \N__11741\
        );

    \I__1664\ : Odrv12
    port map (
            O => \N__11750\,
            I => \RX_ADDR_4\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__11747\,
            I => \RX_ADDR_4\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__11744\,
            I => \RX_ADDR_4\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__11741\,
            I => \RX_ADDR_4\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__11729\,
            I => \N__11726\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__11726\,
            I => \tvp_video_buffer.BUFFER_1_2\
        );

    \I__1657\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11718\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11722\,
            I => \N__11713\
        );

    \I__1655\ : InMux
    port map (
            O => \N__11721\,
            I => \N__11709\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__11718\,
            I => \N__11706\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11703\
        );

    \I__1652\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11700\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__11713\,
            I => \N__11695\
        );

    \I__1650\ : InMux
    port map (
            O => \N__11712\,
            I => \N__11692\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__11709\,
            I => \N__11689\
        );

    \I__1648\ : Span12Mux_s4_v
    port map (
            O => \N__11706\,
            I => \N__11682\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__11703\,
            I => \N__11682\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__11700\,
            I => \N__11682\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11679\
        );

    \I__1644\ : InMux
    port map (
            O => \N__11698\,
            I => \N__11676\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__11695\,
            I => \N__11673\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__11692\,
            I => \N__11670\
        );

    \I__1641\ : Span12Mux_h
    port map (
            O => \N__11689\,
            I => \N__11667\
        );

    \I__1640\ : Span12Mux_v
    port map (
            O => \N__11682\,
            I => \N__11660\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__11679\,
            I => \N__11660\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11676\,
            I => \N__11660\
        );

    \I__1637\ : Span4Mux_v
    port map (
            O => \N__11673\,
            I => \N__11655\
        );

    \I__1636\ : Span4Mux_h
    port map (
            O => \N__11670\,
            I => \N__11655\
        );

    \I__1635\ : Span12Mux_v
    port map (
            O => \N__11667\,
            I => \N__11652\
        );

    \I__1634\ : Span12Mux_v
    port map (
            O => \N__11660\,
            I => \N__11649\
        );

    \I__1633\ : Span4Mux_h
    port map (
            O => \N__11655\,
            I => \N__11646\
        );

    \I__1632\ : Odrv12
    port map (
            O => \N__11652\,
            I => \RX_DATA_0\
        );

    \I__1631\ : Odrv12
    port map (
            O => \N__11649\,
            I => \RX_DATA_0\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__11646\,
            I => \RX_DATA_0\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11639\,
            I => \bfn_13_6_0_\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11636\,
            I => \receive_module.rx_counter.n3156\
        );

    \I__1627\ : InMux
    port map (
            O => \N__11633\,
            I => \receive_module.rx_counter.n3157\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11630\,
            I => \receive_module.rx_counter.n3158\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__11624\,
            I => \N__11621\
        );

    \I__1623\ : Span4Mux_h
    port map (
            O => \N__11621\,
            I => \N__11618\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__11618\,
            I => \transmit_module.Y_DELTA_PATTERN_7\
        );

    \I__1621\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__11612\,
            I => \transmit_module.Y_DELTA_PATTERN_6\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__1617\ : Span12Mux_v
    port map (
            O => \N__11603\,
            I => \N__11600\
        );

    \I__1616\ : Odrv12
    port map (
            O => \N__11600\,
            I => \receive_module.n131\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__11597\,
            I => \N__11593\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__11596\,
            I => \N__11590\
        );

    \I__1613\ : CascadeBuf
    port map (
            O => \N__11593\,
            I => \N__11587\
        );

    \I__1612\ : CascadeBuf
    port map (
            O => \N__11590\,
            I => \N__11584\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__11587\,
            I => \N__11581\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__11584\,
            I => \N__11578\
        );

    \I__1609\ : CascadeBuf
    port map (
            O => \N__11581\,
            I => \N__11575\
        );

    \I__1608\ : CascadeBuf
    port map (
            O => \N__11578\,
            I => \N__11572\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__11575\,
            I => \N__11569\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__11572\,
            I => \N__11566\
        );

    \I__1605\ : CascadeBuf
    port map (
            O => \N__11569\,
            I => \N__11563\
        );

    \I__1604\ : CascadeBuf
    port map (
            O => \N__11566\,
            I => \N__11560\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__11563\,
            I => \N__11557\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__11560\,
            I => \N__11554\
        );

    \I__1601\ : CascadeBuf
    port map (
            O => \N__11557\,
            I => \N__11551\
        );

    \I__1600\ : CascadeBuf
    port map (
            O => \N__11554\,
            I => \N__11548\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__11551\,
            I => \N__11545\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__11548\,
            I => \N__11542\
        );

    \I__1597\ : CascadeBuf
    port map (
            O => \N__11545\,
            I => \N__11539\
        );

    \I__1596\ : CascadeBuf
    port map (
            O => \N__11542\,
            I => \N__11536\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__11539\,
            I => \N__11533\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__11536\,
            I => \N__11530\
        );

    \I__1593\ : CascadeBuf
    port map (
            O => \N__11533\,
            I => \N__11527\
        );

    \I__1592\ : CascadeBuf
    port map (
            O => \N__11530\,
            I => \N__11524\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__11527\,
            I => \N__11521\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__11524\,
            I => \N__11518\
        );

    \I__1589\ : CascadeBuf
    port map (
            O => \N__11521\,
            I => \N__11515\
        );

    \I__1588\ : CascadeBuf
    port map (
            O => \N__11518\,
            I => \N__11512\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__11515\,
            I => \N__11509\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__11512\,
            I => \N__11506\
        );

    \I__1585\ : CascadeBuf
    port map (
            O => \N__11509\,
            I => \N__11503\
        );

    \I__1584\ : CascadeBuf
    port map (
            O => \N__11506\,
            I => \N__11500\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__11503\,
            I => \N__11497\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__11500\,
            I => \N__11494\
        );

    \I__1581\ : CascadeBuf
    port map (
            O => \N__11497\,
            I => \N__11491\
        );

    \I__1580\ : CascadeBuf
    port map (
            O => \N__11494\,
            I => \N__11488\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__11491\,
            I => \N__11485\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__11488\,
            I => \N__11482\
        );

    \I__1577\ : CascadeBuf
    port map (
            O => \N__11485\,
            I => \N__11479\
        );

    \I__1576\ : CascadeBuf
    port map (
            O => \N__11482\,
            I => \N__11476\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__11479\,
            I => \N__11473\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__11476\,
            I => \N__11470\
        );

    \I__1573\ : CascadeBuf
    port map (
            O => \N__11473\,
            I => \N__11467\
        );

    \I__1572\ : CascadeBuf
    port map (
            O => \N__11470\,
            I => \N__11464\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__11467\,
            I => \N__11461\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__11464\,
            I => \N__11458\
        );

    \I__1569\ : CascadeBuf
    port map (
            O => \N__11461\,
            I => \N__11455\
        );

    \I__1568\ : CascadeBuf
    port map (
            O => \N__11458\,
            I => \N__11452\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__11455\,
            I => \N__11449\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__11452\,
            I => \N__11446\
        );

    \I__1565\ : CascadeBuf
    port map (
            O => \N__11449\,
            I => \N__11443\
        );

    \I__1564\ : CascadeBuf
    port map (
            O => \N__11446\,
            I => \N__11440\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__11443\,
            I => \N__11437\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__11440\,
            I => \N__11434\
        );

    \I__1561\ : CascadeBuf
    port map (
            O => \N__11437\,
            I => \N__11431\
        );

    \I__1560\ : CascadeBuf
    port map (
            O => \N__11434\,
            I => \N__11428\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \N__11425\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__11428\,
            I => \N__11422\
        );

    \I__1557\ : CascadeBuf
    port map (
            O => \N__11425\,
            I => \N__11419\
        );

    \I__1556\ : CascadeBuf
    port map (
            O => \N__11422\,
            I => \N__11416\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__11419\,
            I => \N__11413\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__11416\,
            I => \N__11410\
        );

    \I__1553\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11407\
        );

    \I__1552\ : InMux
    port map (
            O => \N__11410\,
            I => \N__11404\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__11407\,
            I => \N__11400\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__11404\,
            I => \N__11397\
        );

    \I__1549\ : InMux
    port map (
            O => \N__11403\,
            I => \N__11394\
        );

    \I__1548\ : Span4Mux_s1_v
    port map (
            O => \N__11400\,
            I => \N__11391\
        );

    \I__1547\ : Span4Mux_s1_v
    port map (
            O => \N__11397\,
            I => \N__11388\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__11394\,
            I => \N__11385\
        );

    \I__1545\ : Span4Mux_h
    port map (
            O => \N__11391\,
            I => \N__11382\
        );

    \I__1544\ : Span4Mux_v
    port map (
            O => \N__11388\,
            I => \N__11379\
        );

    \I__1543\ : Span4Mux_h
    port map (
            O => \N__11385\,
            I => \N__11375\
        );

    \I__1542\ : Sp12to4
    port map (
            O => \N__11382\,
            I => \N__11372\
        );

    \I__1541\ : Sp12to4
    port map (
            O => \N__11379\,
            I => \N__11369\
        );

    \I__1540\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11366\
        );

    \I__1539\ : Span4Mux_v
    port map (
            O => \N__11375\,
            I => \N__11363\
        );

    \I__1538\ : Span12Mux_s5_v
    port map (
            O => \N__11372\,
            I => \N__11358\
        );

    \I__1537\ : Span12Mux_h
    port map (
            O => \N__11369\,
            I => \N__11358\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__11366\,
            I => \RX_ADDR_5\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__11363\,
            I => \RX_ADDR_5\
        );

    \I__1534\ : Odrv12
    port map (
            O => \N__11358\,
            I => \RX_ADDR_5\
        );

    \I__1533\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11348\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__11348\,
            I => \N__11345\
        );

    \I__1531\ : Span4Mux_v
    port map (
            O => \N__11345\,
            I => \N__11342\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__11339\,
            I => \receive_module.n130\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__11336\,
            I => \N__11332\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__11335\,
            I => \N__11329\
        );

    \I__1526\ : CascadeBuf
    port map (
            O => \N__11332\,
            I => \N__11326\
        );

    \I__1525\ : CascadeBuf
    port map (
            O => \N__11329\,
            I => \N__11323\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__11326\,
            I => \N__11320\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__11323\,
            I => \N__11317\
        );

    \I__1522\ : CascadeBuf
    port map (
            O => \N__11320\,
            I => \N__11314\
        );

    \I__1521\ : CascadeBuf
    port map (
            O => \N__11317\,
            I => \N__11311\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__11314\,
            I => \N__11308\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__11311\,
            I => \N__11305\
        );

    \I__1518\ : CascadeBuf
    port map (
            O => \N__11308\,
            I => \N__11302\
        );

    \I__1517\ : CascadeBuf
    port map (
            O => \N__11305\,
            I => \N__11299\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__11302\,
            I => \N__11296\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__11299\,
            I => \N__11293\
        );

    \I__1514\ : CascadeBuf
    port map (
            O => \N__11296\,
            I => \N__11290\
        );

    \I__1513\ : CascadeBuf
    port map (
            O => \N__11293\,
            I => \N__11287\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__11290\,
            I => \N__11284\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__11287\,
            I => \N__11281\
        );

    \I__1510\ : CascadeBuf
    port map (
            O => \N__11284\,
            I => \N__11278\
        );

    \I__1509\ : CascadeBuf
    port map (
            O => \N__11281\,
            I => \N__11275\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__11278\,
            I => \N__11272\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__11275\,
            I => \N__11269\
        );

    \I__1506\ : CascadeBuf
    port map (
            O => \N__11272\,
            I => \N__11266\
        );

    \I__1505\ : CascadeBuf
    port map (
            O => \N__11269\,
            I => \N__11263\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__11266\,
            I => \N__11260\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__11263\,
            I => \N__11257\
        );

    \I__1502\ : CascadeBuf
    port map (
            O => \N__11260\,
            I => \N__11254\
        );

    \I__1501\ : CascadeBuf
    port map (
            O => \N__11257\,
            I => \N__11251\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__11254\,
            I => \N__11248\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__11251\,
            I => \N__11245\
        );

    \I__1498\ : CascadeBuf
    port map (
            O => \N__11248\,
            I => \N__11242\
        );

    \I__1497\ : CascadeBuf
    port map (
            O => \N__11245\,
            I => \N__11239\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__11242\,
            I => \N__11236\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__11239\,
            I => \N__11233\
        );

    \I__1494\ : CascadeBuf
    port map (
            O => \N__11236\,
            I => \N__11230\
        );

    \I__1493\ : CascadeBuf
    port map (
            O => \N__11233\,
            I => \N__11227\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__11230\,
            I => \N__11224\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__11227\,
            I => \N__11221\
        );

    \I__1490\ : CascadeBuf
    port map (
            O => \N__11224\,
            I => \N__11218\
        );

    \I__1489\ : CascadeBuf
    port map (
            O => \N__11221\,
            I => \N__11215\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__11218\,
            I => \N__11212\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__11215\,
            I => \N__11209\
        );

    \I__1486\ : CascadeBuf
    port map (
            O => \N__11212\,
            I => \N__11206\
        );

    \I__1485\ : CascadeBuf
    port map (
            O => \N__11209\,
            I => \N__11203\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__11206\,
            I => \N__11200\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__11203\,
            I => \N__11197\
        );

    \I__1482\ : CascadeBuf
    port map (
            O => \N__11200\,
            I => \N__11194\
        );

    \I__1481\ : CascadeBuf
    port map (
            O => \N__11197\,
            I => \N__11191\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__11194\,
            I => \N__11188\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__11191\,
            I => \N__11185\
        );

    \I__1478\ : CascadeBuf
    port map (
            O => \N__11188\,
            I => \N__11182\
        );

    \I__1477\ : CascadeBuf
    port map (
            O => \N__11185\,
            I => \N__11179\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__11182\,
            I => \N__11176\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__11179\,
            I => \N__11173\
        );

    \I__1474\ : CascadeBuf
    port map (
            O => \N__11176\,
            I => \N__11170\
        );

    \I__1473\ : CascadeBuf
    port map (
            O => \N__11173\,
            I => \N__11167\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__11170\,
            I => \N__11164\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__11167\,
            I => \N__11161\
        );

    \I__1470\ : CascadeBuf
    port map (
            O => \N__11164\,
            I => \N__11158\
        );

    \I__1469\ : CascadeBuf
    port map (
            O => \N__11161\,
            I => \N__11155\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__11158\,
            I => \N__11152\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__11155\,
            I => \N__11149\
        );

    \I__1466\ : InMux
    port map (
            O => \N__11152\,
            I => \N__11146\
        );

    \I__1465\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11142\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__11146\,
            I => \N__11139\
        );

    \I__1463\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11136\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__11142\,
            I => \N__11133\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__11139\,
            I => \N__11130\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__11136\,
            I => \N__11126\
        );

    \I__1459\ : Span4Mux_h
    port map (
            O => \N__11133\,
            I => \N__11123\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__11130\,
            I => \N__11120\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__11129\,
            I => \N__11117\
        );

    \I__1456\ : Span4Mux_h
    port map (
            O => \N__11126\,
            I => \N__11114\
        );

    \I__1455\ : Sp12to4
    port map (
            O => \N__11123\,
            I => \N__11111\
        );

    \I__1454\ : Sp12to4
    port map (
            O => \N__11120\,
            I => \N__11108\
        );

    \I__1453\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11105\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__11114\,
            I => \N__11102\
        );

    \I__1451\ : Span12Mux_v
    port map (
            O => \N__11111\,
            I => \N__11097\
        );

    \I__1450\ : Span12Mux_v
    port map (
            O => \N__11108\,
            I => \N__11097\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__11105\,
            I => \RX_ADDR_6\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__11102\,
            I => \RX_ADDR_6\
        );

    \I__1447\ : Odrv12
    port map (
            O => \N__11097\,
            I => \RX_ADDR_6\
        );

    \I__1446\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1444\ : Sp12to4
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__1443\ : Odrv12
    port map (
            O => \N__11081\,
            I => \receive_module.n129\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__11078\,
            I => \N__11074\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__11077\,
            I => \N__11071\
        );

    \I__1440\ : CascadeBuf
    port map (
            O => \N__11074\,
            I => \N__11068\
        );

    \I__1439\ : CascadeBuf
    port map (
            O => \N__11071\,
            I => \N__11065\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__11068\,
            I => \N__11062\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__11065\,
            I => \N__11059\
        );

    \I__1436\ : CascadeBuf
    port map (
            O => \N__11062\,
            I => \N__11056\
        );

    \I__1435\ : CascadeBuf
    port map (
            O => \N__11059\,
            I => \N__11053\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__11056\,
            I => \N__11050\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__11053\,
            I => \N__11047\
        );

    \I__1432\ : CascadeBuf
    port map (
            O => \N__11050\,
            I => \N__11044\
        );

    \I__1431\ : CascadeBuf
    port map (
            O => \N__11047\,
            I => \N__11041\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__11044\,
            I => \N__11038\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__11041\,
            I => \N__11035\
        );

    \I__1428\ : CascadeBuf
    port map (
            O => \N__11038\,
            I => \N__11032\
        );

    \I__1427\ : CascadeBuf
    port map (
            O => \N__11035\,
            I => \N__11029\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__11032\,
            I => \N__11026\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__11029\,
            I => \N__11023\
        );

    \I__1424\ : CascadeBuf
    port map (
            O => \N__11026\,
            I => \N__11020\
        );

    \I__1423\ : CascadeBuf
    port map (
            O => \N__11023\,
            I => \N__11017\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__11020\,
            I => \N__11014\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__11017\,
            I => \N__11011\
        );

    \I__1420\ : CascadeBuf
    port map (
            O => \N__11014\,
            I => \N__11008\
        );

    \I__1419\ : CascadeBuf
    port map (
            O => \N__11011\,
            I => \N__11005\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__11008\,
            I => \N__11002\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__11005\,
            I => \N__10999\
        );

    \I__1416\ : CascadeBuf
    port map (
            O => \N__11002\,
            I => \N__10996\
        );

    \I__1415\ : CascadeBuf
    port map (
            O => \N__10999\,
            I => \N__10993\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__10996\,
            I => \N__10990\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__10993\,
            I => \N__10987\
        );

    \I__1412\ : CascadeBuf
    port map (
            O => \N__10990\,
            I => \N__10984\
        );

    \I__1411\ : CascadeBuf
    port map (
            O => \N__10987\,
            I => \N__10981\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__10984\,
            I => \N__10978\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__10981\,
            I => \N__10975\
        );

    \I__1408\ : CascadeBuf
    port map (
            O => \N__10978\,
            I => \N__10972\
        );

    \I__1407\ : CascadeBuf
    port map (
            O => \N__10975\,
            I => \N__10969\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__10972\,
            I => \N__10966\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__10969\,
            I => \N__10963\
        );

    \I__1404\ : CascadeBuf
    port map (
            O => \N__10966\,
            I => \N__10960\
        );

    \I__1403\ : CascadeBuf
    port map (
            O => \N__10963\,
            I => \N__10957\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__10960\,
            I => \N__10954\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__10957\,
            I => \N__10951\
        );

    \I__1400\ : CascadeBuf
    port map (
            O => \N__10954\,
            I => \N__10948\
        );

    \I__1399\ : CascadeBuf
    port map (
            O => \N__10951\,
            I => \N__10945\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__10948\,
            I => \N__10942\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__10945\,
            I => \N__10939\
        );

    \I__1396\ : CascadeBuf
    port map (
            O => \N__10942\,
            I => \N__10936\
        );

    \I__1395\ : CascadeBuf
    port map (
            O => \N__10939\,
            I => \N__10933\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__10936\,
            I => \N__10930\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__10933\,
            I => \N__10927\
        );

    \I__1392\ : CascadeBuf
    port map (
            O => \N__10930\,
            I => \N__10924\
        );

    \I__1391\ : CascadeBuf
    port map (
            O => \N__10927\,
            I => \N__10921\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10924\,
            I => \N__10918\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__10921\,
            I => \N__10915\
        );

    \I__1388\ : CascadeBuf
    port map (
            O => \N__10918\,
            I => \N__10912\
        );

    \I__1387\ : CascadeBuf
    port map (
            O => \N__10915\,
            I => \N__10909\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__10912\,
            I => \N__10906\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__10909\,
            I => \N__10903\
        );

    \I__1384\ : CascadeBuf
    port map (
            O => \N__10906\,
            I => \N__10900\
        );

    \I__1383\ : CascadeBuf
    port map (
            O => \N__10903\,
            I => \N__10897\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__10900\,
            I => \N__10894\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__10897\,
            I => \N__10891\
        );

    \I__1380\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10888\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10885\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__10888\,
            I => \N__10882\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10885\,
            I => \N__10879\
        );

    \I__1376\ : Span4Mux_s1_v
    port map (
            O => \N__10882\,
            I => \N__10876\
        );

    \I__1375\ : Span4Mux_s2_v
    port map (
            O => \N__10879\,
            I => \N__10873\
        );

    \I__1374\ : Sp12to4
    port map (
            O => \N__10876\,
            I => \N__10869\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__10873\,
            I => \N__10866\
        );

    \I__1372\ : InMux
    port map (
            O => \N__10872\,
            I => \N__10863\
        );

    \I__1371\ : Span12Mux_h
    port map (
            O => \N__10869\,
            I => \N__10859\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__10866\,
            I => \N__10856\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__10863\,
            I => \N__10853\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10850\
        );

    \I__1367\ : Span12Mux_v
    port map (
            O => \N__10859\,
            I => \N__10847\
        );

    \I__1366\ : Span4Mux_v
    port map (
            O => \N__10856\,
            I => \N__10844\
        );

    \I__1365\ : Odrv12
    port map (
            O => \N__10853\,
            I => \RX_ADDR_7\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__10850\,
            I => \RX_ADDR_7\
        );

    \I__1363\ : Odrv12
    port map (
            O => \N__10847\,
            I => \RX_ADDR_7\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__10844\,
            I => \RX_ADDR_7\
        );

    \I__1361\ : InMux
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1359\ : Odrv12
    port map (
            O => \N__10829\,
            I => \receive_module.n128\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__10826\,
            I => \N__10822\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__10825\,
            I => \N__10819\
        );

    \I__1356\ : CascadeBuf
    port map (
            O => \N__10822\,
            I => \N__10816\
        );

    \I__1355\ : CascadeBuf
    port map (
            O => \N__10819\,
            I => \N__10813\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__10816\,
            I => \N__10810\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__10813\,
            I => \N__10807\
        );

    \I__1352\ : CascadeBuf
    port map (
            O => \N__10810\,
            I => \N__10804\
        );

    \I__1351\ : CascadeBuf
    port map (
            O => \N__10807\,
            I => \N__10801\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__10804\,
            I => \N__10798\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__10801\,
            I => \N__10795\
        );

    \I__1348\ : CascadeBuf
    port map (
            O => \N__10798\,
            I => \N__10792\
        );

    \I__1347\ : CascadeBuf
    port map (
            O => \N__10795\,
            I => \N__10789\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__10792\,
            I => \N__10786\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__10789\,
            I => \N__10783\
        );

    \I__1344\ : CascadeBuf
    port map (
            O => \N__10786\,
            I => \N__10780\
        );

    \I__1343\ : CascadeBuf
    port map (
            O => \N__10783\,
            I => \N__10777\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__10780\,
            I => \N__10774\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__10777\,
            I => \N__10771\
        );

    \I__1340\ : CascadeBuf
    port map (
            O => \N__10774\,
            I => \N__10768\
        );

    \I__1339\ : CascadeBuf
    port map (
            O => \N__10771\,
            I => \N__10765\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__10768\,
            I => \N__10762\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__10765\,
            I => \N__10759\
        );

    \I__1336\ : CascadeBuf
    port map (
            O => \N__10762\,
            I => \N__10756\
        );

    \I__1335\ : CascadeBuf
    port map (
            O => \N__10759\,
            I => \N__10753\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__10756\,
            I => \N__10750\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__10753\,
            I => \N__10747\
        );

    \I__1332\ : CascadeBuf
    port map (
            O => \N__10750\,
            I => \N__10744\
        );

    \I__1331\ : CascadeBuf
    port map (
            O => \N__10747\,
            I => \N__10741\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__10744\,
            I => \N__10738\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__10741\,
            I => \N__10735\
        );

    \I__1328\ : CascadeBuf
    port map (
            O => \N__10738\,
            I => \N__10732\
        );

    \I__1327\ : CascadeBuf
    port map (
            O => \N__10735\,
            I => \N__10729\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__10732\,
            I => \N__10726\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__10729\,
            I => \N__10723\
        );

    \I__1324\ : CascadeBuf
    port map (
            O => \N__10726\,
            I => \N__10720\
        );

    \I__1323\ : CascadeBuf
    port map (
            O => \N__10723\,
            I => \N__10717\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__10720\,
            I => \N__10714\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__10717\,
            I => \N__10711\
        );

    \I__1320\ : CascadeBuf
    port map (
            O => \N__10714\,
            I => \N__10708\
        );

    \I__1319\ : CascadeBuf
    port map (
            O => \N__10711\,
            I => \N__10705\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__10708\,
            I => \N__10702\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__10705\,
            I => \N__10699\
        );

    \I__1316\ : CascadeBuf
    port map (
            O => \N__10702\,
            I => \N__10696\
        );

    \I__1315\ : CascadeBuf
    port map (
            O => \N__10699\,
            I => \N__10693\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__10696\,
            I => \N__10690\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__10693\,
            I => \N__10687\
        );

    \I__1312\ : CascadeBuf
    port map (
            O => \N__10690\,
            I => \N__10684\
        );

    \I__1311\ : CascadeBuf
    port map (
            O => \N__10687\,
            I => \N__10681\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__10684\,
            I => \N__10678\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__10681\,
            I => \N__10675\
        );

    \I__1308\ : CascadeBuf
    port map (
            O => \N__10678\,
            I => \N__10672\
        );

    \I__1307\ : CascadeBuf
    port map (
            O => \N__10675\,
            I => \N__10669\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__10672\,
            I => \N__10666\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__10669\,
            I => \N__10663\
        );

    \I__1304\ : CascadeBuf
    port map (
            O => \N__10666\,
            I => \N__10660\
        );

    \I__1303\ : CascadeBuf
    port map (
            O => \N__10663\,
            I => \N__10657\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__10660\,
            I => \N__10654\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__10657\,
            I => \N__10651\
        );

    \I__1300\ : CascadeBuf
    port map (
            O => \N__10654\,
            I => \N__10648\
        );

    \I__1299\ : CascadeBuf
    port map (
            O => \N__10651\,
            I => \N__10645\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__10648\,
            I => \N__10642\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__10645\,
            I => \N__10639\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10636\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10633\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__10636\,
            I => \N__10629\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__10633\,
            I => \N__10626\
        );

    \I__1292\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10622\
        );

    \I__1291\ : Span4Mux_s3_v
    port map (
            O => \N__10629\,
            I => \N__10619\
        );

    \I__1290\ : Span4Mux_s2_v
    port map (
            O => \N__10626\,
            I => \N__10616\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__10625\,
            I => \N__10613\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__10622\,
            I => \N__10610\
        );

    \I__1287\ : Span4Mux_h
    port map (
            O => \N__10619\,
            I => \N__10607\
        );

    \I__1286\ : Sp12to4
    port map (
            O => \N__10616\,
            I => \N__10604\
        );

    \I__1285\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10601\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__10610\,
            I => \N__10598\
        );

    \I__1283\ : Sp12to4
    port map (
            O => \N__10607\,
            I => \N__10593\
        );

    \I__1282\ : Span12Mux_h
    port map (
            O => \N__10604\,
            I => \N__10593\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__10601\,
            I => \RX_ADDR_8\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__10598\,
            I => \RX_ADDR_8\
        );

    \I__1279\ : Odrv12
    port map (
            O => \N__10593\,
            I => \RX_ADDR_8\
        );

    \I__1278\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10583\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__10583\,
            I => \N__10580\
        );

    \I__1276\ : Odrv12
    port map (
            O => \N__10580\,
            I => \receive_module.n127\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__10577\,
            I => \N__10574\
        );

    \I__1274\ : CascadeBuf
    port map (
            O => \N__10574\,
            I => \N__10570\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__10573\,
            I => \N__10567\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__10570\,
            I => \N__10564\
        );

    \I__1271\ : CascadeBuf
    port map (
            O => \N__10567\,
            I => \N__10561\
        );

    \I__1270\ : CascadeBuf
    port map (
            O => \N__10564\,
            I => \N__10558\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__10561\,
            I => \N__10555\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__10558\,
            I => \N__10552\
        );

    \I__1267\ : CascadeBuf
    port map (
            O => \N__10555\,
            I => \N__10549\
        );

    \I__1266\ : CascadeBuf
    port map (
            O => \N__10552\,
            I => \N__10546\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__10549\,
            I => \N__10543\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__10546\,
            I => \N__10540\
        );

    \I__1263\ : CascadeBuf
    port map (
            O => \N__10543\,
            I => \N__10537\
        );

    \I__1262\ : CascadeBuf
    port map (
            O => \N__10540\,
            I => \N__10534\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__10537\,
            I => \N__10531\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__10534\,
            I => \N__10528\
        );

    \I__1259\ : CascadeBuf
    port map (
            O => \N__10531\,
            I => \N__10525\
        );

    \I__1258\ : CascadeBuf
    port map (
            O => \N__10528\,
            I => \N__10522\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__10525\,
            I => \N__10519\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__10522\,
            I => \N__10516\
        );

    \I__1255\ : CascadeBuf
    port map (
            O => \N__10519\,
            I => \N__10513\
        );

    \I__1254\ : CascadeBuf
    port map (
            O => \N__10516\,
            I => \N__10510\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__10513\,
            I => \N__10507\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__10510\,
            I => \N__10504\
        );

    \I__1251\ : CascadeBuf
    port map (
            O => \N__10507\,
            I => \N__10501\
        );

    \I__1250\ : CascadeBuf
    port map (
            O => \N__10504\,
            I => \N__10498\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__10501\,
            I => \N__10495\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__10498\,
            I => \N__10492\
        );

    \I__1247\ : CascadeBuf
    port map (
            O => \N__10495\,
            I => \N__10489\
        );

    \I__1246\ : CascadeBuf
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__10489\,
            I => \N__10483\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__10486\,
            I => \N__10480\
        );

    \I__1243\ : CascadeBuf
    port map (
            O => \N__10483\,
            I => \N__10477\
        );

    \I__1242\ : CascadeBuf
    port map (
            O => \N__10480\,
            I => \N__10474\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__10477\,
            I => \N__10471\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__10474\,
            I => \N__10468\
        );

    \I__1239\ : CascadeBuf
    port map (
            O => \N__10471\,
            I => \N__10465\
        );

    \I__1238\ : CascadeBuf
    port map (
            O => \N__10468\,
            I => \N__10462\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__10465\,
            I => \N__10459\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__10462\,
            I => \N__10456\
        );

    \I__1235\ : CascadeBuf
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__1234\ : CascadeBuf
    port map (
            O => \N__10456\,
            I => \N__10450\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__10453\,
            I => \N__10447\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__10450\,
            I => \N__10444\
        );

    \I__1231\ : CascadeBuf
    port map (
            O => \N__10447\,
            I => \N__10441\
        );

    \I__1230\ : CascadeBuf
    port map (
            O => \N__10444\,
            I => \N__10438\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__10441\,
            I => \N__10435\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__10438\,
            I => \N__10432\
        );

    \I__1227\ : CascadeBuf
    port map (
            O => \N__10435\,
            I => \N__10429\
        );

    \I__1226\ : CascadeBuf
    port map (
            O => \N__10432\,
            I => \N__10426\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__10429\,
            I => \N__10423\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__10426\,
            I => \N__10420\
        );

    \I__1223\ : CascadeBuf
    port map (
            O => \N__10423\,
            I => \N__10417\
        );

    \I__1222\ : CascadeBuf
    port map (
            O => \N__10420\,
            I => \N__10414\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__10417\,
            I => \N__10411\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__10414\,
            I => \N__10408\
        );

    \I__1219\ : CascadeBuf
    port map (
            O => \N__10411\,
            I => \N__10405\
        );

    \I__1218\ : CascadeBuf
    port map (
            O => \N__10408\,
            I => \N__10402\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__10405\,
            I => \N__10399\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__10402\,
            I => \N__10396\
        );

    \I__1215\ : CascadeBuf
    port map (
            O => \N__10399\,
            I => \N__10393\
        );

    \I__1214\ : InMux
    port map (
            O => \N__10396\,
            I => \N__10390\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__10393\,
            I => \N__10387\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10390\,
            I => \N__10384\
        );

    \I__1211\ : InMux
    port map (
            O => \N__10387\,
            I => \N__10381\
        );

    \I__1210\ : Span4Mux_s2_v
    port map (
            O => \N__10384\,
            I => \N__10378\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__10381\,
            I => \N__10375\
        );

    \I__1208\ : Span4Mux_h
    port map (
            O => \N__10378\,
            I => \N__10372\
        );

    \I__1207\ : Span4Mux_s2_v
    port map (
            O => \N__10375\,
            I => \N__10368\
        );

    \I__1206\ : Span4Mux_h
    port map (
            O => \N__10372\,
            I => \N__10365\
        );

    \I__1205\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10362\
        );

    \I__1204\ : Span4Mux_h
    port map (
            O => \N__10368\,
            I => \N__10357\
        );

    \I__1203\ : Span4Mux_h
    port map (
            O => \N__10365\,
            I => \N__10357\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__10362\,
            I => \N__10353\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__10357\,
            I => \N__10350\
        );

    \I__1200\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10347\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__10353\,
            I => \N__10344\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__10350\,
            I => \N__10341\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__10347\,
            I => \RX_ADDR_9\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__10344\,
            I => \RX_ADDR_9\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__10341\,
            I => \RX_ADDR_9\
        );

    \I__1194\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1192\ : Odrv12
    port map (
            O => \N__10328\,
            I => \receive_module.n136\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__10325\,
            I => \N__10321\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__10324\,
            I => \N__10318\
        );

    \I__1189\ : CascadeBuf
    port map (
            O => \N__10321\,
            I => \N__10315\
        );

    \I__1188\ : CascadeBuf
    port map (
            O => \N__10318\,
            I => \N__10312\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__10315\,
            I => \N__10309\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__10312\,
            I => \N__10306\
        );

    \I__1185\ : CascadeBuf
    port map (
            O => \N__10309\,
            I => \N__10303\
        );

    \I__1184\ : CascadeBuf
    port map (
            O => \N__10306\,
            I => \N__10300\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__10303\,
            I => \N__10297\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__10300\,
            I => \N__10294\
        );

    \I__1181\ : CascadeBuf
    port map (
            O => \N__10297\,
            I => \N__10291\
        );

    \I__1180\ : CascadeBuf
    port map (
            O => \N__10294\,
            I => \N__10288\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__10291\,
            I => \N__10285\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__10288\,
            I => \N__10282\
        );

    \I__1177\ : CascadeBuf
    port map (
            O => \N__10285\,
            I => \N__10279\
        );

    \I__1176\ : CascadeBuf
    port map (
            O => \N__10282\,
            I => \N__10276\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__10279\,
            I => \N__10273\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__10276\,
            I => \N__10270\
        );

    \I__1173\ : CascadeBuf
    port map (
            O => \N__10273\,
            I => \N__10267\
        );

    \I__1172\ : CascadeBuf
    port map (
            O => \N__10270\,
            I => \N__10264\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__10267\,
            I => \N__10261\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__10264\,
            I => \N__10258\
        );

    \I__1169\ : CascadeBuf
    port map (
            O => \N__10261\,
            I => \N__10255\
        );

    \I__1168\ : CascadeBuf
    port map (
            O => \N__10258\,
            I => \N__10252\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__10255\,
            I => \N__10249\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__10252\,
            I => \N__10246\
        );

    \I__1165\ : CascadeBuf
    port map (
            O => \N__10249\,
            I => \N__10243\
        );

    \I__1164\ : CascadeBuf
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__10243\,
            I => \N__10237\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__10240\,
            I => \N__10234\
        );

    \I__1161\ : CascadeBuf
    port map (
            O => \N__10237\,
            I => \N__10231\
        );

    \I__1160\ : CascadeBuf
    port map (
            O => \N__10234\,
            I => \N__10228\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__10228\,
            I => \N__10222\
        );

    \I__1157\ : CascadeBuf
    port map (
            O => \N__10225\,
            I => \N__10219\
        );

    \I__1156\ : CascadeBuf
    port map (
            O => \N__10222\,
            I => \N__10216\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__10219\,
            I => \N__10213\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__10216\,
            I => \N__10210\
        );

    \I__1153\ : CascadeBuf
    port map (
            O => \N__10213\,
            I => \N__10207\
        );

    \I__1152\ : CascadeBuf
    port map (
            O => \N__10210\,
            I => \N__10204\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__10207\,
            I => \N__10201\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__10204\,
            I => \N__10198\
        );

    \I__1149\ : CascadeBuf
    port map (
            O => \N__10201\,
            I => \N__10195\
        );

    \I__1148\ : CascadeBuf
    port map (
            O => \N__10198\,
            I => \N__10192\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__10195\,
            I => \N__10189\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__10192\,
            I => \N__10186\
        );

    \I__1145\ : CascadeBuf
    port map (
            O => \N__10189\,
            I => \N__10183\
        );

    \I__1144\ : CascadeBuf
    port map (
            O => \N__10186\,
            I => \N__10180\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__10183\,
            I => \N__10177\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__10180\,
            I => \N__10174\
        );

    \I__1141\ : CascadeBuf
    port map (
            O => \N__10177\,
            I => \N__10171\
        );

    \I__1140\ : CascadeBuf
    port map (
            O => \N__10174\,
            I => \N__10168\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__10168\,
            I => \N__10162\
        );

    \I__1137\ : CascadeBuf
    port map (
            O => \N__10165\,
            I => \N__10159\
        );

    \I__1136\ : CascadeBuf
    port map (
            O => \N__10162\,
            I => \N__10156\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__10159\,
            I => \N__10153\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__10156\,
            I => \N__10150\
        );

    \I__1133\ : CascadeBuf
    port map (
            O => \N__10153\,
            I => \N__10147\
        );

    \I__1132\ : CascadeBuf
    port map (
            O => \N__10150\,
            I => \N__10144\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__10147\,
            I => \N__10141\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__10144\,
            I => \N__10138\
        );

    \I__1129\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10135\
        );

    \I__1128\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10132\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__10135\,
            I => \N__10129\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__10132\,
            I => \N__10125\
        );

    \I__1125\ : Span4Mux_s1_v
    port map (
            O => \N__10129\,
            I => \N__10122\
        );

    \I__1124\ : InMux
    port map (
            O => \N__10128\,
            I => \N__10119\
        );

    \I__1123\ : Span4Mux_s2_v
    port map (
            O => \N__10125\,
            I => \N__10116\
        );

    \I__1122\ : Span4Mux_h
    port map (
            O => \N__10122\,
            I => \N__10113\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__10119\,
            I => \N__10110\
        );

    \I__1120\ : Span4Mux_h
    port map (
            O => \N__10116\,
            I => \N__10107\
        );

    \I__1119\ : Sp12to4
    port map (
            O => \N__10113\,
            I => \N__10103\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__10110\,
            I => \N__10100\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__10107\,
            I => \N__10097\
        );

    \I__1116\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10094\
        );

    \I__1115\ : Span12Mux_v
    port map (
            O => \N__10103\,
            I => \N__10091\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__10100\,
            I => \N__10086\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__10097\,
            I => \N__10086\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__10094\,
            I => \RX_ADDR_0\
        );

    \I__1111\ : Odrv12
    port map (
            O => \N__10091\,
            I => \RX_ADDR_0\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__10086\,
            I => \RX_ADDR_0\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__1108\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__1106\ : Odrv12
    port map (
            O => \N__10070\,
            I => \receive_module.n135\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__10067\,
            I => \N__10063\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__10066\,
            I => \N__10060\
        );

    \I__1103\ : CascadeBuf
    port map (
            O => \N__10063\,
            I => \N__10057\
        );

    \I__1102\ : CascadeBuf
    port map (
            O => \N__10060\,
            I => \N__10054\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__10057\,
            I => \N__10051\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__10054\,
            I => \N__10048\
        );

    \I__1099\ : CascadeBuf
    port map (
            O => \N__10051\,
            I => \N__10045\
        );

    \I__1098\ : CascadeBuf
    port map (
            O => \N__10048\,
            I => \N__10042\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__10045\,
            I => \N__10039\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__10042\,
            I => \N__10036\
        );

    \I__1095\ : CascadeBuf
    port map (
            O => \N__10039\,
            I => \N__10033\
        );

    \I__1094\ : CascadeBuf
    port map (
            O => \N__10036\,
            I => \N__10030\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__10033\,
            I => \N__10027\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__10030\,
            I => \N__10024\
        );

    \I__1091\ : CascadeBuf
    port map (
            O => \N__10027\,
            I => \N__10021\
        );

    \I__1090\ : CascadeBuf
    port map (
            O => \N__10024\,
            I => \N__10018\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__10021\,
            I => \N__10015\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__10018\,
            I => \N__10012\
        );

    \I__1087\ : CascadeBuf
    port map (
            O => \N__10015\,
            I => \N__10009\
        );

    \I__1086\ : CascadeBuf
    port map (
            O => \N__10012\,
            I => \N__10006\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__10009\,
            I => \N__10003\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__10006\,
            I => \N__10000\
        );

    \I__1083\ : CascadeBuf
    port map (
            O => \N__10003\,
            I => \N__9997\
        );

    \I__1082\ : CascadeBuf
    port map (
            O => \N__10000\,
            I => \N__9994\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__9997\,
            I => \N__9991\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__9994\,
            I => \N__9988\
        );

    \I__1079\ : CascadeBuf
    port map (
            O => \N__9991\,
            I => \N__9985\
        );

    \I__1078\ : CascadeBuf
    port map (
            O => \N__9988\,
            I => \N__9982\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__9985\,
            I => \N__9979\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__9982\,
            I => \N__9976\
        );

    \I__1075\ : CascadeBuf
    port map (
            O => \N__9979\,
            I => \N__9973\
        );

    \I__1074\ : CascadeBuf
    port map (
            O => \N__9976\,
            I => \N__9970\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__9973\,
            I => \N__9967\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__9970\,
            I => \N__9964\
        );

    \I__1071\ : CascadeBuf
    port map (
            O => \N__9967\,
            I => \N__9961\
        );

    \I__1070\ : CascadeBuf
    port map (
            O => \N__9964\,
            I => \N__9958\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__9961\,
            I => \N__9955\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__9958\,
            I => \N__9952\
        );

    \I__1067\ : CascadeBuf
    port map (
            O => \N__9955\,
            I => \N__9949\
        );

    \I__1066\ : CascadeBuf
    port map (
            O => \N__9952\,
            I => \N__9946\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__9949\,
            I => \N__9943\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__9946\,
            I => \N__9940\
        );

    \I__1063\ : CascadeBuf
    port map (
            O => \N__9943\,
            I => \N__9937\
        );

    \I__1062\ : CascadeBuf
    port map (
            O => \N__9940\,
            I => \N__9934\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__9937\,
            I => \N__9931\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__9934\,
            I => \N__9928\
        );

    \I__1059\ : CascadeBuf
    port map (
            O => \N__9931\,
            I => \N__9925\
        );

    \I__1058\ : CascadeBuf
    port map (
            O => \N__9928\,
            I => \N__9922\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__9925\,
            I => \N__9919\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__9922\,
            I => \N__9916\
        );

    \I__1055\ : CascadeBuf
    port map (
            O => \N__9919\,
            I => \N__9913\
        );

    \I__1054\ : CascadeBuf
    port map (
            O => \N__9916\,
            I => \N__9910\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__9913\,
            I => \N__9907\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__9910\,
            I => \N__9904\
        );

    \I__1051\ : CascadeBuf
    port map (
            O => \N__9907\,
            I => \N__9901\
        );

    \I__1050\ : CascadeBuf
    port map (
            O => \N__9904\,
            I => \N__9898\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__9901\,
            I => \N__9895\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__9898\,
            I => \N__9892\
        );

    \I__1047\ : CascadeBuf
    port map (
            O => \N__9895\,
            I => \N__9889\
        );

    \I__1046\ : CascadeBuf
    port map (
            O => \N__9892\,
            I => \N__9886\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__9889\,
            I => \N__9883\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__9886\,
            I => \N__9880\
        );

    \I__1043\ : InMux
    port map (
            O => \N__9883\,
            I => \N__9877\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9874\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__9877\,
            I => \N__9871\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__9874\,
            I => \N__9867\
        );

    \I__1039\ : Span4Mux_s2_v
    port map (
            O => \N__9871\,
            I => \N__9864\
        );

    \I__1038\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9861\
        );

    \I__1037\ : Span12Mux_s1_v
    port map (
            O => \N__9867\,
            I => \N__9858\
        );

    \I__1036\ : Span4Mux_h
    port map (
            O => \N__9864\,
            I => \N__9855\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__9861\,
            I => \N__9852\
        );

    \I__1034\ : Span12Mux_v
    port map (
            O => \N__9858\,
            I => \N__9848\
        );

    \I__1033\ : Span4Mux_v
    port map (
            O => \N__9855\,
            I => \N__9845\
        );

    \I__1032\ : Span12Mux_v
    port map (
            O => \N__9852\,
            I => \N__9842\
        );

    \I__1031\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9839\
        );

    \I__1030\ : Span12Mux_h
    port map (
            O => \N__9848\,
            I => \N__9836\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__9845\,
            I => \N__9833\
        );

    \I__1028\ : Odrv12
    port map (
            O => \N__9842\,
            I => \RX_ADDR_1\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9839\,
            I => \RX_ADDR_1\
        );

    \I__1026\ : Odrv12
    port map (
            O => \N__9836\,
            I => \RX_ADDR_1\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__9833\,
            I => \RX_ADDR_1\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9821\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__1022\ : Span12Mux_v
    port map (
            O => \N__9818\,
            I => \N__9815\
        );

    \I__1021\ : Odrv12
    port map (
            O => \N__9815\,
            I => \line_buffer.n593\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9812\,
            I => \N__9809\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__9809\,
            I => \N__9806\
        );

    \I__1018\ : Span12Mux_v
    port map (
            O => \N__9806\,
            I => \N__9803\
        );

    \I__1017\ : Odrv12
    port map (
            O => \N__9803\,
            I => \line_buffer.n585\
        );

    \I__1016\ : InMux
    port map (
            O => \N__9800\,
            I => \transmit_module.video_signal_controller.n3133\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9797\,
            I => \transmit_module.video_signal_controller.n3134\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9794\,
            I => \transmit_module.video_signal_controller.n3135\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9788\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__9788\,
            I => \transmit_module.Y_DELTA_PATTERN_2\
        );

    \I__1011\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9782\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9782\,
            I => \transmit_module.Y_DELTA_PATTERN_3\
        );

    \I__1009\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9776\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__9776\,
            I => \transmit_module.Y_DELTA_PATTERN_5\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9770\,
            I => \transmit_module.Y_DELTA_PATTERN_4\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9767\,
            I => \bfn_12_15_0_\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9764\,
            I => \transmit_module.video_signal_controller.n3125\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9761\,
            I => \transmit_module.video_signal_controller.n3126\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9758\,
            I => \transmit_module.video_signal_controller.n3127\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9755\,
            I => \transmit_module.video_signal_controller.n3128\
        );

    \I__1000\ : InMux
    port map (
            O => \N__9752\,
            I => \transmit_module.video_signal_controller.n3129\
        );

    \I__999\ : InMux
    port map (
            O => \N__9749\,
            I => \transmit_module.video_signal_controller.n3130\
        );

    \I__998\ : InMux
    port map (
            O => \N__9746\,
            I => \transmit_module.video_signal_controller.n3131\
        );

    \I__997\ : InMux
    port map (
            O => \N__9743\,
            I => \bfn_12_16_0_\
        );

    \I__996\ : InMux
    port map (
            O => \N__9740\,
            I => \receive_module.n3102\
        );

    \I__995\ : InMux
    port map (
            O => \N__9737\,
            I => \receive_module.n3103\
        );

    \I__994\ : CEMux
    port map (
            O => \N__9734\,
            I => \N__9731\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__992\ : Span4Mux_h
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__9725\,
            I => \receive_module.n3632\
        );

    \I__990\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__9719\,
            I => \transmit_module.Y_DELTA_PATTERN_53\
        );

    \I__988\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__9713\,
            I => \transmit_module.Y_DELTA_PATTERN_52\
        );

    \I__986\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9707\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__9707\,
            I => \transmit_module.Y_DELTA_PATTERN_56\
        );

    \I__984\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__9701\,
            I => \transmit_module.Y_DELTA_PATTERN_55\
        );

    \I__982\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9695\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__9695\,
            I => \transmit_module.Y_DELTA_PATTERN_54\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__9692\,
            I => \transmit_module.video_signal_controller.n3629_cascade_\
        );

    \I__979\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__9686\,
            I => \transmit_module.video_signal_controller.n2901\
        );

    \I__977\ : InMux
    port map (
            O => \N__9683\,
            I => \receive_module.n3093\
        );

    \I__976\ : InMux
    port map (
            O => \N__9680\,
            I => \receive_module.n3094\
        );

    \I__975\ : InMux
    port map (
            O => \N__9677\,
            I => \receive_module.n3095\
        );

    \I__974\ : InMux
    port map (
            O => \N__9674\,
            I => \receive_module.n3096\
        );

    \I__973\ : InMux
    port map (
            O => \N__9671\,
            I => \receive_module.n3097\
        );

    \I__972\ : InMux
    port map (
            O => \N__9668\,
            I => \bfn_12_12_0_\
        );

    \I__971\ : InMux
    port map (
            O => \N__9665\,
            I => \receive_module.n3099\
        );

    \I__970\ : InMux
    port map (
            O => \N__9662\,
            I => \receive_module.n3100\
        );

    \I__969\ : InMux
    port map (
            O => \N__9659\,
            I => \receive_module.n3101\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__9656\,
            I => \receive_module.rx_counter.n4_cascade_\
        );

    \I__967\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9650\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9650\,
            I => \receive_module.rx_counter.n3400\
        );

    \I__965\ : SRMux
    port map (
            O => \N__9647\,
            I => \N__9644\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__963\ : Span4Mux_v
    port map (
            O => \N__9641\,
            I => \N__9637\
        );

    \I__962\ : SRMux
    port map (
            O => \N__9640\,
            I => \N__9633\
        );

    \I__961\ : Span4Mux_v
    port map (
            O => \N__9637\,
            I => \N__9630\
        );

    \I__960\ : SRMux
    port map (
            O => \N__9636\,
            I => \N__9627\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__9633\,
            I => \N__9624\
        );

    \I__958\ : Span4Mux_v
    port map (
            O => \N__9630\,
            I => \N__9619\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__9627\,
            I => \N__9619\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__9624\,
            I => \N__9613\
        );

    \I__955\ : Span4Mux_v
    port map (
            O => \N__9619\,
            I => \N__9613\
        );

    \I__954\ : SRMux
    port map (
            O => \N__9618\,
            I => \N__9610\
        );

    \I__953\ : Sp12to4
    port map (
            O => \N__9613\,
            I => \N__9605\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9610\,
            I => \N__9605\
        );

    \I__951\ : Odrv12
    port map (
            O => \N__9605\,
            I => \line_buffer.n565\
        );

    \I__950\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9597\
        );

    \I__949\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9592\
        );

    \I__948\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9592\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9597\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__9592\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__945\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9582\
        );

    \I__944\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9577\
        );

    \I__943\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9577\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__9582\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__9577\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__940\ : InMux
    port map (
            O => \N__9572\,
            I => \N__9567\
        );

    \I__939\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9562\
        );

    \I__938\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9562\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9567\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__9562\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__935\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9552\
        );

    \I__934\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9547\
        );

    \I__933\ : InMux
    port map (
            O => \N__9555\,
            I => \N__9547\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__9552\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__9547\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__9542\,
            I => \receive_module.rx_counter.n6_cascade_\
        );

    \I__929\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9534\
        );

    \I__928\ : InMux
    port map (
            O => \N__9538\,
            I => \N__9529\
        );

    \I__927\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9529\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9534\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__9529\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__924\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9521\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__9521\,
            I => \receive_module.rx_counter.n3385\
        );

    \I__922\ : InMux
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__920\ : Odrv4
    port map (
            O => \N__9512\,
            I => \receive_module.rx_counter.old_HS\
        );

    \I__919\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9505\
        );

    \I__918\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9501\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__9505\,
            I => \N__9498\
        );

    \I__916\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9495\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__9501\,
            I => \TVP_HSYNC_buff\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__9498\,
            I => \TVP_HSYNC_buff\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__9495\,
            I => \TVP_HSYNC_buff\
        );

    \I__912\ : InMux
    port map (
            O => \N__9488\,
            I => \bfn_12_11_0_\
        );

    \I__911\ : InMux
    port map (
            O => \N__9485\,
            I => \receive_module.n3091\
        );

    \I__910\ : InMux
    port map (
            O => \N__9482\,
            I => \receive_module.n3092\
        );

    \I__909\ : IoInMux
    port map (
            O => \N__9479\,
            I => \N__9476\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__9476\,
            I => \N__9473\
        );

    \I__907\ : Span4Mux_s2_h
    port map (
            O => \N__9473\,
            I => \N__9470\
        );

    \I__906\ : Span4Mux_h
    port map (
            O => \N__9470\,
            I => \N__9466\
        );

    \I__905\ : InMux
    port map (
            O => \N__9469\,
            I => \N__9463\
        );

    \I__904\ : Span4Mux_h
    port map (
            O => \N__9466\,
            I => \N__9458\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__9463\,
            I => \N__9458\
        );

    \I__902\ : Span4Mux_h
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__901\ : Span4Mux_v
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__9452\,
            I => \DEBUG_c_0_c\
        );

    \I__899\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__9446\,
            I => \TVP_VSYNC_buff_I_0.BUFFER_0_0\
        );

    \I__897\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9439\
        );

    \I__896\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9436\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__9439\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__9436\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__9431\,
            I => \N__9427\
        );

    \I__892\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9424\
        );

    \I__891\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9421\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__9424\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__9421\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__888\ : SRMux
    port map (
            O => \N__9416\,
            I => \N__9412\
        );

    \I__887\ : SRMux
    port map (
            O => \N__9415\,
            I => \N__9409\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__9412\,
            I => \N__9406\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__9409\,
            I => \N__9403\
        );

    \I__884\ : Sp12to4
    port map (
            O => \N__9406\,
            I => \N__9400\
        );

    \I__883\ : Span4Mux_h
    port map (
            O => \N__9403\,
            I => \N__9397\
        );

    \I__882\ : Odrv12
    port map (
            O => \N__9400\,
            I => \receive_module.rx_counter.n3630\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__9397\,
            I => \receive_module.rx_counter.n3630\
        );

    \I__880\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9389\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__9389\,
            I => \N__9386\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__9386\,
            I => \TVP_VSYNC_buff_I_0.BUFFER_1_0\
        );

    \I__877\ : SRMux
    port map (
            O => \N__9383\,
            I => \N__9379\
        );

    \I__876\ : SRMux
    port map (
            O => \N__9382\,
            I => \N__9376\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__9379\,
            I => \N__9370\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__9376\,
            I => \N__9370\
        );

    \I__873\ : SRMux
    port map (
            O => \N__9375\,
            I => \N__9367\
        );

    \I__872\ : Span4Mux_v
    port map (
            O => \N__9370\,
            I => \N__9362\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__9367\,
            I => \N__9362\
        );

    \I__870\ : Span4Mux_h
    port map (
            O => \N__9362\,
            I => \N__9358\
        );

    \I__869\ : SRMux
    port map (
            O => \N__9361\,
            I => \N__9355\
        );

    \I__868\ : Span4Mux_v
    port map (
            O => \N__9358\,
            I => \N__9352\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__9355\,
            I => \N__9349\
        );

    \I__866\ : Span4Mux_v
    port map (
            O => \N__9352\,
            I => \N__9346\
        );

    \I__865\ : Span4Mux_v
    port map (
            O => \N__9349\,
            I => \N__9343\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__9346\,
            I => \N__9340\
        );

    \I__863\ : Sp12to4
    port map (
            O => \N__9343\,
            I => \N__9337\
        );

    \I__862\ : Span4Mux_v
    port map (
            O => \N__9340\,
            I => \N__9334\
        );

    \I__861\ : Span12Mux_h
    port map (
            O => \N__9337\,
            I => \N__9331\
        );

    \I__860\ : Odrv4
    port map (
            O => \N__9334\,
            I => \line_buffer.n467\
        );

    \I__859\ : Odrv12
    port map (
            O => \N__9331\,
            I => \line_buffer.n467\
        );

    \I__858\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__9323\,
            I => \transmit_module.Y_DELTA_PATTERN_43\
        );

    \I__856\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__854\ : Odrv12
    port map (
            O => \N__9314\,
            I => \transmit_module.Y_DELTA_PATTERN_59\
        );

    \I__853\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9308\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__9308\,
            I => \transmit_module.Y_DELTA_PATTERN_45\
        );

    \I__851\ : InMux
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__9302\,
            I => \transmit_module.Y_DELTA_PATTERN_44\
        );

    \I__849\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__9293\,
            I => \transmit_module.Y_DELTA_PATTERN_47\
        );

    \I__846\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__9287\,
            I => \transmit_module.Y_DELTA_PATTERN_46\
        );

    \I__844\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9281\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__9281\,
            I => \transmit_module.Y_DELTA_PATTERN_61\
        );

    \I__842\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__9275\,
            I => \transmit_module.Y_DELTA_PATTERN_60\
        );

    \I__840\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__9269\,
            I => \transmit_module.Y_DELTA_PATTERN_77\
        );

    \I__838\ : InMux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__9263\,
            I => \transmit_module.Y_DELTA_PATTERN_76\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__835\ : CascadeBuf
    port map (
            O => \N__9257\,
            I => \N__9253\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__9256\,
            I => \N__9250\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__9253\,
            I => \N__9247\
        );

    \I__832\ : CascadeBuf
    port map (
            O => \N__9250\,
            I => \N__9244\
        );

    \I__831\ : CascadeBuf
    port map (
            O => \N__9247\,
            I => \N__9241\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__9244\,
            I => \N__9238\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__9241\,
            I => \N__9235\
        );

    \I__828\ : CascadeBuf
    port map (
            O => \N__9238\,
            I => \N__9232\
        );

    \I__827\ : CascadeBuf
    port map (
            O => \N__9235\,
            I => \N__9229\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__9232\,
            I => \N__9226\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__9229\,
            I => \N__9223\
        );

    \I__824\ : CascadeBuf
    port map (
            O => \N__9226\,
            I => \N__9220\
        );

    \I__823\ : CascadeBuf
    port map (
            O => \N__9223\,
            I => \N__9217\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__9220\,
            I => \N__9214\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__9217\,
            I => \N__9211\
        );

    \I__820\ : CascadeBuf
    port map (
            O => \N__9214\,
            I => \N__9208\
        );

    \I__819\ : CascadeBuf
    port map (
            O => \N__9211\,
            I => \N__9205\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__9208\,
            I => \N__9202\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__9205\,
            I => \N__9199\
        );

    \I__816\ : CascadeBuf
    port map (
            O => \N__9202\,
            I => \N__9196\
        );

    \I__815\ : CascadeBuf
    port map (
            O => \N__9199\,
            I => \N__9193\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__9196\,
            I => \N__9190\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__9193\,
            I => \N__9187\
        );

    \I__812\ : CascadeBuf
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__811\ : CascadeBuf
    port map (
            O => \N__9187\,
            I => \N__9181\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__9184\,
            I => \N__9178\
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__9181\,
            I => \N__9175\
        );

    \I__808\ : CascadeBuf
    port map (
            O => \N__9178\,
            I => \N__9172\
        );

    \I__807\ : CascadeBuf
    port map (
            O => \N__9175\,
            I => \N__9169\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__9172\,
            I => \N__9166\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__9169\,
            I => \N__9163\
        );

    \I__804\ : CascadeBuf
    port map (
            O => \N__9166\,
            I => \N__9160\
        );

    \I__803\ : CascadeBuf
    port map (
            O => \N__9163\,
            I => \N__9157\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__9160\,
            I => \N__9154\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__9157\,
            I => \N__9151\
        );

    \I__800\ : CascadeBuf
    port map (
            O => \N__9154\,
            I => \N__9148\
        );

    \I__799\ : CascadeBuf
    port map (
            O => \N__9151\,
            I => \N__9145\
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__9148\,
            I => \N__9142\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__9145\,
            I => \N__9139\
        );

    \I__796\ : CascadeBuf
    port map (
            O => \N__9142\,
            I => \N__9136\
        );

    \I__795\ : CascadeBuf
    port map (
            O => \N__9139\,
            I => \N__9133\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__9136\,
            I => \N__9130\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__9133\,
            I => \N__9127\
        );

    \I__792\ : CascadeBuf
    port map (
            O => \N__9130\,
            I => \N__9124\
        );

    \I__791\ : CascadeBuf
    port map (
            O => \N__9127\,
            I => \N__9121\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__9124\,
            I => \N__9118\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__9121\,
            I => \N__9115\
        );

    \I__788\ : CascadeBuf
    port map (
            O => \N__9118\,
            I => \N__9112\
        );

    \I__787\ : CascadeBuf
    port map (
            O => \N__9115\,
            I => \N__9109\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__9112\,
            I => \N__9106\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__9109\,
            I => \N__9103\
        );

    \I__784\ : CascadeBuf
    port map (
            O => \N__9106\,
            I => \N__9100\
        );

    \I__783\ : CascadeBuf
    port map (
            O => \N__9103\,
            I => \N__9097\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__9100\,
            I => \N__9094\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__9097\,
            I => \N__9091\
        );

    \I__780\ : CascadeBuf
    port map (
            O => \N__9094\,
            I => \N__9088\
        );

    \I__779\ : CascadeBuf
    port map (
            O => \N__9091\,
            I => \N__9085\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__9088\,
            I => \N__9082\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__9085\,
            I => \N__9079\
        );

    \I__776\ : CascadeBuf
    port map (
            O => \N__9082\,
            I => \N__9076\
        );

    \I__775\ : InMux
    port map (
            O => \N__9079\,
            I => \N__9073\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__9076\,
            I => \N__9070\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__9073\,
            I => \N__9067\
        );

    \I__772\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9064\
        );

    \I__771\ : Span12Mux_h
    port map (
            O => \N__9067\,
            I => \N__9061\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__9064\,
            I => \N__9058\
        );

    \I__769\ : Odrv12
    port map (
            O => \N__9061\,
            I => n24
        );

    \I__768\ : Odrv4
    port map (
            O => \N__9058\,
            I => n24
        );

    \I__767\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__765\ : Span4Mux_h
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__9044\,
            I => \TVP_VIDEO_c_4\
        );

    \I__763\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__9038\,
            I => \transmit_module.Y_DELTA_PATTERN_99\
        );

    \I__761\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__9032\,
            I => \transmit_module.Y_DELTA_PATTERN_10\
        );

    \I__759\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__9026\,
            I => \transmit_module.Y_DELTA_PATTERN_9\
        );

    \I__757\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9020\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__9020\,
            I => \transmit_module.Y_DELTA_PATTERN_12\
        );

    \I__755\ : InMux
    port map (
            O => \N__9017\,
            I => \N__9014\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__9014\,
            I => \transmit_module.Y_DELTA_PATTERN_11\
        );

    \I__753\ : InMux
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__751\ : Odrv4
    port map (
            O => \N__9005\,
            I => \transmit_module.Y_DELTA_PATTERN_38\
        );

    \I__750\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__8999\,
            I => \transmit_module.Y_DELTA_PATTERN_40\
        );

    \I__748\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__8993\,
            I => \transmit_module.Y_DELTA_PATTERN_39\
        );

    \I__746\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8987\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8987\,
            I => \transmit_module.Y_DELTA_PATTERN_41\
        );

    \I__744\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__8981\,
            I => \transmit_module.Y_DELTA_PATTERN_42\
        );

    \I__742\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8975\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__8975\,
            I => \transmit_module.Y_DELTA_PATTERN_24\
        );

    \I__740\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__8969\,
            I => \transmit_module.Y_DELTA_PATTERN_23\
        );

    \I__738\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__8963\,
            I => \transmit_module.Y_DELTA_PATTERN_28\
        );

    \I__736\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8957\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__8957\,
            I => \transmit_module.Y_DELTA_PATTERN_27\
        );

    \I__734\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8951\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8951\,
            I => \transmit_module.Y_DELTA_PATTERN_13\
        );

    \I__732\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__8945\,
            I => \transmit_module.Y_DELTA_PATTERN_15\
        );

    \I__730\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__8939\,
            I => \transmit_module.Y_DELTA_PATTERN_14\
        );

    \I__728\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__8933\,
            I => \transmit_module.Y_DELTA_PATTERN_26\
        );

    \I__726\ : InMux
    port map (
            O => \N__8930\,
            I => \N__8927\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__8927\,
            I => \transmit_module.Y_DELTA_PATTERN_25\
        );

    \I__724\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__8921\,
            I => \transmit_module.Y_DELTA_PATTERN_8\
        );

    \I__722\ : InMux
    port map (
            O => \N__8918\,
            I => \N__8915\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__8915\,
            I => \transmit_module.Y_DELTA_PATTERN_50\
        );

    \I__720\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__8909\,
            I => \transmit_module.Y_DELTA_PATTERN_51\
        );

    \I__718\ : InMux
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__8903\,
            I => \transmit_module.Y_DELTA_PATTERN_58\
        );

    \I__716\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__8897\,
            I => \transmit_module.Y_DELTA_PATTERN_57\
        );

    \I__714\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__8891\,
            I => \transmit_module.Y_DELTA_PATTERN_22\
        );

    \I__712\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8885\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__8885\,
            I => \transmit_module.Y_DELTA_PATTERN_21\
        );

    \I__710\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8879\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__8879\,
            I => \receive_module.rx_counter.n9_adj_612\
        );

    \I__708\ : InMux
    port map (
            O => \N__8876\,
            I => \receive_module.rx_counter.n3147\
        );

    \I__707\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__8870\,
            I => \receive_module.rx_counter.n8_adj_611\
        );

    \I__705\ : InMux
    port map (
            O => \N__8867\,
            I => \receive_module.rx_counter.n3148\
        );

    \I__704\ : InMux
    port map (
            O => \N__8864\,
            I => \receive_module.rx_counter.n3149\
        );

    \I__703\ : InMux
    port map (
            O => \N__8861\,
            I => \receive_module.rx_counter.n3150\
        );

    \I__702\ : InMux
    port map (
            O => \N__8858\,
            I => \receive_module.rx_counter.n3151\
        );

    \I__701\ : InMux
    port map (
            O => \N__8855\,
            I => \receive_module.rx_counter.n3152\
        );

    \I__700\ : InMux
    port map (
            O => \N__8852\,
            I => \receive_module.rx_counter.n3153\
        );

    \I__699\ : InMux
    port map (
            O => \N__8849\,
            I => \bfn_11_10_0_\
        );

    \I__698\ : InMux
    port map (
            O => \N__8846\,
            I => \receive_module.rx_counter.n3155\
        );

    \I__697\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__8840\,
            I => \transmit_module.Y_DELTA_PATTERN_75\
        );

    \I__695\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__8834\,
            I => \transmit_module.Y_DELTA_PATTERN_62\
        );

    \I__693\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__8825\,
            I => \transmit_module.Y_DELTA_PATTERN_78\
        );

    \I__690\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__8819\,
            I => \tvp_video_buffer.BUFFER_0_2\
        );

    \I__688\ : IoInMux
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__686\ : Span12Mux_s6_v
    port map (
            O => \N__8810\,
            I => \N__8806\
        );

    \I__685\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8803\
        );

    \I__684\ : Odrv12
    port map (
            O => \N__8806\,
            I => \LED_c\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__8803\,
            I => \LED_c\
        );

    \I__682\ : IoInMux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__680\ : IoSpan4Mux
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__679\ : Span4Mux_s3_h
    port map (
            O => \N__8789\,
            I => \N__8785\
        );

    \I__678\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8782\
        );

    \I__677\ : Span4Mux_h
    port map (
            O => \N__8785\,
            I => \N__8779\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__8782\,
            I => \N__8776\
        );

    \I__675\ : Span4Mux_h
    port map (
            O => \N__8779\,
            I => \N__8771\
        );

    \I__674\ : Span4Mux_v
    port map (
            O => \N__8776\,
            I => \N__8771\
        );

    \I__673\ : Span4Mux_h
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__672\ : Span4Mux_h
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__8765\,
            I => \DEBUG_c_1_c\
        );

    \I__670\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__8759\,
            I => \tvp_hs_buffer.BUFFER_0_0\
        );

    \I__668\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8753\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__8753\,
            I => \tvp_hs_buffer.BUFFER_1_0\
        );

    \I__666\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__8747\,
            I => \receive_module.rx_counter.n10\
        );

    \I__664\ : InMux
    port map (
            O => \N__8744\,
            I => \bfn_11_9_0_\
        );

    \I__663\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__661\ : Odrv4
    port map (
            O => \N__8735\,
            I => \transmit_module.Y_DELTA_PATTERN_33\
        );

    \I__660\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8729\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__8729\,
            I => \transmit_module.Y_DELTA_PATTERN_29\
        );

    \I__658\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__8723\,
            I => \transmit_module.Y_DELTA_PATTERN_32\
        );

    \I__656\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__8717\,
            I => \transmit_module.Y_DELTA_PATTERN_31\
        );

    \I__654\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__8711\,
            I => \transmit_module.Y_DELTA_PATTERN_30\
        );

    \I__652\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__8705\,
            I => \transmit_module.Y_DELTA_PATTERN_74\
        );

    \I__650\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__8696\,
            I => \transmit_module.Y_DELTA_PATTERN_73\
        );

    \I__647\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__8690\,
            I => \transmit_module.Y_DELTA_PATTERN_65\
        );

    \I__645\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__8684\,
            I => \transmit_module.Y_DELTA_PATTERN_64\
        );

    \I__643\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__8678\,
            I => \transmit_module.Y_DELTA_PATTERN_63\
        );

    \I__641\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__8672\,
            I => \transmit_module.Y_DELTA_PATTERN_91\
        );

    \I__639\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__8666\,
            I => \transmit_module.Y_DELTA_PATTERN_93\
        );

    \I__637\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__8660\,
            I => \transmit_module.Y_DELTA_PATTERN_92\
        );

    \I__635\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__8654\,
            I => \transmit_module.Y_DELTA_PATTERN_94\
        );

    \I__633\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__8648\,
            I => \transmit_module.Y_DELTA_PATTERN_97\
        );

    \I__631\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__8642\,
            I => \transmit_module.Y_DELTA_PATTERN_98\
        );

    \I__629\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__8636\,
            I => \transmit_module.Y_DELTA_PATTERN_96\
        );

    \I__627\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__8630\,
            I => \transmit_module.Y_DELTA_PATTERN_95\
        );

    \I__625\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__623\ : IoSpan4Mux
    port map (
            O => \N__8621\,
            I => \N__8618\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__8618\,
            I => \TVP_VIDEO_c_2\
        );

    \I__621\ : SRMux
    port map (
            O => \N__8615\,
            I => \N__8610\
        );

    \I__620\ : SRMux
    port map (
            O => \N__8614\,
            I => \N__8607\
        );

    \I__619\ : SRMux
    port map (
            O => \N__8613\,
            I => \N__8604\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8600\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__8607\,
            I => \N__8595\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8595\
        );

    \I__615\ : SRMux
    port map (
            O => \N__8603\,
            I => \N__8592\
        );

    \I__614\ : Span4Mux_h
    port map (
            O => \N__8600\,
            I => \N__8589\
        );

    \I__613\ : Span4Mux_v
    port map (
            O => \N__8595\,
            I => \N__8584\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__8592\,
            I => \N__8584\
        );

    \I__611\ : Sp12to4
    port map (
            O => \N__8589\,
            I => \N__8581\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__8584\,
            I => \N__8578\
        );

    \I__609\ : Span12Mux_v
    port map (
            O => \N__8581\,
            I => \N__8575\
        );

    \I__608\ : Span4Mux_h
    port map (
            O => \N__8578\,
            I => \N__8572\
        );

    \I__607\ : Odrv12
    port map (
            O => \N__8575\,
            I => \line_buffer.n533\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__8572\,
            I => \line_buffer.n533\
        );

    \I__605\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__603\ : Span4Mux_h
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__8558\,
            I => \tvp_video_buffer.BUFFER_0_3\
        );

    \I__601\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__599\ : Span4Mux_v
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__598\ : Odrv4
    port map (
            O => \N__8546\,
            I => \transmit_module.Y_DELTA_PATTERN_82\
        );

    \I__597\ : InMux
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__595\ : Span4Mux_v
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__594\ : Odrv4
    port map (
            O => \N__8534\,
            I => \transmit_module.Y_DELTA_PATTERN_49\
        );

    \I__593\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__8528\,
            I => \transmit_module.Y_DELTA_PATTERN_84\
        );

    \I__591\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8522\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__8522\,
            I => \transmit_module.Y_DELTA_PATTERN_83\
        );

    \I__589\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__8516\,
            I => \transmit_module.Y_DELTA_PATTERN_85\
        );

    \I__587\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__8510\,
            I => \transmit_module.Y_DELTA_PATTERN_87\
        );

    \I__585\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__8504\,
            I => \transmit_module.Y_DELTA_PATTERN_86\
        );

    \I__583\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__8498\,
            I => \transmit_module.Y_DELTA_PATTERN_81\
        );

    \I__581\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__8492\,
            I => \transmit_module.Y_DELTA_PATTERN_80\
        );

    \I__579\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__8486\,
            I => \transmit_module.Y_DELTA_PATTERN_37\
        );

    \I__577\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__8480\,
            I => \transmit_module.Y_DELTA_PATTERN_79\
        );

    \I__575\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__8474\,
            I => \transmit_module.Y_DELTA_PATTERN_66\
        );

    \I__573\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__571\ : Span4Mux_v
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__8462\,
            I => \transmit_module.Y_DELTA_PATTERN_69\
        );

    \I__569\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8456\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__8456\,
            I => \transmit_module.Y_DELTA_PATTERN_68\
        );

    \I__567\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8450\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__8450\,
            I => \transmit_module.Y_DELTA_PATTERN_67\
        );

    \I__565\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__8444\,
            I => \transmit_module.Y_DELTA_PATTERN_48\
        );

    \I__563\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__8438\,
            I => \transmit_module.Y_DELTA_PATTERN_34\
        );

    \I__561\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8432\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__8429\,
            I => \transmit_module.Y_DELTA_PATTERN_72\
        );

    \I__558\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8423\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__8423\,
            I => \transmit_module.Y_DELTA_PATTERN_90\
        );

    \I__556\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8417\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__8417\,
            I => \transmit_module.Y_DELTA_PATTERN_89\
        );

    \I__554\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__8411\,
            I => \transmit_module.Y_DELTA_PATTERN_88\
        );

    \I__552\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__8402\,
            I => \transmit_module.Y_DELTA_PATTERN_36\
        );

    \I__549\ : IoInMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__8396\,
            I => \N__8392\
        );

    \I__547\ : IoInMux
    port map (
            O => \N__8395\,
            I => \N__8389\
        );

    \I__546\ : IoSpan4Mux
    port map (
            O => \N__8392\,
            I => \N__8386\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__8389\,
            I => \N__8383\
        );

    \I__544\ : Span4Mux_s3_v
    port map (
            O => \N__8386\,
            I => \N__8380\
        );

    \I__543\ : Span4Mux_s2_h
    port map (
            O => \N__8383\,
            I => \N__8377\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__8380\,
            I => \N__8374\
        );

    \I__541\ : Sp12to4
    port map (
            O => \N__8377\,
            I => \N__8371\
        );

    \I__540\ : Sp12to4
    port map (
            O => \N__8374\,
            I => \N__8366\
        );

    \I__539\ : Span12Mux_v
    port map (
            O => \N__8371\,
            I => \N__8366\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__8366\,
            I => \GB_BUFFER_DEBUG_c_2_c_THRU_CO\
        );

    \I__537\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8360\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__8360\,
            I => \transmit_module.Y_DELTA_PATTERN_70\
        );

    \I__535\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8354\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__8354\,
            I => \N__8351\
        );

    \I__533\ : Odrv12
    port map (
            O => \N__8351\,
            I => \TVP_VIDEO_c_3\
        );

    \I__532\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8345\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__8345\,
            I => \transmit_module.Y_DELTA_PATTERN_71\
        );

    \I__530\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__8339\,
            I => \transmit_module.Y_DELTA_PATTERN_35\
        );

    \INVTVP_VSYNC_buff_I_0.WIRE_OUT_0__9C\ : INV
    port map (
            O => \INVTVP_VSYNC_buff_I_0.WIRE_OUT_0__9C_net\,
            I => \N__24595\
        );

    \INVTVP_VSYNC_buff_I_0.BUFFER_0__i2C\ : INV
    port map (
            O => \INVTVP_VSYNC_buff_I_0.BUFFER_0__i2C_net\,
            I => \N__24586\
        );

    \INVTVP_VSYNC_buff_I_0.BUFFER_0__i1C\ : INV
    port map (
            O => \INVTVP_VSYNC_buff_I_0.BUFFER_0__i1C_net\,
            I => \N__24582\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3143\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3132\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.n3111\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3124\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3154\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.n3098\,
            carryinitout => \bfn_12_12_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \GB_BUFFER_DEBUG_c_2_c_THRU_LUT4_0_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24641\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_DEBUG_c_2_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i70_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8348\,
            lcout => \transmit_module.Y_DELTA_PATTERN_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23482\,
            ce => \N__15257\,
            sr => \N__20409\
        );

    \transmit_module.Y_DELTA_PATTERN_i69_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8363\,
            lcout => \transmit_module.Y_DELTA_PATTERN_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23500\,
            ce => \N__15251\,
            sr => \N__20285\
        );

    \tvp_video_buffer.BUFFER_0__i2_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8357\,
            lcout => \tvp_video_buffer.BUFFER_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i71_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8435\,
            lcout => \transmit_module.Y_DELTA_PATTERN_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23457\,
            ce => \N__15255\,
            sr => \N__20354\
        );

    \transmit_module.Y_DELTA_PATTERN_i35_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8408\,
            lcout => \transmit_module.Y_DELTA_PATTERN_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23317\,
            ce => \N__15250\,
            sr => \N__20298\
        );

    \transmit_module.Y_DELTA_PATTERN_i34_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8342\,
            lcout => \transmit_module.Y_DELTA_PATTERN_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23317\,
            ce => \N__15250\,
            sr => \N__20298\
        );

    \transmit_module.Y_DELTA_PATTERN_i33_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8441\,
            lcout => \transmit_module.Y_DELTA_PATTERN_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23319\,
            ce => \N__15248\,
            sr => \N__20414\
        );

    \transmit_module.Y_DELTA_PATTERN_i72_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8702\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23316\,
            ce => \N__15221\,
            sr => \N__20385\
        );

    \transmit_module.Y_DELTA_PATTERN_i87_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8414\,
            lcout => \transmit_module.Y_DELTA_PATTERN_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23506\,
            ce => \N__18406\,
            sr => \N__20416\
        );

    \transmit_module.Y_DELTA_PATTERN_i89_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8426\,
            lcout => \transmit_module.Y_DELTA_PATTERN_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23498\,
            ce => \N__18392\,
            sr => \N__20327\
        );

    \transmit_module.Y_DELTA_PATTERN_i90_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8675\,
            lcout => \transmit_module.Y_DELTA_PATTERN_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23498\,
            ce => \N__18392\,
            sr => \N__20327\
        );

    \transmit_module.Y_DELTA_PATTERN_i88_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8420\,
            lcout => \transmit_module.Y_DELTA_PATTERN_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23498\,
            ce => \N__18392\,
            sr => \N__20327\
        );

    \transmit_module.Y_DELTA_PATTERN_i96_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8651\,
            lcout => \transmit_module.Y_DELTA_PATTERN_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23422\,
            ce => \N__21047\,
            sr => \N__20413\
        );

    \transmit_module.Y_DELTA_PATTERN_i36_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8489\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23505\,
            ce => \N__15256\,
            sr => \N__20338\
        );

    \transmit_module.Y_DELTA_PATTERN_i79_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8495\,
            lcout => \transmit_module.Y_DELTA_PATTERN_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23505\,
            ce => \N__15256\,
            sr => \N__20338\
        );

    \transmit_module.Y_DELTA_PATTERN_i81_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8555\,
            lcout => \transmit_module.Y_DELTA_PATTERN_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23505\,
            ce => \N__15256\,
            sr => \N__20338\
        );

    \transmit_module.Y_DELTA_PATTERN_i80_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8501\,
            lcout => \transmit_module.Y_DELTA_PATTERN_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23505\,
            ce => \N__15256\,
            sr => \N__20338\
        );

    \transmit_module.Y_DELTA_PATTERN_i37_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9011\,
            lcout => \transmit_module.Y_DELTA_PATTERN_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23435\,
            ce => \N__15244\,
            sr => \N__20393\
        );

    \transmit_module.Y_DELTA_PATTERN_i78_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8483\,
            lcout => \transmit_module.Y_DELTA_PATTERN_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23435\,
            ce => \N__15244\,
            sr => \N__20393\
        );

    \transmit_module.Y_DELTA_PATTERN_i66_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8453\,
            lcout => \transmit_module.Y_DELTA_PATTERN_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23372\,
            ce => \N__15220\,
            sr => \N__20384\
        );

    \transmit_module.Y_DELTA_PATTERN_i48_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8543\,
            lcout => \transmit_module.Y_DELTA_PATTERN_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23372\,
            ce => \N__15220\,
            sr => \N__20384\
        );

    \transmit_module.Y_DELTA_PATTERN_i65_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8477\,
            lcout => \transmit_module.Y_DELTA_PATTERN_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23372\,
            ce => \N__15220\,
            sr => \N__20384\
        );

    \transmit_module.Y_DELTA_PATTERN_i68_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8471\,
            lcout => \transmit_module.Y_DELTA_PATTERN_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23372\,
            ce => \N__15220\,
            sr => \N__20384\
        );

    \transmit_module.Y_DELTA_PATTERN_i67_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8459\,
            lcout => \transmit_module.Y_DELTA_PATTERN_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23372\,
            ce => \N__15220\,
            sr => \N__20384\
        );

    \transmit_module.Y_DELTA_PATTERN_i47_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8447\,
            lcout => \transmit_module.Y_DELTA_PATTERN_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23372\,
            ce => \N__15220\,
            sr => \N__20384\
        );

    \tvp_video_buffer.BUFFER_0__i1_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8627\,
            lcout => \tvp_video_buffer.BUFFER_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14812\,
            in1 => \N__14668\,
            in2 => \N__14575\,
            in3 => \N__14474\,
            lcout => \line_buffer.n533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i10_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8567\,
            lcout => \tvp_video_buffer.BUFFER_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8525\,
            lcout => \transmit_module.Y_DELTA_PATTERN_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23516\,
            ce => \N__15254\,
            sr => \N__20336\
        );

    \transmit_module.Y_DELTA_PATTERN_i49_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8918\,
            lcout => \transmit_module.Y_DELTA_PATTERN_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23516\,
            ce => \N__15254\,
            sr => \N__20336\
        );

    \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8519\,
            lcout => \transmit_module.Y_DELTA_PATTERN_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23455\,
            ce => \N__18407\,
            sr => \N__20295\
        );

    \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8531\,
            lcout => \transmit_module.Y_DELTA_PATTERN_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23455\,
            ce => \N__18407\,
            sr => \N__20295\
        );

    \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8507\,
            lcout => \transmit_module.Y_DELTA_PATTERN_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23455\,
            ce => \N__18407\,
            sr => \N__20295\
        );

    \transmit_module.Y_DELTA_PATTERN_i86_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8513\,
            lcout => \transmit_module.Y_DELTA_PATTERN_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23455\,
            ce => \N__18407\,
            sr => \N__20295\
        );

    \transmit_module.Y_DELTA_PATTERN_i93_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8657\,
            lcout => \transmit_module.Y_DELTA_PATTERN_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23458\,
            ce => \N__18402\,
            sr => \N__20284\
        );

    \transmit_module.Y_DELTA_PATTERN_i91_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8663\,
            lcout => \transmit_module.Y_DELTA_PATTERN_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23458\,
            ce => \N__18402\,
            sr => \N__20284\
        );

    \transmit_module.Y_DELTA_PATTERN_i92_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8669\,
            lcout => \transmit_module.Y_DELTA_PATTERN_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23458\,
            ce => \N__18402\,
            sr => \N__20284\
        );

    \transmit_module.Y_DELTA_PATTERN_i94_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8633\,
            lcout => \transmit_module.Y_DELTA_PATTERN_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23303\,
            ce => \N__18391\,
            sr => \N__20293\
        );

    \transmit_module.Y_DELTA_PATTERN_i97_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8645\,
            lcout => \transmit_module.Y_DELTA_PATTERN_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23303\,
            ce => \N__18391\,
            sr => \N__20293\
        );

    \transmit_module.Y_DELTA_PATTERN_i98_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9041\,
            lcout => \transmit_module.Y_DELTA_PATTERN_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23303\,
            ce => \N__18391\,
            sr => \N__20293\
        );

    \transmit_module.Y_DELTA_PATTERN_i95_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8639\,
            lcout => \transmit_module.Y_DELTA_PATTERN_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23303\,
            ce => \N__18391\,
            sr => \N__20293\
        );

    \transmit_module.Y_DELTA_PATTERN_i28_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8732\,
            lcout => \transmit_module.Y_DELTA_PATTERN_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23468\,
            ce => \N__21032\,
            sr => \N__20337\
        );

    \transmit_module.Y_DELTA_PATTERN_i7_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8924\,
            lcout => \transmit_module.Y_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23468\,
            ce => \N__21032\,
            sr => \N__20337\
        );

    \transmit_module.Y_DELTA_PATTERN_i32_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8741\,
            lcout => \transmit_module.Y_DELTA_PATTERN_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23436\,
            ce => \N__21022\,
            sr => \N__20397\
        );

    \transmit_module.Y_DELTA_PATTERN_i29_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8714\,
            lcout => \transmit_module.Y_DELTA_PATTERN_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23436\,
            ce => \N__21022\,
            sr => \N__20397\
        );

    \transmit_module.Y_DELTA_PATTERN_i31_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8726\,
            lcout => \transmit_module.Y_DELTA_PATTERN_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23436\,
            ce => \N__21022\,
            sr => \N__20397\
        );

    \transmit_module.Y_DELTA_PATTERN_i30_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8720\,
            lcout => \transmit_module.Y_DELTA_PATTERN_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23436\,
            ce => \N__21022\,
            sr => \N__20397\
        );

    \transmit_module.Y_DELTA_PATTERN_i74_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23376\,
            ce => \N__15164\,
            sr => \N__20267\
        );

    \transmit_module.Y_DELTA_PATTERN_i73_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8708\,
            lcout => \transmit_module.Y_DELTA_PATTERN_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23376\,
            ce => \N__15164\,
            sr => \N__20267\
        );

    \transmit_module.Y_DELTA_PATTERN_i64_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8693\,
            lcout => \transmit_module.Y_DELTA_PATTERN_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23376\,
            ce => \N__15164\,
            sr => \N__20267\
        );

    \transmit_module.Y_DELTA_PATTERN_i62_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8681\,
            lcout => \transmit_module.Y_DELTA_PATTERN_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23161\,
            ce => \N__15240\,
            sr => \N__20297\
        );

    \transmit_module.Y_DELTA_PATTERN_i63_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8687\,
            lcout => \transmit_module.Y_DELTA_PATTERN_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23161\,
            ce => \N__15240\,
            sr => \N__20297\
        );

    \transmit_module.Y_DELTA_PATTERN_i75_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9266\,
            lcout => \transmit_module.Y_DELTA_PATTERN_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23161\,
            ce => \N__15240\,
            sr => \N__20297\
        );

    \transmit_module.Y_DELTA_PATTERN_i61_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8837\,
            lcout => \transmit_module.Y_DELTA_PATTERN_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23161\,
            ce => \N__15240\,
            sr => \N__20297\
        );

    \transmit_module.Y_DELTA_PATTERN_i77_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23161\,
            ce => \N__15240\,
            sr => \N__20297\
        );

    \tvp_video_buffer.BUFFER_0__i9_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8822\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.PULSE_1HZ_49_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8809\,
            in2 => \_gnd_net_\,
            in3 => \N__12530\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24590\,
            ce => \N__12622\,
            sr => \_gnd_net_\
        );

    \tvp_hs_buffer.BUFFER_0__i2_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8762\,
            lcout => \tvp_hs_buffer.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_hs_buffer.BUFFER_0__i1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8788\,
            lcout => \tvp_hs_buffer.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_hs_buffer.WIRE_OUT_0__9_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8756\,
            lcout => \TVP_HSYNC_buff\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.X_243__i0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8750\,
            in2 => \_gnd_net_\,
            in3 => \N__8744\,
            lcout => \receive_module.rx_counter.n10\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \receive_module.rx_counter.n3147\,
            clk => \N__24599\,
            ce => 'H',
            sr => \N__9415\
        );

    \receive_module.rx_counter.X_243__i1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8882\,
            in2 => \_gnd_net_\,
            in3 => \N__8876\,
            lcout => \receive_module.rx_counter.n9_adj_612\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3147\,
            carryout => \receive_module.rx_counter.n3148\,
            clk => \N__24599\,
            ce => 'H',
            sr => \N__9415\
        );

    \receive_module.rx_counter.X_243__i2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8873\,
            in2 => \_gnd_net_\,
            in3 => \N__8867\,
            lcout => \receive_module.rx_counter.n8_adj_611\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3148\,
            carryout => \receive_module.rx_counter.n3149\,
            clk => \N__24599\,
            ce => 'H',
            sr => \N__9415\
        );

    \receive_module.rx_counter.X_243__i3_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9572\,
            in2 => \_gnd_net_\,
            in3 => \N__8864\,
            lcout => \receive_module.rx_counter.X_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3149\,
            carryout => \receive_module.rx_counter.n3150\,
            clk => \N__24599\,
            ce => 'H',
            sr => \N__9415\
        );

    \receive_module.rx_counter.X_243__i4_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9587\,
            in2 => \_gnd_net_\,
            in3 => \N__8861\,
            lcout => \receive_module.rx_counter.X_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3150\,
            carryout => \receive_module.rx_counter.n3151\,
            clk => \N__24599\,
            ce => 'H',
            sr => \N__9415\
        );

    \receive_module.rx_counter.X_243__i5_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9602\,
            in2 => \_gnd_net_\,
            in3 => \N__8858\,
            lcout => \receive_module.rx_counter.X_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3151\,
            carryout => \receive_module.rx_counter.n3152\,
            clk => \N__24599\,
            ce => 'H',
            sr => \N__9415\
        );

    \receive_module.rx_counter.X_243__i6_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9557\,
            in2 => \_gnd_net_\,
            in3 => \N__8855\,
            lcout => \receive_module.rx_counter.X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3152\,
            carryout => \receive_module.rx_counter.n3153\,
            clk => \N__24599\,
            ce => 'H',
            sr => \N__9415\
        );

    \receive_module.rx_counter.X_243__i7_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9539\,
            in2 => \_gnd_net_\,
            in3 => \N__8852\,
            lcout => \receive_module.rx_counter.X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3153\,
            carryout => \receive_module.rx_counter.n3154\,
            clk => \N__24599\,
            ce => 'H',
            sr => \N__9415\
        );

    \receive_module.rx_counter.X_243__i8_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9443\,
            in2 => \_gnd_net_\,
            in3 => \N__8849\,
            lcout => \receive_module.rx_counter.X_8\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \receive_module.rx_counter.n3155\,
            clk => \N__24602\,
            ce => 'H',
            sr => \N__9416\
        );

    \receive_module.rx_counter.X_243__i9_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9430\,
            in2 => \_gnd_net_\,
            in3 => \N__8846\,
            lcout => \receive_module.rx_counter.X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24602\,
            ce => 'H',
            sr => \N__9416\
        );

    \receive_module.i246_2_lut_rep_26_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14675\,
            in2 => \_gnd_net_\,
            in3 => \N__13089\,
            lcout => \receive_module.n3632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8906\,
            lcout => \transmit_module.Y_DELTA_PATTERN_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23459\,
            ce => \N__15253\,
            sr => \N__20335\
        );

    \transmit_module.Y_DELTA_PATTERN_i50_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8912\,
            lcout => \transmit_module.Y_DELTA_PATTERN_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23459\,
            ce => \N__15253\,
            sr => \N__20335\
        );

    \transmit_module.Y_DELTA_PATTERN_i51_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9716\,
            lcout => \transmit_module.Y_DELTA_PATTERN_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23459\,
            ce => \N__15253\,
            sr => \N__20335\
        );

    \transmit_module.Y_DELTA_PATTERN_i58_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9320\,
            lcout => \transmit_module.Y_DELTA_PATTERN_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23459\,
            ce => \N__15253\,
            sr => \N__20335\
        );

    \transmit_module.Y_DELTA_PATTERN_i56_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8900\,
            lcout => \transmit_module.Y_DELTA_PATTERN_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23305\,
            ce => \N__15252\,
            sr => \N__20294\
        );

    \transmit_module.Y_DELTA_PATTERN_i22_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8972\,
            lcout => \transmit_module.Y_DELTA_PATTERN_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23472\,
            ce => \N__21033\,
            sr => \N__20251\
        );

    \transmit_module.Y_DELTA_PATTERN_i21_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8894\,
            lcout => \transmit_module.Y_DELTA_PATTERN_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23472\,
            ce => \N__21033\,
            sr => \N__20251\
        );

    \transmit_module.Y_DELTA_PATTERN_i20_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8888\,
            lcout => \transmit_module.Y_DELTA_PATTERN_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23472\,
            ce => \N__21033\,
            sr => \N__20251\
        );

    \transmit_module.Y_DELTA_PATTERN_i24_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8930\,
            lcout => \transmit_module.Y_DELTA_PATTERN_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23472\,
            ce => \N__21033\,
            sr => \N__20251\
        );

    \transmit_module.Y_DELTA_PATTERN_i23_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8978\,
            lcout => \transmit_module.Y_DELTA_PATTERN_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23472\,
            ce => \N__21033\,
            sr => \N__20251\
        );

    \transmit_module.Y_DELTA_PATTERN_i27_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8966\,
            lcout => \transmit_module.Y_DELTA_PATTERN_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23484\,
            ce => \N__21046\,
            sr => \N__20292\
        );

    \transmit_module.Y_DELTA_PATTERN_i26_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8960\,
            lcout => \transmit_module.Y_DELTA_PATTERN_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23484\,
            ce => \N__21046\,
            sr => \N__20292\
        );

    \transmit_module.Y_DELTA_PATTERN_i15_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18311\,
            lcout => \transmit_module.Y_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23484\,
            ce => \N__21046\,
            sr => \N__20292\
        );

    \transmit_module.Y_DELTA_PATTERN_i12_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8954\,
            lcout => \transmit_module.Y_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23484\,
            ce => \N__21046\,
            sr => \N__20292\
        );

    \transmit_module.Y_DELTA_PATTERN_i13_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8942\,
            lcout => \transmit_module.Y_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23484\,
            ce => \N__21046\,
            sr => \N__20292\
        );

    \transmit_module.Y_DELTA_PATTERN_i14_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8948\,
            lcout => \transmit_module.Y_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23484\,
            ce => \N__21046\,
            sr => \N__20292\
        );

    \transmit_module.Y_DELTA_PATTERN_i25_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8936\,
            lcout => \transmit_module.Y_DELTA_PATTERN_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23484\,
            ce => \N__21046\,
            sr => \N__20292\
        );

    \transmit_module.Y_DELTA_PATTERN_i8_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9029\,
            lcout => \transmit_module.Y_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23377\,
            ce => \N__21009\,
            sr => \N__20164\
        );

    \transmit_module.Y_DELTA_PATTERN_i99_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20657\,
            lcout => \transmit_module.Y_DELTA_PATTERN_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23377\,
            ce => \N__21009\,
            sr => \N__20164\
        );

    \transmit_module.Y_DELTA_PATTERN_i10_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9017\,
            lcout => \transmit_module.Y_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23377\,
            ce => \N__21009\,
            sr => \N__20164\
        );

    \transmit_module.Y_DELTA_PATTERN_i9_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9035\,
            lcout => \transmit_module.Y_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23377\,
            ce => \N__21009\,
            sr => \N__20164\
        );

    \transmit_module.Y_DELTA_PATTERN_i11_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9023\,
            lcout => \transmit_module.Y_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23377\,
            ce => \N__21009\,
            sr => \N__20164\
        );

    \transmit_module.Y_DELTA_PATTERN_i40_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8990\,
            lcout => \transmit_module.Y_DELTA_PATTERN_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23434\,
            ce => \N__15212\,
            sr => \N__20392\
        );

    \transmit_module.Y_DELTA_PATTERN_i38_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8996\,
            lcout => \transmit_module.Y_DELTA_PATTERN_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23434\,
            ce => \N__15212\,
            sr => \N__20392\
        );

    \transmit_module.Y_DELTA_PATTERN_i39_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9002\,
            lcout => \transmit_module.Y_DELTA_PATTERN_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23434\,
            ce => \N__15212\,
            sr => \N__20392\
        );

    \transmit_module.Y_DELTA_PATTERN_i41_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8984\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23434\,
            ce => \N__15212\,
            sr => \N__20392\
        );

    \transmit_module.Y_DELTA_PATTERN_i42_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9326\,
            lcout => \transmit_module.Y_DELTA_PATTERN_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23371\,
            ce => \N__15199\,
            sr => \N__20339\
        );

    \transmit_module.Y_DELTA_PATTERN_i45_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9290\,
            lcout => \transmit_module.Y_DELTA_PATTERN_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23371\,
            ce => \N__15199\,
            sr => \N__20339\
        );

    \transmit_module.Y_DELTA_PATTERN_i43_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9305\,
            lcout => \transmit_module.Y_DELTA_PATTERN_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23371\,
            ce => \N__15199\,
            sr => \N__20339\
        );

    \transmit_module.Y_DELTA_PATTERN_i59_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9278\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23371\,
            ce => \N__15199\,
            sr => \N__20339\
        );

    \transmit_module.Y_DELTA_PATTERN_i44_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9311\,
            lcout => \transmit_module.Y_DELTA_PATTERN_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23371\,
            ce => \N__15199\,
            sr => \N__20339\
        );

    \transmit_module.Y_DELTA_PATTERN_i46_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9299\,
            lcout => \transmit_module.Y_DELTA_PATTERN_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23371\,
            ce => \N__15199\,
            sr => \N__20339\
        );

    \transmit_module.Y_DELTA_PATTERN_i60_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9284\,
            lcout => \transmit_module.Y_DELTA_PATTERN_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23154\,
            ce => \N__15219\,
            sr => \N__20296\
        );

    \transmit_module.Y_DELTA_PATTERN_i76_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9272\,
            lcout => \transmit_module.Y_DELTA_PATTERN_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23154\,
            ce => \N__15219\,
            sr => \N__20296\
        );

    \transmit_module.i1613_4_lut_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20877\,
            in1 => \N__20557\,
            in2 => \N__20408\,
            in3 => \N__18245\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i3_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9053\,
            lcout => \tvp_video_buffer.BUFFER_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TVP_VSYNC_buff_I_0.BUFFER_0__i1_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9469\,
            lcout => \TVP_VSYNC_buff_I_0.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVTVP_VSYNC_buff_I_0.BUFFER_0__i1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i130_2_lut_rep_17_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12521\,
            lcout => \receive_module.rx_counter.n3623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TVP_VSYNC_buff_I_0.BUFFER_0__i2_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9449\,
            lcout => \TVP_VSYNC_buff_I_0.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVTVP_VSYNC_buff_I_0.BUFFER_0__i2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_HS_51_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9508\,
            lcout => \receive_module.rx_counter.old_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i59_4_lut_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011100101"
        )
    port map (
            in0 => \N__9442\,
            in1 => \N__9653\,
            in2 => \N__9431\,
            in3 => \N__9524\,
            lcout => \receive_module.rx_counter.n55_adj_606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_1_lut_rep_24_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.rx_counter.n3630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TVP_VSYNC_buff_I_0.WIRE_OUT_0__9_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9392\,
            lcout => \TVP_VSYNC_buff\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVTVP_VSYNC_buff_I_0.WIRE_OUT_0__9C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__14794\,
            in1 => \N__14643\,
            in2 => \N__14560\,
            in3 => \N__14455\,
            lcout => \line_buffer.n467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_18_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9570\,
            in2 => \_gnd_net_\,
            in3 => \N__9585\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_adj_19_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__9601\,
            in1 => \N__9555\,
            in2 => \N__9656\,
            in3 => \N__9537\,
            lcout => \receive_module.rx_counter.n3400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14649\,
            in1 => \N__14795\,
            in2 => \N__14561\,
            in3 => \N__14467\,
            lcout => \line_buffer.n565\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_adj_20_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9600\,
            in2 => \_gnd_net_\,
            in3 => \N__9586\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2042_4_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__9571\,
            in1 => \N__9556\,
            in2 => \N__9542\,
            in3 => \N__9538\,
            lcout => \receive_module.rx_counter.n3385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.O_VS_I_0_1_lut_rep_25_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13067\,
            lcout => \receive_module.n3631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i249_3_lut_3_lut_3_lut_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__13068\,
            in1 => \N__9518\,
            in2 => \_gnd_net_\,
            in3 => \N__9509\,
            lcout => \receive_module.rx_counter.n2063\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_2_lut_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10128\,
            in2 => \_gnd_net_\,
            in3 => \N__9488\,
            lcout => \receive_module.n136\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \receive_module.n3091\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_3_lut_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9870\,
            in2 => \_gnd_net_\,
            in3 => \N__9485\,
            lcout => \receive_module.n135\,
            ltout => OPEN,
            carryin => \receive_module.n3091\,
            carryout => \receive_module.n3092\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_4_lut_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12831\,
            in2 => \_gnd_net_\,
            in3 => \N__9482\,
            lcout => \receive_module.n134\,
            ltout => OPEN,
            carryin => \receive_module.n3092\,
            carryout => \receive_module.n3093\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_5_lut_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12045\,
            in2 => \_gnd_net_\,
            in3 => \N__9683\,
            lcout => \receive_module.n133\,
            ltout => OPEN,
            carryin => \receive_module.n3093\,
            carryout => \receive_module.n3094\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_6_lut_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11787\,
            in2 => \_gnd_net_\,
            in3 => \N__9680\,
            lcout => \receive_module.n132\,
            ltout => OPEN,
            carryin => \receive_module.n3094\,
            carryout => \receive_module.n3095\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_7_lut_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11403\,
            in2 => \_gnd_net_\,
            in3 => \N__9677\,
            lcout => \receive_module.n131\,
            ltout => OPEN,
            carryin => \receive_module.n3095\,
            carryout => \receive_module.n3096\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_8_lut_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11145\,
            in2 => \_gnd_net_\,
            in3 => \N__9674\,
            lcout => \receive_module.n130\,
            ltout => OPEN,
            carryin => \receive_module.n3096\,
            carryout => \receive_module.n3097\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_9_lut_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10872\,
            in2 => \_gnd_net_\,
            in3 => \N__9671\,
            lcout => \receive_module.n129\,
            ltout => OPEN,
            carryin => \receive_module.n3097\,
            carryout => \receive_module.n3098\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_10_lut_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10632\,
            in2 => \_gnd_net_\,
            in3 => \N__9668\,
            lcout => \receive_module.n128\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \receive_module.n3099\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_11_lut_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10371\,
            in2 => \_gnd_net_\,
            in3 => \N__9665\,
            lcout => \receive_module.n127\,
            ltout => OPEN,
            carryin => \receive_module.n3099\,
            carryout => \receive_module.n3100\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_12_lut_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12294\,
            in2 => \_gnd_net_\,
            in3 => \N__9662\,
            lcout => \receive_module.n126\,
            ltout => OPEN,
            carryin => \receive_module.n3100\,
            carryout => \receive_module.n3101\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i11_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14430\,
            in2 => \_gnd_net_\,
            in3 => \N__9659\,
            lcout => \RX_ADDR_11\,
            ltout => OPEN,
            carryin => \receive_module.n3101\,
            carryout => \receive_module.n3102\,
            clk => \N__24605\,
            ce => \N__9734\,
            sr => \N__12761\
        );

    \receive_module.BRAM_ADDR__i12_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14778\,
            in2 => \_gnd_net_\,
            in3 => \N__9740\,
            lcout => \RX_ADDR_12\,
            ltout => OPEN,
            carryin => \receive_module.n3102\,
            carryout => \receive_module.n3103\,
            clk => \N__24605\,
            ce => \N__9734\,
            sr => \N__12761\
        );

    \receive_module.BRAM_ADDR__i13_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14532\,
            in2 => \_gnd_net_\,
            in3 => \N__9737\,
            lcout => \RX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24605\,
            ce => \N__9734\,
            sr => \N__12761\
        );

    \transmit_module.Y_DELTA_PATTERN_i53_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9698\,
            lcout => \transmit_module.Y_DELTA_PATTERN_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23486\,
            ce => \N__15249\,
            sr => \N__20415\
        );

    \transmit_module.Y_DELTA_PATTERN_i52_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9722\,
            lcout => \transmit_module.Y_DELTA_PATTERN_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23486\,
            ce => \N__15249\,
            sr => \N__20415\
        );

    \transmit_module.Y_DELTA_PATTERN_i55_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9710\,
            lcout => \transmit_module.Y_DELTA_PATTERN_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23486\,
            ce => \N__15249\,
            sr => \N__20415\
        );

    \transmit_module.Y_DELTA_PATTERN_i54_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9704\,
            lcout => \transmit_module.Y_DELTA_PATTERN_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23486\,
            ce => \N__15249\,
            sr => \N__20415\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15299\,
            in2 => \_gnd_net_\,
            in3 => \N__13632\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3629_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__9689\,
            in1 => \N__13656\,
            in2 => \N__9692\,
            in3 => \N__13340\,
            lcout => \transmit_module.video_signal_controller.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1653_2_lut_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13291\,
            in2 => \_gnd_net_\,
            in3 => \N__13312\,
            lcout => \transmit_module.video_signal_controller.n2901\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_X_i0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13292\,
            in2 => \_gnd_net_\,
            in3 => \N__9767\,
            lcout => \transmit_module.video_signal_controller.VGA_X_0\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \transmit_module.video_signal_controller.n3125\,
            clk => \N__23132\,
            ce => 'H',
            sr => \N__14248\
        );

    \transmit_module.video_signal_controller.VGA_X_i1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13313\,
            in2 => \_gnd_net_\,
            in3 => \N__9764\,
            lcout => \transmit_module.video_signal_controller.VGA_X_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3125\,
            carryout => \transmit_module.video_signal_controller.n3126\,
            clk => \N__23132\,
            ce => 'H',
            sr => \N__14248\
        );

    \transmit_module.video_signal_controller.VGA_X_i2_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13341\,
            in2 => \_gnd_net_\,
            in3 => \N__9761\,
            lcout => \transmit_module.video_signal_controller.VGA_X_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3126\,
            carryout => \transmit_module.video_signal_controller.n3127\,
            clk => \N__23132\,
            ce => 'H',
            sr => \N__14248\
        );

    \transmit_module.video_signal_controller.VGA_X_i3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13657\,
            in2 => \_gnd_net_\,
            in3 => \N__9758\,
            lcout => \transmit_module.video_signal_controller.VGA_X_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3127\,
            carryout => \transmit_module.video_signal_controller.n3128\,
            clk => \N__23132\,
            ce => 'H',
            sr => \N__14248\
        );

    \transmit_module.video_signal_controller.VGA_X_i4_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13514\,
            in2 => \_gnd_net_\,
            in3 => \N__9755\,
            lcout => \transmit_module.video_signal_controller.VGA_X_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3128\,
            carryout => \transmit_module.video_signal_controller.n3129\,
            clk => \N__23132\,
            ce => 'H',
            sr => \N__14248\
        );

    \transmit_module.video_signal_controller.VGA_X_i5_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13634\,
            in2 => \_gnd_net_\,
            in3 => \N__9752\,
            lcout => \transmit_module.video_signal_controller.VGA_X_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3129\,
            carryout => \transmit_module.video_signal_controller.n3130\,
            clk => \N__23132\,
            ce => 'H',
            sr => \N__14248\
        );

    \transmit_module.video_signal_controller.VGA_X_i6_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15300\,
            in2 => \_gnd_net_\,
            in3 => \N__9749\,
            lcout => \transmit_module.video_signal_controller.VGA_X_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3130\,
            carryout => \transmit_module.video_signal_controller.n3131\,
            clk => \N__23132\,
            ce => 'H',
            sr => \N__14248\
        );

    \transmit_module.video_signal_controller.VGA_X_i7_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13539\,
            in2 => \_gnd_net_\,
            in3 => \N__9746\,
            lcout => \transmit_module.video_signal_controller.VGA_X_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3131\,
            carryout => \transmit_module.video_signal_controller.n3132\,
            clk => \N__23132\,
            ce => 'H',
            sr => \N__14248\
        );

    \transmit_module.video_signal_controller.VGA_X_i8_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15350\,
            in2 => \_gnd_net_\,
            in3 => \N__9743\,
            lcout => \transmit_module.video_signal_controller.VGA_X_8\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \transmit_module.video_signal_controller.n3133\,
            clk => \N__23404\,
            ce => 'H',
            sr => \N__14252\
        );

    \transmit_module.video_signal_controller.VGA_X_i9_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13602\,
            in2 => \_gnd_net_\,
            in3 => \N__9800\,
            lcout => \transmit_module.video_signal_controller.VGA_X_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3133\,
            carryout => \transmit_module.video_signal_controller.n3134\,
            clk => \N__23404\,
            ce => 'H',
            sr => \N__14252\
        );

    \transmit_module.video_signal_controller.VGA_X_i10_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13573\,
            in2 => \_gnd_net_\,
            in3 => \N__9797\,
            lcout => \transmit_module.video_signal_controller.VGA_X_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3134\,
            carryout => \transmit_module.video_signal_controller.n3135\,
            clk => \N__23404\,
            ce => 'H',
            sr => \N__14252\
        );

    \transmit_module.video_signal_controller.VGA_X_i11_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16716\,
            in2 => \_gnd_net_\,
            in3 => \N__9794\,
            lcout => \transmit_module.video_signal_controller.VGA_X_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23404\,
            ce => 'H',
            sr => \N__14252\
        );

    \transmit_module.i123_2_lut_4_lut_rep_29_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__16403\,
            in1 => \N__16427\,
            in2 => \N__20326\,
            in3 => \N__16369\,
            lcout => \transmit_module.n3635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9791\,
            lcout => \transmit_module.Y_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23229\,
            ce => \N__20990\,
            sr => \N__20260\
        );

    \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9785\,
            lcout => \transmit_module.Y_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23229\,
            ce => \N__20990\,
            sr => \N__20260\
        );

    \transmit_module.Y_DELTA_PATTERN_i3_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9773\,
            lcout => \transmit_module.Y_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23229\,
            ce => \N__20990\,
            sr => \N__20260\
        );

    \transmit_module.Y_DELTA_PATTERN_i5_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11615\,
            lcout => \transmit_module.Y_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23229\,
            ce => \N__20990\,
            sr => \N__20260\
        );

    \transmit_module.Y_DELTA_PATTERN_i4_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9779\,
            lcout => \transmit_module.Y_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23229\,
            ce => \N__20990\,
            sr => \N__20260\
        );

    \transmit_module.Y_DELTA_PATTERN_i6_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11627\,
            lcout => \transmit_module.Y_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23229\,
            ce => \N__20990\,
            sr => \N__20260\
        );

    \receive_module.BRAM_ADDR__i5_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__11609\,
            in1 => \N__11378\,
            in2 => \N__14732\,
            in3 => \N__13118\,
            lcout => \RX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24614\,
            ce => 'H',
            sr => \N__12786\
        );

    \receive_module.BRAM_ADDR__i6_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__13119\,
            in1 => \N__14718\,
            in2 => \N__11129\,
            in3 => \N__11351\,
            lcout => \RX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24614\,
            ce => 'H',
            sr => \N__12786\
        );

    \receive_module.BRAM_ADDR__i7_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__10862\,
            in1 => \N__11090\,
            in2 => \N__14733\,
            in3 => \N__13120\,
            lcout => \RX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24614\,
            ce => 'H',
            sr => \N__12786\
        );

    \receive_module.BRAM_ADDR__i8_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__13121\,
            in1 => \N__14722\,
            in2 => \N__10625\,
            in3 => \N__10835\,
            lcout => \RX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24614\,
            ce => 'H',
            sr => \N__12786\
        );

    \receive_module.BRAM_ADDR__i9_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__10356\,
            in1 => \N__10586\,
            in2 => \N__14734\,
            in3 => \N__13122\,
            lcout => \RX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24614\,
            ce => 'H',
            sr => \N__12786\
        );

    \receive_module.BRAM_ADDR__i0_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__10334\,
            in1 => \N__10106\,
            in2 => \N__14731\,
            in3 => \N__13116\,
            lcout => \RX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24614\,
            ce => 'H',
            sr => \N__12786\
        );

    \receive_module.BRAM_ADDR__i1_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__13117\,
            in1 => \N__14714\,
            in2 => \N__10079\,
            in3 => \N__9851\,
            lcout => \RX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24614\,
            ce => 'H',
            sr => \N__12786\
        );

    \line_buffer.i2158_3_lut_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24358\,
            in1 => \N__9824\,
            in2 => \_gnd_net_\,
            in3 => \N__9812\,
            lcout => \line_buffer.n3501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i10_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__12269\,
            in1 => \N__12494\,
            in2 => \N__14738\,
            in3 => \N__13129\,
            lcout => \RX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24619\,
            ce => 'H',
            sr => \N__12795\
        );

    \receive_module.BRAM_ADDR__i3_LC_12_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__12239\,
            in1 => \N__12017\,
            in2 => \N__14729\,
            in3 => \N__13141\,
            lcout => \RX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24626\,
            ce => 'H',
            sr => \N__12808\
        );

    \receive_module.BRAM_ADDR__i4_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__11990\,
            in1 => \N__11759\,
            in2 => \N__14730\,
            in3 => \N__13142\,
            lcout => \RX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24628\,
            ce => 'H',
            sr => \N__12809\
        );

    \tvp_video_buffer.WIRE_OUT_i0_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11732\,
            lcout => \RX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12563\,
            in2 => \_gnd_net_\,
            in3 => \N__11639\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_0\,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \receive_module.rx_counter.n3156\,
            clk => \N__24576\,
            ce => \N__12623\,
            sr => \N__12506\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12575\,
            in2 => \_gnd_net_\,
            in3 => \N__11636\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3156\,
            carryout => \receive_module.rx_counter.n3157\,
            clk => \N__24576\,
            ce => \N__12623\,
            sr => \N__12506\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12599\,
            in2 => \_gnd_net_\,
            in3 => \N__11633\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3157\,
            carryout => \receive_module.rx_counter.n3158\,
            clk => \N__24576\,
            ce => \N__12623\,
            sr => \N__12506\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12551\,
            in2 => \_gnd_net_\,
            in3 => \N__11630\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3158\,
            carryout => \receive_module.rx_counter.n3159\,
            clk => \N__24576\,
            ce => \N__12623\,
            sr => \N__12506\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12611\,
            in2 => \_gnd_net_\,
            in3 => \N__12629\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3159\,
            carryout => \receive_module.rx_counter.n3160\,
            clk => \N__24576\,
            ce => \N__12623\,
            sr => \N__12506\
        );

    \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12587\,
            in2 => \_gnd_net_\,
            in3 => \N__12626\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24576\,
            ce => \N__12623\,
            sr => \N__12506\
        );

    \receive_module.rx_counter.i1_4_lut_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__13868\,
            in1 => \N__13708\,
            in2 => \N__13898\,
            in3 => \N__12701\,
            lcout => \receive_module.rx_counter.n4_adj_605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_22_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12610\,
            in2 => \_gnd_net_\,
            in3 => \N__12598\,
            lcout => \receive_module.rx_counter.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_VS_52_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.rx_counter.old_VS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2130_2_lut_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12586\,
            in2 => \_gnd_net_\,
            in3 => \N__12574\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3473_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_4_lut_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__12562\,
            in1 => \N__12550\,
            in2 => \N__12539\,
            in3 => \N__12536\,
            lcout => \receive_module.rx_counter.n11\,
            ltout => \receive_module.rx_counter.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1281_2_lut_3_lut_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12520\,
            in2 => \N__12509\,
            in3 => \N__13086\,
            lcout => \receive_module.rx_counter.n2529\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__12641\,
            in1 => \N__12713\,
            in2 => \N__13769\,
            in3 => \N__12707\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3422_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.O_VISIBLE_53_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__12728\,
            in1 => \N__13768\,
            in2 => \N__12722\,
            in3 => \N__12719\,
            lcout => \RX_WE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13736\,
            in1 => \N__13838\,
            in2 => \_gnd_net_\,
            in3 => \N__13788\,
            lcout => \receive_module.rx_counter.n3394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_3_lut_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13210\,
            in1 => \N__13862\,
            in2 => \_gnd_net_\,
            in3 => \N__13192\,
            lcout => \receive_module.rx_counter.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__13735\,
            in1 => \N__13811\,
            in2 => \N__13841\,
            in3 => \N__13787\,
            lcout => \receive_module.rx_counter.n3413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__14620\,
            in1 => \N__14810\,
            in2 => \N__14573\,
            in3 => \N__14471\,
            lcout => \line_buffer.n596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i595_2_lut_rep_27_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13191\,
            in2 => \_gnd_net_\,
            in3 => \N__13209\,
            lcout => \receive_module.rx_counter.n3633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_21_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13889\,
            lcout => \receive_module.rx_counter.n4_adj_604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.Y__i0_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13733\,
            in2 => \_gnd_net_\,
            in3 => \N__12635\,
            lcout => \receive_module.rx_counter.Y_0\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \receive_module.rx_counter.n3117\,
            clk => \N__24592\,
            ce => \N__13166\,
            sr => \N__12771\
        );

    \receive_module.rx_counter.Y__i1_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13839\,
            in2 => \_gnd_net_\,
            in3 => \N__12632\,
            lcout => \receive_module.rx_counter.Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3117\,
            carryout => \receive_module.rx_counter.n3118\,
            clk => \N__24592\,
            ce => \N__13166\,
            sr => \N__12771\
        );

    \receive_module.rx_counter.Y__i2_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13789\,
            in2 => \_gnd_net_\,
            in3 => \N__13220\,
            lcout => \receive_module.rx_counter.Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3118\,
            carryout => \receive_module.rx_counter.n3119\,
            clk => \N__24592\,
            ce => \N__13166\,
            sr => \N__12771\
        );

    \receive_module.rx_counter.Y__i3_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13813\,
            in2 => \_gnd_net_\,
            in3 => \N__13217\,
            lcout => \receive_module.rx_counter.Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3119\,
            carryout => \receive_module.rx_counter.n3120\,
            clk => \N__24592\,
            ce => \N__13166\,
            sr => \N__12771\
        );

    \receive_module.rx_counter.Y__i4_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13890\,
            in2 => \_gnd_net_\,
            in3 => \N__13214\,
            lcout => \receive_module.rx_counter.Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3120\,
            carryout => \receive_module.rx_counter.n3121\,
            clk => \N__24592\,
            ce => \N__13166\,
            sr => \N__12771\
        );

    \receive_module.rx_counter.Y__i5_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13211\,
            in2 => \_gnd_net_\,
            in3 => \N__13196\,
            lcout => \receive_module.rx_counter.Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3121\,
            carryout => \receive_module.rx_counter.n3122\,
            clk => \N__24592\,
            ce => \N__13166\,
            sr => \N__12771\
        );

    \receive_module.rx_counter.Y__i6_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13193\,
            in2 => \_gnd_net_\,
            in3 => \N__13175\,
            lcout => \receive_module.rx_counter.Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3122\,
            carryout => \receive_module.rx_counter.n3123\,
            clk => \N__24592\,
            ce => \N__13166\,
            sr => \N__12771\
        );

    \receive_module.rx_counter.Y__i7_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13867\,
            in2 => \_gnd_net_\,
            in3 => \N__13172\,
            lcout => \receive_module.rx_counter.Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3123\,
            carryout => \receive_module.rx_counter.n3124\,
            clk => \N__24592\,
            ce => \N__13166\,
            sr => \N__12771\
        );

    \receive_module.rx_counter.Y__i8_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13763\,
            in2 => \_gnd_net_\,
            in3 => \N__13169\,
            lcout => \receive_module.rx_counter.Y_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24596\,
            ce => \N__13165\,
            sr => \N__12760\
        );

    \receive_module.BRAM_ADDR__i2_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__13148\,
            in1 => \N__12830\,
            in2 => \N__14669\,
            in3 => \N__13095\,
            lcout => \RX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24600\,
            ce => 'H',
            sr => \N__12772\
        );

    \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14873\,
            in2 => \_gnd_net_\,
            in3 => \N__12731\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_0\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \transmit_module.video_signal_controller.n3136\,
            clk => \N__23501\,
            ce => \N__14247\,
            sr => \N__14203\
        );

    \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14896\,
            in2 => \_gnd_net_\,
            in3 => \N__13247\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3136\,
            carryout => \transmit_module.video_signal_controller.n3137\,
            clk => \N__23501\,
            ce => \N__14247\,
            sr => \N__14203\
        );

    \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15381\,
            in2 => \_gnd_net_\,
            in3 => \N__13244\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3137\,
            carryout => \transmit_module.video_signal_controller.n3138\,
            clk => \N__23501\,
            ce => \N__14247\,
            sr => \N__14203\
        );

    \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14922\,
            in2 => \_gnd_net_\,
            in3 => \N__13241\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3138\,
            carryout => \transmit_module.video_signal_controller.n3139\,
            clk => \N__23501\,
            ce => \N__14247\,
            sr => \N__14203\
        );

    \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15528\,
            in2 => \_gnd_net_\,
            in3 => \N__13238\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3139\,
            carryout => \transmit_module.video_signal_controller.n3140\,
            clk => \N__23501\,
            ce => \N__14247\,
            sr => \N__14203\
        );

    \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14955\,
            in2 => \_gnd_net_\,
            in3 => \N__13235\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3140\,
            carryout => \transmit_module.video_signal_controller.n3141\,
            clk => \N__23501\,
            ce => \N__14247\,
            sr => \N__14203\
        );

    \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15012\,
            in2 => \_gnd_net_\,
            in3 => \N__13232\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3141\,
            carryout => \transmit_module.video_signal_controller.n3142\,
            clk => \N__23501\,
            ce => \N__14247\,
            sr => \N__14203\
        );

    \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15048\,
            in2 => \_gnd_net_\,
            in3 => \N__13229\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3142\,
            carryout => \transmit_module.video_signal_controller.n3143\,
            clk => \N__23501\,
            ce => \N__14247\,
            sr => \N__14203\
        );

    \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15073\,
            in2 => \_gnd_net_\,
            in3 => \N__13226\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_8\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \transmit_module.video_signal_controller.n3144\,
            clk => \N__23364\,
            ce => \N__14246\,
            sr => \N__14207\
        );

    \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15488\,
            in2 => \_gnd_net_\,
            in3 => \N__13223\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3144\,
            carryout => \transmit_module.video_signal_controller.n3145\,
            clk => \N__23364\,
            ce => \N__14246\,
            sr => \N__14207\
        );

    \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15429\,
            in2 => \_gnd_net_\,
            in3 => \N__13406\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3145\,
            carryout => \transmit_module.video_signal_controller.n3146\,
            clk => \N__23364\,
            ce => \N__14246\,
            sr => \N__14207\
        );

    \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14983\,
            in2 => \_gnd_net_\,
            in3 => \N__13403\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23364\,
            ce => \N__14246\,
            sr => \N__14207\
        );

    \transmit_module.video_signal_controller.i485_4_lut_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__13349\,
            in1 => \N__13256\,
            in2 => \N__13274\,
            in3 => \N__15352\,
            lcout => \transmit_module.video_signal_controller.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__14653\,
            in1 => \N__14803\,
            in2 => \N__14565\,
            in3 => \N__14456\,
            lcout => \line_buffer.n564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_adj_26_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13511\,
            in2 => \_gnd_net_\,
            in3 => \N__13655\,
            lcout => \transmit_module.video_signal_controller.n3313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__15304\,
            in1 => \N__13631\,
            in2 => \_gnd_net_\,
            in3 => \N__13538\,
            lcout => \transmit_module.video_signal_controller.n2001\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1585_2_lut_rep_18_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__13310\,
            in1 => \_gnd_net_\,
            in2 => \N__13342\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.video_signal_controller.n3624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1669_2_lut_3_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13343\,
            in1 => \N__13311\,
            in2 => \_gnd_net_\,
            in3 => \N__13290\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2917_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1699_4_lut_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__13270\,
            in1 => \N__15351\,
            in2 => \N__13259\,
            in3 => \N__13255\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2947_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1705_4_lut_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__16717\,
            in1 => \N__13604\,
            in2 => \N__13697\,
            in3 => \N__13577\,
            lcout => \transmit_module.video_signal_controller.n2036\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3591_bdd_4_lut_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__23806\,
            in1 => \N__13412\,
            in2 => \N__13694\,
            in3 => \N__13676\,
            lcout => \line_buffer.n3594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__13541\,
            in1 => \N__13512\,
            in2 => \N__13661\,
            in3 => \N__13633\,
            lcout => \transmit_module.video_signal_controller.n4_adj_617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101010110"
        )
    port map (
            in0 => \N__13572\,
            in1 => \N__13610\,
            in2 => \N__13603\,
            in3 => \N__16711\,
            lcout => \transmit_module.video_signal_controller.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_rep_19_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13595\,
            in1 => \N__13568\,
            in2 => \_gnd_net_\,
            in3 => \N__16712\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2128_4_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__13547\,
            in1 => \N__13540\,
            in2 => \N__13517\,
            in3 => \N__13513\,
            lcout => \transmit_module.video_signal_controller.n3471\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14654\,
            in1 => \N__14799\,
            in2 => \N__14566\,
            in3 => \N__14460\,
            lcout => \line_buffer.n597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2245_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24339\,
            in1 => \N__13445\,
            in2 => \N__23841\,
            in3 => \N__13427\,
            lcout => \line_buffer.n3591\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14900\,
            in2 => \_gnd_net_\,
            in3 => \N__15385\,
            lcout => \transmit_module.video_signal_controller.n3628\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__14811\,
            in1 => \N__14655\,
            in2 => \N__14574\,
            in3 => \N__14472\,
            lcout => \line_buffer.n468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i4_3_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20635\,
            in1 => \N__13916\,
            in2 => \_gnd_net_\,
            in3 => \N__16501\,
            lcout => \transmit_module.n113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1612_4_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20763\,
            in1 => \N__20016\,
            in2 => \N__14857\,
            in3 => \N__15268\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16505\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22976\,
            ce => \N__20454\,
            sr => \N__20240\
        );

    \tvp_video_buffer.BUFFER_0__i11_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13910\,
            lcout => \tvp_video_buffer.BUFFER_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24565\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13891\,
            in2 => \_gnd_net_\,
            in3 => \N__13863\,
            lcout => \receive_module.rx_counter.n10_adj_610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i6_4_lut_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__13840\,
            in1 => \N__13814\,
            in2 => \N__13793\,
            in3 => \N__13764\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.SYNC_46_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13742\,
            in1 => \N__13734\,
            in2 => \N__13712\,
            in3 => \N__13709\,
            lcout => \RX_TX_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.BUFFER_0__i2_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14819\,
            lcout => \sync_buffer.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.BUFFER_0__i1_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14825\,
            lcout => \sync_buffer.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__14813\,
            in1 => \N__14621\,
            in2 => \N__14576\,
            in3 => \N__14473\,
            lcout => \line_buffer.n532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i1_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14360\,
            lcout => \RX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.WIRE_OUT_0__9_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14267\,
            lcout => \RX_TX_SYNC_BUFF\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1138_2_lut_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14258\,
            in2 => \_gnd_net_\,
            in3 => \N__14239\,
            lcout => \transmit_module.video_signal_controller.n2378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_28_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14916\,
            in1 => \N__14891\,
            in2 => \_gnd_net_\,
            in3 => \N__15377\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__15527\,
            in1 => \N__14954\,
            in2 => \N__14186\,
            in3 => \N__15005\,
            lcout => \transmit_module.video_signal_controller.n3412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i0_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20855\,
            in1 => \N__16097\,
            in2 => \N__20288\,
            in3 => \N__16081\,
            lcout => \transmit_module.TX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14872\,
            lcout => \transmit_module.video_signal_controller.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i1_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__15851\,
            in1 => \N__15826\,
            in2 => \N__20875\,
            in3 => \N__20259\,
            lcout => \transmit_module.TX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i2_3_lut_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21612\,
            in1 => \_gnd_net_\,
            in2 => \N__16520\,
            in3 => \N__18282\,
            lcout => \transmit_module.n146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2124_2_lut_rep_16_3_lut_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__15052\,
            in1 => \_gnd_net_\,
            in2 => \N__15017\,
            in3 => \N__15072\,
            lcout => \transmit_module.video_signal_controller.n3622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i3_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20869\,
            in1 => \N__14861\,
            in2 => \N__20258\,
            in3 => \N__15275\,
            lcout => \transmit_module.TX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i6_3_lut_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21613\,
            in1 => \N__16451\,
            in2 => \_gnd_net_\,
            in3 => \N__17015\,
            lcout => \transmit_module.n142\,
            ltout => \transmit_module.n142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i5_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__20870\,
            in1 => \N__20189\,
            in2 => \N__14840\,
            in3 => \N__16991\,
            lcout => \transmit_module.TX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i1_3_lut_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21611\,
            in1 => \N__16526\,
            in2 => \_gnd_net_\,
            in3 => \N__16551\,
            lcout => \transmit_module.n147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i6_4_lut_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15532\,
            in1 => \N__14959\,
            in2 => \N__14837\,
            in3 => \N__14982\,
            lcout => \transmit_module.video_signal_controller.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__15026\,
            in1 => \N__15460\,
            in2 => \N__15496\,
            in3 => \N__15083\,
            lcout => \transmit_module.video_signal_controller.n3333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1608_2_lut_rep_20_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15074\,
            in2 => \_gnd_net_\,
            in3 => \N__15053\,
            lcout => \transmit_module.video_signal_controller.n3626\,
            ltout => \transmit_module.video_signal_controller.n3626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2134_3_lut_4_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15492\,
            in1 => \N__15016\,
            in2 => \N__14987\,
            in3 => \N__14930\,
            lcout => \transmit_module.video_signal_controller.n3477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14984\,
            in2 => \_gnd_net_\,
            in3 => \N__15430\,
            lcout => \transmit_module.video_signal_controller.n3331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i11_3_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21585\,
            in1 => \N__16665\,
            in2 => \_gnd_net_\,
            in3 => \N__16610\,
            lcout => \transmit_module.n137\,
            ltout => \transmit_module.n137_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i10_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__20123\,
            in1 => \N__20824\,
            in2 => \N__14963\,
            in3 => \N__16642\,
            lcout => \transmit_module.TX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23131\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16553\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23397\,
            ce => \N__20444\,
            sr => \N__20186\
        );

    \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16667\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23397\,
            ce => \N__20444\,
            sr => \N__20186\
        );

    \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17021\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23397\,
            ce => \N__20444\,
            sr => \N__20186\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_27_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__14960\,
            in1 => \N__14929\,
            in2 => \N__15536\,
            in3 => \N__15503\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n7_adj_618_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i5_4_lut_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15497\,
            in1 => \N__15464\,
            in2 => \N__15449\,
            in3 => \N__15446\,
            lcout => \transmit_module.video_signal_controller.VGA_VISIBLE_N_580\,
            ltout => \transmit_module.video_signal_controller.VGA_VISIBLE_N_580_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15437\,
            in3 => \N__16736\,
            lcout => \transmit_module.VGA_VISIBLE_Y\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VS_67_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15434\,
            in1 => \N__15410\,
            in2 => \N__15401\,
            in3 => \N__15389\,
            lcout => \ADV_VSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i123_2_lut_4_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__16423\,
            in1 => \N__16399\,
            in2 => \N__20121\,
            in3 => \N__16361\,
            lcout => \transmit_module.n2167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.old_VGA_HS_40_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16362\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.old_VGA_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_HS_66_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__15356\,
            in1 => \N__15329\,
            in2 => \N__15320\,
            in3 => \N__15308\,
            lcout => \ADV_HSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i4_3_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21607\,
            in1 => \N__16469\,
            in2 => \_gnd_net_\,
            in3 => \N__16494\,
            lcout => \transmit_module.n144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i123_2_lut_4_lut_rep_30_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__16422\,
            in1 => \N__16398\,
            in2 => \N__20122\,
            in3 => \N__16360\,
            lcout => \transmit_module.n3636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i1_3_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20634\,
            in1 => \N__16439\,
            in2 => \_gnd_net_\,
            in3 => \N__16552\,
            lcout => \transmit_module.n116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i2_3_lut_rep_21_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16421\,
            in1 => \N__16397\,
            in2 => \_gnd_net_\,
            in3 => \N__16359\,
            lcout => \transmit_module.n3627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1619_4_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__16643\,
            in1 => \N__20015\,
            in2 => \N__20817\,
            in3 => \N__16334\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1603_4_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20769\,
            in1 => \N__16093\,
            in2 => \N__20163\,
            in3 => \N__16082\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i2_3_lut_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20655\,
            in1 => \N__18263\,
            in2 => \_gnd_net_\,
            in3 => \N__18295\,
            lcout => \transmit_module.n115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1610_4_lut_LC_14_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20878\,
            in1 => \N__15850\,
            in2 => \N__20328\,
            in3 => \N__15830\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i4_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24566\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i5_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15565\,
            lcout => \tvp_video_buffer.BUFFER_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i14_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16559\,
            lcout => \tvp_video_buffer.BUFFER_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i6_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16576\,
            lcout => \tvp_video_buffer.BUFFER_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_2_lut_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16544\,
            in2 => \N__19673\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n132\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \transmit_module.n3104\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_3_lut_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18288\,
            in3 => \N__16511\,
            lcout => \transmit_module.n131\,
            ltout => OPEN,
            carryin => \transmit_module.n3104\,
            carryout => \transmit_module.n3105\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_4_lut_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19215\,
            in3 => \N__16508\,
            lcout => \transmit_module.n130\,
            ltout => OPEN,
            carryin => \transmit_module.n3105\,
            carryout => \transmit_module.n3106\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_5_lut_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16493\,
            in3 => \N__16457\,
            lcout => \transmit_module.n129\,
            ltout => OPEN,
            carryin => \transmit_module.n3106\,
            carryout => \transmit_module.n3107\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_6_lut_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20523\,
            in3 => \N__16454\,
            lcout => \transmit_module.n128\,
            ltout => OPEN,
            carryin => \transmit_module.n3107\,
            carryout => \transmit_module.n3108\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_7_lut_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17020\,
            in3 => \N__16445\,
            lcout => \transmit_module.n127\,
            ltout => OPEN,
            carryin => \transmit_module.n3108\,
            carryout => \transmit_module.n3109\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_8_lut_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19262\,
            in3 => \N__16442\,
            lcout => \transmit_module.n126\,
            ltout => OPEN,
            carryin => \transmit_module.n3109\,
            carryout => \transmit_module.n3110\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_9_lut_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19328\,
            in3 => \N__16619\,
            lcout => \transmit_module.n125\,
            ltout => OPEN,
            carryin => \transmit_module.n3110\,
            carryout => \transmit_module.n3111\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_10_lut_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17271\,
            in3 => \N__16616\,
            lcout => \transmit_module.n124\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \transmit_module.n3112\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_11_lut_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19169\,
            in3 => \N__16613\,
            lcout => \transmit_module.n123\,
            ltout => OPEN,
            carryin => \transmit_module.n3112\,
            carryout => \transmit_module.n3113\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_12_lut_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16664\,
            in2 => \_gnd_net_\,
            in3 => \N__16604\,
            lcout => \transmit_module.n122\,
            ltout => OPEN,
            carryin => \transmit_module.n3113\,
            carryout => \transmit_module.n3114\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_13_lut_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24310\,
            in2 => \_gnd_net_\,
            in3 => \N__16601\,
            lcout => \transmit_module.n121\,
            ltout => OPEN,
            carryin => \transmit_module.n3114\,
            carryout => \transmit_module.n3115\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_14_lut_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23783\,
            in2 => \_gnd_net_\,
            in3 => \N__16598\,
            lcout => \transmit_module.n120\,
            ltout => OPEN,
            carryin => \transmit_module.n3115\,
            carryout => \transmit_module.n3116\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_15_lut_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23950\,
            in2 => \_gnd_net_\,
            in3 => \N__16595\,
            lcout => \transmit_module.n119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17264\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23393\,
            ce => \N__20455\,
            sr => \N__20352\
        );

    \transmit_module.BRAM_ADDR__i9_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__19142\,
            in1 => \N__20821\,
            in2 => \N__20286\,
            in3 => \N__19127\,
            lcout => \transmit_module.TX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i4_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20819\,
            in1 => \N__20171\,
            in2 => \N__20558\,
            in3 => \N__18238\,
            lcout => \transmit_module.TX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i8_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20820\,
            in1 => \N__20172\,
            in2 => \N__19601\,
            in3 => \N__19580\,
            lcout => \transmit_module.TX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i6_3_lut_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17027\,
            in1 => \N__20656\,
            in2 => \_gnd_net_\,
            in3 => \N__17016\,
            lcout => \transmit_module.n111\,
            ltout => \transmit_module.n111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1614_4_lut_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__20170\,
            in1 => \N__20818\,
            in2 => \N__16985\,
            in3 => \N__16982\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16742\,
            in1 => \N__16735\,
            in2 => \N__16721\,
            in3 => \N__16685\,
            lcout => \transmit_module.VGA_VISIBLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i11_3_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20652\,
            in1 => \N__16673\,
            in2 => \_gnd_net_\,
            in3 => \N__16666\,
            lcout => \transmit_module.n106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1_3_lut_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__20654\,
            in1 => \N__20179\,
            in2 => \_gnd_net_\,
            in3 => \N__20822\,
            lcout => \transmit_module.n2069\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1625_4_lut_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110010"
        )
    port map (
            in0 => \N__20823\,
            in1 => \N__20653\,
            in2 => \N__20287\,
            in3 => \N__21602\,
            lcout => \transmit_module.n2057\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i12_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18584\,
            in1 => \N__20770\,
            in2 => \_gnd_net_\,
            in3 => \N__16628\,
            lcout => \TX_ADDR_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => \N__17558\,
            sr => \N__20356\
        );

    \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18578\,
            in1 => \N__20772\,
            in2 => \_gnd_net_\,
            in3 => \N__17576\,
            lcout => \TX_ADDR_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => \N__17558\,
            sr => \N__20356\
        );

    \transmit_module.BRAM_ADDR__i13_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18593\,
            in1 => \N__20771\,
            in2 => \_gnd_net_\,
            in3 => \N__17567\,
            lcout => \TX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22937\,
            ce => \N__17558\,
            sr => \N__20356\
        );

    \transmit_module.mux_14_i9_3_lut_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21606\,
            in1 => \N__17272\,
            in2 => \_gnd_net_\,
            in3 => \N__17549\,
            lcout => \transmit_module.n139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i7_3_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21604\,
            in1 => \N__19272\,
            in2 => \_gnd_net_\,
            in3 => \N__17540\,
            lcout => \transmit_module.n141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i10_3_lut_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21603\,
            in1 => \N__19170\,
            in2 => \_gnd_net_\,
            in3 => \N__17531\,
            lcout => \transmit_module.n138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i8_3_lut_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21605\,
            in1 => \N__19334\,
            in2 => \_gnd_net_\,
            in3 => \N__17522\,
            lcout => \transmit_module.n140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1615_4_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20764\,
            in1 => \N__19237\,
            in2 => \N__20187\,
            in3 => \N__18418\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i9_3_lut_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20621\,
            in1 => \N__17285\,
            in2 => \_gnd_net_\,
            in3 => \N__17276\,
            lcout => \transmit_module.n108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1616_4_lut_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20765\,
            in1 => \N__19294\,
            in2 => \N__20188\,
            in3 => \N__18331\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19277\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22779\,
            ce => \N__20479\,
            sr => \N__20168\
        );

    \transmit_module.ADDR_Y_COMPONENT__i1_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18299\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22779\,
            ce => \N__20479\,
            sr => \N__20168\
        );

    \transmit_module.mux_14_i5_3_lut_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18257\,
            in1 => \N__21618\,
            in2 => \_gnd_net_\,
            in3 => \N__20516\,
            lcout => \transmit_module.n143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i3_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17807\,
            lcout => \RX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i12_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17813\,
            lcout => \tvp_video_buffer.BUFFER_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i13_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17801\,
            lcout => \tvp_video_buffer.BUFFER_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i4_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17795\,
            lcout => \RX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i5_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17693\,
            lcout => \RX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24572\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i6_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18431\,
            lcout => \RX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i7_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18454\,
            lcout => \tvp_video_buffer.BUFFER_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i15_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18437\,
            lcout => \tvp_video_buffer.BUFFER_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i6_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20868\,
            in1 => \N__19241\,
            in2 => \N__20353\,
            in3 => \N__18425\,
            lcout => \transmit_module.TX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i0_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21179\,
            lcout => \transmit_module.X_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23130\,
            ce => \N__21129\,
            sr => \N__18382\
        );

    \transmit_module.BRAM_ADDR__i7_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__19298\,
            in1 => \N__20237\,
            in2 => \N__20879\,
            in3 => \N__18338\,
            lcout => \transmit_module.TX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i3_3_lut_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19208\,
            in1 => \N__21614\,
            in2 => \_gnd_net_\,
            in3 => \N__18320\,
            lcout => \transmit_module.n145\,
            ltout => \transmit_module.n145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i2_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__20236\,
            in1 => \N__20871\,
            in2 => \N__18314\,
            in3 => \N__18889\,
            lcout => \transmit_module.TX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i16_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18626\,
            lcout => \transmit_module.Y_DELTA_PATTERN_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22700\,
            ce => \N__21062\,
            sr => \N__20239\
        );

    \transmit_module.Y_DELTA_PATTERN_i17_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18599\,
            lcout => \transmit_module.Y_DELTA_PATTERN_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22700\,
            ce => \N__21062\,
            sr => \N__20239\
        );

    \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18620\,
            lcout => \transmit_module.Y_DELTA_PATTERN_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23194\,
            ce => \N__21056\,
            sr => \N__20250\
        );

    \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18605\,
            lcout => \transmit_module.Y_DELTA_PATTERN_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23194\,
            ce => \N__21056\,
            sr => \N__20250\
        );

    \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19178\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => \N__20472\,
            sr => \N__20238\
        );

    \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19217\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => \N__20472\,
            sr => \N__20238\
        );

    \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23949\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => \N__20472\,
            sr => \N__20238\
        );

    \transmit_module.ADDR_Y_COMPONENT__i12_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23733\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => \N__20472\,
            sr => \N__20238\
        );

    \transmit_module.ADDR_Y_COMPONENT__i11_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24261\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => \N__20472\,
            sr => \N__20238\
        );

    \transmit_module.ADDR_Y_COMPONENT__i7_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19333\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22936\,
            ce => \N__20472\,
            sr => \N__20238\
        );

    \transmit_module.Y_DELTA_PATTERN_i0_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19610\,
            lcout => \transmit_module.Y_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23031\,
            ce => \N__21061\,
            sr => \N__20268\
        );

    \transmit_module.i1617_4_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20839\,
            in1 => \N__19591\,
            in2 => \N__20355\,
            in3 => \N__19576\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i8_3_lut_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20611\,
            in1 => \N__19343\,
            in2 => \_gnd_net_\,
            in3 => \N__19332\,
            lcout => \transmit_module.n109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i7_3_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20613\,
            in1 => \N__19283\,
            in2 => \_gnd_net_\,
            in3 => \N__19273\,
            lcout => \transmit_module.n110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i3_3_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20610\,
            in1 => \N__19226\,
            in2 => \_gnd_net_\,
            in3 => \N__19216\,
            lcout => \transmit_module.n114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i10_3_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20612\,
            in1 => \N__19187\,
            in2 => \_gnd_net_\,
            in3 => \N__19177\,
            lcout => \transmit_module.n107\,
            ltout => \transmit_module.n107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1618_4_lut_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20840\,
            in1 => \N__20305\,
            in2 => \N__19130\,
            in3 => \N__19123\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1611_4_lut_LC_16_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20876\,
            in1 => \N__18890\,
            in2 => \N__20407\,
            in3 => \N__18869\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i2_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18641\,
            lcout => \RX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19672\,
            lcout => \transmit_module.X_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23378\,
            ce => \N__21119\,
            sr => \N__21063\
        );

    \transmit_module.X_DELTA_PATTERN_i9_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19658\,
            lcout => \transmit_module.X_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23125\,
            ce => \N__21111\,
            sr => \N__21057\
        );

    \transmit_module.X_DELTA_PATTERN_i10_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19628\,
            lcout => \transmit_module.X_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23125\,
            ce => \N__21111\,
            sr => \N__21057\
        );

    \transmit_module.X_DELTA_PATTERN_i13_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19646\,
            lcout => \transmit_module.X_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23125\,
            ce => \N__21111\,
            sr => \N__21057\
        );

    \transmit_module.X_DELTA_PATTERN_i14_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19652\,
            lcout => \transmit_module.X_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23125\,
            ce => \N__21111\,
            sr => \N__21057\
        );

    \transmit_module.X_DELTA_PATTERN_i12_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19640\,
            lcout => \transmit_module.X_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23125\,
            ce => \N__21111\,
            sr => \N__21057\
        );

    \transmit_module.X_DELTA_PATTERN_i11_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19634\,
            lcout => \transmit_module.X_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23125\,
            ce => \N__21111\,
            sr => \N__21057\
        );

    \transmit_module.X_DELTA_PATTERN_i7_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19616\,
            lcout => \transmit_module.X_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23391\,
            ce => \N__21118\,
            sr => \N__21054\
        );

    \transmit_module.X_DELTA_PATTERN_i8_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19622\,
            lcout => \transmit_module.X_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23391\,
            ce => \N__21118\,
            sr => \N__21054\
        );

    \transmit_module.X_DELTA_PATTERN_i5_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21137\,
            lcout => \transmit_module.X_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23391\,
            ce => \N__21118\,
            sr => \N__21054\
        );

    \transmit_module.i2_3_lut_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20229\,
            in1 => \N__20841\,
            in2 => \_gnd_net_\,
            in3 => \N__21622\,
            lcout => \transmit_module.n2115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2176_3_lut_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20687\,
            in1 => \N__20669\,
            in2 => \_gnd_net_\,
            in3 => \N__24335\,
            lcout => \line_buffer.n3519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i5_3_lut_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20524\,
            in1 => \N__20620\,
            in2 => \_gnd_net_\,
            in3 => \N__20486\,
            lcout => \transmit_module.n112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i4_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23262\,
            ce => \N__20480\,
            sr => \N__20169\
        );

    \line_buffer.i2157_3_lut_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24373\,
            in1 => \N__19826\,
            in2 => \_gnd_net_\,
            in3 => \N__19811\,
            lcout => OPEN,
            ltout => \line_buffer.n3500_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2210_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__23827\,
            in1 => \N__24010\,
            in2 => \N__19796\,
            in3 => \N__19793\,
            lcout => OPEN,
            ltout => \line_buffer.n3537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i6_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__21239\,
            in1 => \N__21461\,
            in2 => \N__19781\,
            in3 => \N__24011\,
            lcout => \TX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2154_3_lut_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21272\,
            in1 => \N__21257\,
            in2 => \_gnd_net_\,
            in3 => \N__24385\,
            lcout => \line_buffer.n3497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2178_3_lut_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24384\,
            in1 => \N__21233\,
            in2 => \_gnd_net_\,
            in3 => \N__21215\,
            lcout => \line_buffer.n3521\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2182_3_lut_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21206\,
            in1 => \N__21188\,
            in2 => \_gnd_net_\,
            in3 => \N__24357\,
            lcout => \line_buffer.n3525\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i1_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21167\,
            lcout => \transmit_module.X_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23389\,
            ce => \N__21131\,
            sr => \N__21064\
        );

    \transmit_module.X_DELTA_PATTERN_i2_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21161\,
            lcout => \transmit_module.X_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23389\,
            ce => \N__21131\,
            sr => \N__21064\
        );

    \transmit_module.X_DELTA_PATTERN_i3_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21149\,
            lcout => \transmit_module.X_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23389\,
            ce => \N__21131\,
            sr => \N__21064\
        );

    \transmit_module.X_DELTA_PATTERN_i4_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21155\,
            lcout => \transmit_module.X_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23147\,
            ce => \N__21117\,
            sr => \N__21065\
        );

    \transmit_module.X_DELTA_PATTERN_i6_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21143\,
            lcout => \transmit_module.X_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23464\,
            ce => \N__21130\,
            sr => \N__21055\
        );

    \line_buffer.i2181_3_lut_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20909\,
            in1 => \N__20894\,
            in2 => \_gnd_net_\,
            in3 => \N__24367\,
            lcout => OPEN,
            ltout => \line_buffer.n3524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i5_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__23974\,
            in1 => \N__21530\,
            in2 => \N__21521\,
            in3 => \N__21725\,
            lcout => \TX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2215_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23826\,
            in1 => \N__22343\,
            in2 => \N__24009\,
            in3 => \N__21518\,
            lcout => OPEN,
            ltout => \line_buffer.n3555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i1_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__23997\,
            in1 => \N__24161\,
            in2 => \N__21509\,
            in3 => \N__21506\,
            lcout => \TX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2155_3_lut_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24341\,
            in1 => \N__21500\,
            in2 => \_gnd_net_\,
            in3 => \N__21482\,
            lcout => \line_buffer.n3498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2250_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24340\,
            in1 => \N__21455\,
            in2 => \N__23846\,
            in3 => \N__21446\,
            lcout => \line_buffer.n3597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i1_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21629\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n1814,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23019\,
            ce => 'H',
            sr => \N__24784\
        );

    \transmit_module.VGA_R__i2_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21386\,
            lcout => n1813,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23061\,
            ce => 'H',
            sr => \N__24796\
        );

    \transmit_module.VGA_R__i6_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21326\,
            lcout => n1809,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22772\,
            ce => 'H',
            sr => \N__24798\
        );

    \transmit_module.VGA_R__i7_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21878\,
            lcout => n1808,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22911\,
            ce => 'H',
            sr => \N__24797\
        );

    \line_buffer.i2145_3_lut_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24378\,
            in1 => \N__21815\,
            in2 => \_gnd_net_\,
            in3 => \N__21800\,
            lcout => \line_buffer.n3488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i7_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23998\,
            in1 => \N__21785\,
            in2 => \_gnd_net_\,
            in3 => \N__22037\,
            lcout => \TX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2146_3_lut_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24369\,
            in1 => \N__21776\,
            in2 => \_gnd_net_\,
            in3 => \N__21761\,
            lcout => \line_buffer.n3489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2220_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23819\,
            in1 => \N__21740\,
            in2 => \N__24008\,
            in3 => \N__21734\,
            lcout => \line_buffer.n3561\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2230_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24290\,
            in1 => \N__21719\,
            in2 => \N__23842\,
            in3 => \N__21704\,
            lcout => \line_buffer.n3573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3597_bdd_4_lut_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__21683\,
            in1 => \N__23833\,
            in2 => \N__21659\,
            in3 => \N__21638\,
            lcout => OPEN,
            ltout => \line_buffer.n3600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i0_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23996\,
            in2 => \N__21632\,
            in3 => \N__22286\,
            lcout => \TX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1118_1_lut_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21623\,
            lcout => \transmit_module.n2367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i8_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22220\,
            lcout => \ADV_B_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23123\,
            ce => 'H',
            sr => \N__24792\
        );

    \tvp_video_buffer.WIRE_OUT_i7_LC_20_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24728\,
            lcout => \RX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3585_bdd_4_lut_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__22073\,
            in1 => \N__23840\,
            in2 => \N__22055\,
            in3 => \N__24056\,
            lcout => \line_buffer.n3588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2225_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24337\,
            in1 => \N__22031\,
            in2 => \N__23849\,
            in3 => \N__22019\,
            lcout => \line_buffer.n3549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3549_bdd_4_lut_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__22004\,
            in1 => \N__23816\,
            in2 => \N__21989\,
            in3 => \N__21965\,
            lcout => OPEN,
            ltout => \line_buffer.n3552_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i2_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23986\,
            in2 => \N__21956\,
            in3 => \N__22469\,
            lcout => \TX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3573_bdd_4_lut_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__21953\,
            in1 => \N__23817\,
            in2 => \N__21938\,
            in3 => \N__21917\,
            lcout => \line_buffer.n3576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24344\,
            in1 => \N__21911\,
            in2 => \N__23844\,
            in3 => \N__21896\,
            lcout => OPEN,
            ltout => \line_buffer.n3603_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3603_bdd_4_lut_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__22502\,
            in1 => \N__22487\,
            in2 => \N__22472\,
            in3 => \N__23818\,
            lcout => \line_buffer.n3606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3543_bdd_4_lut_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__23831\,
            in1 => \N__22463\,
            in2 => \N__22448\,
            in3 => \N__23657\,
            lcout => OPEN,
            ltout => \line_buffer.n3546_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i4_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24016\,
            in2 => \N__22430\,
            in3 => \N__22427\,
            lcout => \TX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2235_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24368\,
            in1 => \N__22421\,
            in2 => \N__23847\,
            in3 => \N__22409\,
            lcout => \line_buffer.n3579\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2139_3_lut_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22400\,
            in1 => \N__22385\,
            in2 => \_gnd_net_\,
            in3 => \N__24380\,
            lcout => \line_buffer.n3482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2179_3_lut_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24379\,
            in1 => \N__22370\,
            in2 => \_gnd_net_\,
            in3 => \N__22358\,
            lcout => \line_buffer.n3522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3579_bdd_4_lut_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__22334\,
            in1 => \N__23832\,
            in2 => \N__22319\,
            in3 => \N__22295\,
            lcout => \line_buffer.n3582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i3_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22280\,
            lcout => n1812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22932\,
            ce => 'H',
            sr => \N__24785\
        );

    \transmit_module.VGA_R__i5_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24152\,
            lcout => n1810,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23092\,
            ce => 'H',
            sr => \N__24799\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2240_LC_21_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__24336\,
            in1 => \N__24086\,
            in2 => \N__23848\,
            in3 => \N__24071\,
            lcout => \line_buffer.n3585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2140_3_lut_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24377\,
            in1 => \N__24050\,
            in2 => \_gnd_net_\,
            in3 => \N__24032\,
            lcout => \line_buffer.n3483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__23845\,
            in1 => \N__24689\,
            in2 => \N__24017\,
            in3 => \N__23624\,
            lcout => OPEN,
            ltout => \line_buffer.n3567_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i3_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__24015\,
            in1 => \N__23888\,
            in2 => \N__23879\,
            in3 => \N__23876\,
            lcout => \TX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2205_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24342\,
            in1 => \N__23870\,
            in2 => \N__23843\,
            in3 => \N__23669\,
            lcout => \line_buffer.n3543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2137_3_lut_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__24343\,
            in1 => \N__23651\,
            in2 => \_gnd_net_\,
            in3 => \N__23636\,
            lcout => \line_buffer.n3480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i4_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23618\,
            lcout => n1811,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23184\,
            ce => 'H',
            sr => \N__24803\
        );

    \tvp_video_buffer.BUFFER_0__i16_LC_22_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24647\,
            lcout => \tvp_video_buffer.BUFFER_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2136_3_lut_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24719\,
            in1 => \N__24338\,
            in2 => \_gnd_net_\,
            in3 => \N__24704\,
            lcout => \line_buffer.n3479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i8_LC_23_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24664\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2175_3_lut_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24413\,
            in1 => \N__24401\,
            in2 => \_gnd_net_\,
            in3 => \N__24386\,
            lcout => \line_buffer.n3518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
