// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Oct 7 2018 19:45:30

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "main" view "INTERFACE"

module main (
    TVP_VIDEO,
    ADV_B,
    ADV_G,
    ADV_R,
    DEBUG,
    TVP_CLK,
    ADV_CLK,
    TVP_HSYNC,
    ADV_HSYNC,
    TVP_VSYNC,
    ADV_VSYNC,
    ADV_BLANK_N,
    LED,
    ADV_SYNC_N);

    input [9:0] TVP_VIDEO;
    output [7:0] ADV_B;
    output [7:0] ADV_G;
    output [7:0] ADV_R;
    inout [7:0] DEBUG;
    input TVP_CLK;
    output ADV_CLK;
    input TVP_HSYNC;
    output ADV_HSYNC;
    input TVP_VSYNC;
    output ADV_VSYNC;
    output ADV_BLANK_N;
    output LED;
    output ADV_SYNC_N;

    wire N__25265;
    wire N__25264;
    wire N__25263;
    wire N__25254;
    wire N__25253;
    wire N__25252;
    wire N__25245;
    wire N__25244;
    wire N__25243;
    wire N__25236;
    wire N__25235;
    wire N__25234;
    wire N__25227;
    wire N__25226;
    wire N__25225;
    wire N__25218;
    wire N__25217;
    wire N__25216;
    wire N__25209;
    wire N__25208;
    wire N__25207;
    wire N__25200;
    wire N__25199;
    wire N__25198;
    wire N__25191;
    wire N__25190;
    wire N__25189;
    wire N__25182;
    wire N__25181;
    wire N__25180;
    wire N__25173;
    wire N__25172;
    wire N__25171;
    wire N__25164;
    wire N__25163;
    wire N__25162;
    wire N__25155;
    wire N__25154;
    wire N__25153;
    wire N__25146;
    wire N__25145;
    wire N__25144;
    wire N__25137;
    wire N__25136;
    wire N__25135;
    wire N__25128;
    wire N__25127;
    wire N__25126;
    wire N__25119;
    wire N__25118;
    wire N__25117;
    wire N__25110;
    wire N__25109;
    wire N__25108;
    wire N__25101;
    wire N__25100;
    wire N__25099;
    wire N__25092;
    wire N__25091;
    wire N__25090;
    wire N__25083;
    wire N__25082;
    wire N__25081;
    wire N__25074;
    wire N__25073;
    wire N__25072;
    wire N__25065;
    wire N__25064;
    wire N__25063;
    wire N__25056;
    wire N__25055;
    wire N__25054;
    wire N__25047;
    wire N__25046;
    wire N__25045;
    wire N__25038;
    wire N__25037;
    wire N__25036;
    wire N__25029;
    wire N__25028;
    wire N__25027;
    wire N__25020;
    wire N__25019;
    wire N__25018;
    wire N__25011;
    wire N__25010;
    wire N__25009;
    wire N__25002;
    wire N__25001;
    wire N__25000;
    wire N__24993;
    wire N__24992;
    wire N__24991;
    wire N__24984;
    wire N__24983;
    wire N__24982;
    wire N__24975;
    wire N__24974;
    wire N__24973;
    wire N__24966;
    wire N__24965;
    wire N__24964;
    wire N__24957;
    wire N__24956;
    wire N__24955;
    wire N__24948;
    wire N__24947;
    wire N__24946;
    wire N__24939;
    wire N__24938;
    wire N__24937;
    wire N__24930;
    wire N__24929;
    wire N__24928;
    wire N__24921;
    wire N__24920;
    wire N__24919;
    wire N__24912;
    wire N__24911;
    wire N__24910;
    wire N__24903;
    wire N__24902;
    wire N__24901;
    wire N__24894;
    wire N__24893;
    wire N__24892;
    wire N__24885;
    wire N__24884;
    wire N__24883;
    wire N__24876;
    wire N__24875;
    wire N__24874;
    wire N__24867;
    wire N__24866;
    wire N__24865;
    wire N__24858;
    wire N__24857;
    wire N__24856;
    wire N__24849;
    wire N__24848;
    wire N__24847;
    wire N__24840;
    wire N__24839;
    wire N__24838;
    wire N__24831;
    wire N__24830;
    wire N__24829;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24799;
    wire N__24798;
    wire N__24797;
    wire N__24796;
    wire N__24795;
    wire N__24794;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24786;
    wire N__24785;
    wire N__24784;
    wire N__24781;
    wire N__24780;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24765;
    wire N__24764;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24749;
    wire N__24746;
    wire N__24745;
    wire N__24744;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24733;
    wire N__24732;
    wire N__24727;
    wire N__24724;
    wire N__24719;
    wire N__24716;
    wire N__24715;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24686;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24642;
    wire N__24641;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24625;
    wire N__24618;
    wire N__24613;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24523;
    wire N__24522;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24514;
    wire N__24513;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24505;
    wire N__24500;
    wire N__24497;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24489;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24474;
    wire N__24471;
    wire N__24470;
    wire N__24469;
    wire N__24468;
    wire N__24463;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24455;
    wire N__24454;
    wire N__24447;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24425;
    wire N__24424;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24412;
    wire N__24411;
    wire N__24410;
    wire N__24409;
    wire N__24408;
    wire N__24407;
    wire N__24404;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24378;
    wire N__24377;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24344;
    wire N__24343;
    wire N__24342;
    wire N__24339;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24323;
    wire N__24322;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24270;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24227;
    wire N__24220;
    wire N__24217;
    wire N__24210;
    wire N__24205;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24167;
    wire N__24166;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24162;
    wire N__24161;
    wire N__24160;
    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24156;
    wire N__24155;
    wire N__24154;
    wire N__24153;
    wire N__24152;
    wire N__24149;
    wire N__24148;
    wire N__24147;
    wire N__24146;
    wire N__24145;
    wire N__24144;
    wire N__24143;
    wire N__24142;
    wire N__24141;
    wire N__24140;
    wire N__24139;
    wire N__24138;
    wire N__24137;
    wire N__24136;
    wire N__24135;
    wire N__24134;
    wire N__24133;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24129;
    wire N__24128;
    wire N__24127;
    wire N__24126;
    wire N__24125;
    wire N__24124;
    wire N__24123;
    wire N__24122;
    wire N__24121;
    wire N__24120;
    wire N__24119;
    wire N__24118;
    wire N__24117;
    wire N__24116;
    wire N__24115;
    wire N__24114;
    wire N__24113;
    wire N__24112;
    wire N__24111;
    wire N__24110;
    wire N__24109;
    wire N__24108;
    wire N__24107;
    wire N__24106;
    wire N__24105;
    wire N__24104;
    wire N__24103;
    wire N__24102;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24098;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23945;
    wire N__23944;
    wire N__23941;
    wire N__23940;
    wire N__23939;
    wire N__23938;
    wire N__23937;
    wire N__23934;
    wire N__23933;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23920;
    wire N__23919;
    wire N__23918;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23891;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23864;
    wire N__23861;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23839;
    wire N__23836;
    wire N__23827;
    wire N__23822;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23791;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23738;
    wire N__23735;
    wire N__23734;
    wire N__23731;
    wire N__23730;
    wire N__23729;
    wire N__23728;
    wire N__23725;
    wire N__23724;
    wire N__23723;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23715;
    wire N__23714;
    wire N__23711;
    wire N__23710;
    wire N__23709;
    wire N__23708;
    wire N__23705;
    wire N__23704;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23689;
    wire N__23688;
    wire N__23687;
    wire N__23686;
    wire N__23681;
    wire N__23678;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23667;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23649;
    wire N__23648;
    wire N__23647;
    wire N__23646;
    wire N__23641;
    wire N__23638;
    wire N__23637;
    wire N__23636;
    wire N__23635;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23621;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23613;
    wire N__23608;
    wire N__23605;
    wire N__23604;
    wire N__23603;
    wire N__23602;
    wire N__23601;
    wire N__23600;
    wire N__23599;
    wire N__23598;
    wire N__23595;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23571;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23553;
    wire N__23552;
    wire N__23551;
    wire N__23550;
    wire N__23547;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23532;
    wire N__23531;
    wire N__23528;
    wire N__23527;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23488;
    wire N__23487;
    wire N__23486;
    wire N__23483;
    wire N__23482;
    wire N__23479;
    wire N__23478;
    wire N__23475;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23467;
    wire N__23466;
    wire N__23457;
    wire N__23452;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23440;
    wire N__23439;
    wire N__23436;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23418;
    wire N__23417;
    wire N__23414;
    wire N__23413;
    wire N__23410;
    wire N__23409;
    wire N__23406;
    wire N__23405;
    wire N__23404;
    wire N__23403;
    wire N__23400;
    wire N__23395;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23358;
    wire N__23357;
    wire N__23350;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23336;
    wire N__23335;
    wire N__23332;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23302;
    wire N__23299;
    wire N__23298;
    wire N__23295;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23278;
    wire N__23271;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23257;
    wire N__23254;
    wire N__23253;
    wire N__23250;
    wire N__23249;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23232;
    wire N__23229;
    wire N__23228;
    wire N__23227;
    wire N__23216;
    wire N__23213;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23201;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23184;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23157;
    wire N__23154;
    wire N__23149;
    wire N__23144;
    wire N__23137;
    wire N__23134;
    wire N__23133;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23125;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23083;
    wire N__23080;
    wire N__23075;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23051;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23039;
    wire N__23038;
    wire N__23037;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23023;
    wire N__23020;
    wire N__23015;
    wire N__23012;
    wire N__23003;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22987;
    wire N__22982;
    wire N__22979;
    wire N__22972;
    wire N__22969;
    wire N__22964;
    wire N__22961;
    wire N__22956;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22936;
    wire N__22931;
    wire N__22928;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22912;
    wire N__22909;
    wire N__22908;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22887;
    wire N__22880;
    wire N__22877;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22807;
    wire N__22800;
    wire N__22797;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22761;
    wire N__22758;
    wire N__22753;
    wire N__22746;
    wire N__22737;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22716;
    wire N__22707;
    wire N__22694;
    wire N__22693;
    wire N__22692;
    wire N__22689;
    wire N__22688;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22649;
    wire N__22646;
    wire N__22641;
    wire N__22634;
    wire N__22631;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22519;
    wire N__22518;
    wire N__22517;
    wire N__22514;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22483;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22445;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22423;
    wire N__22418;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22393;
    wire N__22392;
    wire N__22391;
    wire N__22390;
    wire N__22389;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22381;
    wire N__22378;
    wire N__22377;
    wire N__22376;
    wire N__22375;
    wire N__22374;
    wire N__22373;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22350;
    wire N__22347;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22339;
    wire N__22338;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22306;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22269;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22249;
    wire N__22242;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22200;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21955;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21475;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21431;
    wire N__21430;
    wire N__21429;
    wire N__21428;
    wire N__21427;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21407;
    wire N__21406;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21382;
    wire N__21381;
    wire N__21378;
    wire N__21373;
    wire N__21366;
    wire N__21363;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21355;
    wire N__21354;
    wire N__21351;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21322;
    wire N__21319;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21287;
    wire N__21278;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20965;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20879;
    wire N__20876;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20806;
    wire N__20805;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20773;
    wire N__20772;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20757;
    wire N__20752;
    wire N__20749;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20683;
    wire N__20682;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20676;
    wire N__20673;
    wire N__20672;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20661;
    wire N__20656;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20648;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20626;
    wire N__20625;
    wire N__20620;
    wire N__20615;
    wire N__20612;
    wire N__20605;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20579;
    wire N__20578;
    wire N__20577;
    wire N__20574;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20552;
    wire N__20549;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20263;
    wire N__20262;
    wire N__20261;
    wire N__20260;
    wire N__20259;
    wire N__20258;
    wire N__20257;
    wire N__20256;
    wire N__20255;
    wire N__20254;
    wire N__20253;
    wire N__20252;
    wire N__20251;
    wire N__20248;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20209;
    wire N__20206;
    wire N__20201;
    wire N__20196;
    wire N__20195;
    wire N__20194;
    wire N__20193;
    wire N__20190;
    wire N__20185;
    wire N__20182;
    wire N__20181;
    wire N__20180;
    wire N__20179;
    wire N__20172;
    wire N__20167;
    wire N__20164;
    wire N__20163;
    wire N__20162;
    wire N__20161;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20130;
    wire N__20129;
    wire N__20128;
    wire N__20127;
    wire N__20122;
    wire N__20119;
    wire N__20112;
    wire N__20109;
    wire N__20104;
    wire N__20091;
    wire N__20084;
    wire N__20069;
    wire N__20068;
    wire N__20067;
    wire N__20066;
    wire N__20065;
    wire N__20062;
    wire N__20061;
    wire N__20060;
    wire N__20059;
    wire N__20058;
    wire N__20057;
    wire N__20056;
    wire N__20055;
    wire N__20054;
    wire N__20051;
    wire N__20050;
    wire N__20049;
    wire N__20046;
    wire N__20045;
    wire N__20044;
    wire N__20043;
    wire N__20042;
    wire N__20041;
    wire N__20038;
    wire N__20037;
    wire N__20036;
    wire N__20035;
    wire N__20034;
    wire N__20033;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20019;
    wire N__20018;
    wire N__20017;
    wire N__20014;
    wire N__20013;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20007;
    wire N__20006;
    wire N__20003;
    wire N__20002;
    wire N__20001;
    wire N__19998;
    wire N__19997;
    wire N__19996;
    wire N__19995;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19964;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19952;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19935;
    wire N__19932;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19912;
    wire N__19911;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19876;
    wire N__19875;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19852;
    wire N__19849;
    wire N__19842;
    wire N__19839;
    wire N__19838;
    wire N__19837;
    wire N__19836;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19791;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19758;
    wire N__19751;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19739;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19727;
    wire N__19724;
    wire N__19723;
    wire N__19722;
    wire N__19721;
    wire N__19718;
    wire N__19709;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19694;
    wire N__19693;
    wire N__19692;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19674;
    wire N__19671;
    wire N__19660;
    wire N__19653;
    wire N__19638;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19616;
    wire N__19613;
    wire N__19612;
    wire N__19609;
    wire N__19608;
    wire N__19607;
    wire N__19604;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19586;
    wire N__19583;
    wire N__19568;
    wire N__19561;
    wire N__19552;
    wire N__19547;
    wire N__19540;
    wire N__19517;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19499;
    wire N__19496;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19481;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19264;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19213;
    wire N__19210;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19147;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19136;
    wire N__19135;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19120;
    wire N__19119;
    wire N__19112;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19082;
    wire N__19081;
    wire N__19078;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19056;
    wire N__19051;
    wire N__19048;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19035;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19021;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19006;
    wire N__19003;
    wire N__19002;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18963;
    wire N__18960;
    wire N__18959;
    wire N__18956;
    wire N__18951;
    wire N__18944;
    wire N__18941;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18925;
    wire N__18920;
    wire N__18919;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18908;
    wire N__18901;
    wire N__18898;
    wire N__18897;
    wire N__18896;
    wire N__18895;
    wire N__18894;
    wire N__18893;
    wire N__18892;
    wire N__18887;
    wire N__18880;
    wire N__18873;
    wire N__18872;
    wire N__18871;
    wire N__18870;
    wire N__18863;
    wire N__18862;
    wire N__18855;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18844;
    wire N__18843;
    wire N__18840;
    wire N__18835;
    wire N__18832;
    wire N__18827;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18798;
    wire N__18793;
    wire N__18790;
    wire N__18785;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18777;
    wire N__18772;
    wire N__18769;
    wire N__18768;
    wire N__18767;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18756;
    wire N__18755;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18737;
    wire N__18734;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18713;
    wire N__18710;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18686;
    wire N__18683;
    wire N__18682;
    wire N__18681;
    wire N__18680;
    wire N__18675;
    wire N__18670;
    wire N__18669;
    wire N__18666;
    wire N__18665;
    wire N__18664;
    wire N__18663;
    wire N__18662;
    wire N__18661;
    wire N__18660;
    wire N__18659;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18635;
    wire N__18632;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18592;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18581;
    wire N__18580;
    wire N__18579;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18558;
    wire N__18557;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18525;
    wire N__18520;
    wire N__18517;
    wire N__18512;
    wire N__18509;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18416;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18404;
    wire N__18401;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18389;
    wire N__18386;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18374;
    wire N__18371;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18359;
    wire N__18356;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18326;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18063;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__18001;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17920;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17890;
    wire N__17887;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17863;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17827;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17794;
    wire N__17791;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17625;
    wire N__17622;
    wire N__17619;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17570;
    wire N__17567;
    wire N__17566;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17556;
    wire N__17555;
    wire N__17554;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17542;
    wire N__17541;
    wire N__17538;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17517;
    wire N__17514;
    wire N__17513;
    wire N__17510;
    wire N__17505;
    wire N__17502;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17462;
    wire N__17461;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16846;
    wire N__16843;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16780;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16738;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16725;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16683;
    wire N__16680;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16657;
    wire N__16654;
    wire N__16651;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16594;
    wire N__16591;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16543;
    wire N__16540;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16464;
    wire N__16461;
    wire N__16458;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16425;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16405;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16128;
    wire N__16121;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16085;
    wire N__16084;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16074;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15853;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15832;
    wire N__15829;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15795;
    wire N__15792;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15496;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15379;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15367;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15343;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15255;
    wire N__15252;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15175;
    wire N__15174;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15156;
    wire N__15153;
    wire N__15146;
    wire N__15145;
    wire N__15144;
    wire N__15143;
    wire N__15142;
    wire N__15141;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15127;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15119;
    wire N__15116;
    wire N__15115;
    wire N__15114;
    wire N__15111;
    wire N__15106;
    wire N__15103;
    wire N__15098;
    wire N__15097;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15024;
    wire N__15019;
    wire N__15016;
    wire N__15015;
    wire N__15010;
    wire N__15007;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14992;
    wire N__14989;
    wire N__14988;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14923;
    wire N__14922;
    wire N__14921;
    wire N__14920;
    wire N__14919;
    wire N__14918;
    wire N__14917;
    wire N__14916;
    wire N__14913;
    wire N__14910;
    wire N__14903;
    wire N__14896;
    wire N__14893;
    wire N__14882;
    wire N__14881;
    wire N__14880;
    wire N__14879;
    wire N__14876;
    wire N__14869;
    wire N__14868;
    wire N__14867;
    wire N__14866;
    wire N__14865;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14847;
    wire N__14844;
    wire N__14839;
    wire N__14828;
    wire N__14827;
    wire N__14826;
    wire N__14825;
    wire N__14824;
    wire N__14823;
    wire N__14822;
    wire N__14821;
    wire N__14818;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14776;
    wire N__14771;
    wire N__14768;
    wire N__14753;
    wire N__14750;
    wire N__14749;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14706;
    wire N__14703;
    wire N__14698;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14578;
    wire N__14575;
    wire N__14574;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14539;
    wire N__14536;
    wire N__14535;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14523;
    wire N__14520;
    wire N__14513;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14503;
    wire N__14502;
    wire N__14499;
    wire N__14496;
    wire N__14493;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14461;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14451;
    wire N__14450;
    wire N__14443;
    wire N__14440;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14360;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14344;
    wire N__14341;
    wire N__14336;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14294;
    wire N__14291;
    wire N__14288;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14277;
    wire N__14274;
    wire N__14273;
    wire N__14270;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14247;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14212;
    wire N__14211;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14190;
    wire N__14187;
    wire N__14180;
    wire N__14177;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14165;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14114;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13895;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13834;
    wire N__13831;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13669;
    wire N__13666;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13615;
    wire N__13612;
    wire N__13609;
    wire N__13604;
    wire N__13601;
    wire N__13600;
    wire N__13597;
    wire N__13594;
    wire N__13591;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13534;
    wire N__13533;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13486;
    wire N__13483;
    wire N__13482;
    wire N__13479;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13414;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13404;
    wire N__13403;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13384;
    wire N__13381;
    wire N__13378;
    wire N__13375;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13309;
    wire N__13306;
    wire N__13305;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13293;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13268;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13219;
    wire N__13218;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13206;
    wire N__13199;
    wire N__13198;
    wire N__13195;
    wire N__13194;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13169;
    wire N__13166;
    wire N__13165;
    wire N__13164;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13152;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13135;
    wire N__13134;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13122;
    wire N__13115;
    wire N__13114;
    wire N__13111;
    wire N__13110;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13072;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13061;
    wire N__13054;
    wire N__13051;
    wire N__13048;
    wire N__13045;
    wire N__13040;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13028;
    wire N__13025;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13017;
    wire N__13016;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__12998;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12971;
    wire N__12970;
    wire N__12969;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12953;
    wire N__12952;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12913;
    wire N__12910;
    wire N__12907;
    wire N__12902;
    wire N__12901;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12890;
    wire N__12887;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12871;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12853;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12836;
    wire N__12835;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12811;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12794;
    wire N__12793;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12727;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12640;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12578;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12566;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12554;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12535;
    wire N__12534;
    wire N__12531;
    wire N__12526;
    wire N__12521;
    wire N__12520;
    wire N__12519;
    wire N__12516;
    wire N__12511;
    wire N__12506;
    wire N__12503;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12493;
    wire N__12490;
    wire N__12485;
    wire N__12484;
    wire N__12483;
    wire N__12480;
    wire N__12477;
    wire N__12474;
    wire N__12473;
    wire N__12468;
    wire N__12463;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12444;
    wire N__12439;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12416;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12408;
    wire N__12407;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12384;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12359;
    wire N__12356;
    wire N__12355;
    wire N__12352;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12103;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12043;
    wire N__12040;
    wire N__12037;
    wire N__12034;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__11998;
    wire N__11995;
    wire N__11992;
    wire N__11989;
    wire N__11986;
    wire N__11983;
    wire N__11980;
    wire N__11977;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11920;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11873;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11861;
    wire N__11860;
    wire N__11857;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11829;
    wire N__11826;
    wire N__11819;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11804;
    wire N__11801;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11767;
    wire N__11764;
    wire N__11761;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11686;
    wire N__11683;
    wire N__11680;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11555;
    wire N__11554;
    wire N__11549;
    wire N__11548;
    wire N__11545;
    wire N__11544;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11288;
    wire N__11285;
    wire N__11284;
    wire N__11283;
    wire N__11278;
    wire N__11275;
    wire N__11274;
    wire N__11271;
    wire N__11266;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11251;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11015;
    wire N__11014;
    wire N__11013;
    wire N__11010;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10964;
    wire N__10963;
    wire N__10962;
    wire N__10959;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10870;
    wire N__10865;
    wire N__10862;
    wire N__10861;
    wire N__10860;
    wire N__10857;
    wire N__10852;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10819;
    wire N__10818;
    wire N__10815;
    wire N__10810;
    wire N__10809;
    wire N__10808;
    wire N__10807;
    wire N__10804;
    wire N__10801;
    wire N__10794;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10728;
    wire N__10725;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10717;
    wire N__10716;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10708;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10689;
    wire N__10686;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10665;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10609;
    wire N__10606;
    wire N__10603;
    wire N__10602;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10596;
    wire N__10595;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10565;
    wire N__10560;
    wire N__10557;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10541;
    wire N__10536;
    wire N__10531;
    wire N__10528;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10500;
    wire N__10497;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10482;
    wire N__10477;
    wire N__10476;
    wire N__10475;
    wire N__10472;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10446;
    wire N__10439;
    wire N__10436;
    wire N__10431;
    wire N__10428;
    wire N__10423;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10399;
    wire N__10396;
    wire N__10395;
    wire N__10394;
    wire N__10391;
    wire N__10384;
    wire N__10379;
    wire N__10378;
    wire N__10377;
    wire N__10376;
    wire N__10373;
    wire N__10366;
    wire N__10361;
    wire N__10358;
    wire N__10357;
    wire N__10356;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10344;
    wire N__10341;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10327;
    wire N__10326;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10314;
    wire N__10311;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10294;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10264;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10220;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10132;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9988;
    wire N__9985;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9968;
    wire N__9965;
    wire N__9964;
    wire N__9961;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9920;
    wire N__9917;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9894;
    wire N__9893;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9865;
    wire N__9862;
    wire N__9861;
    wire N__9860;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9839;
    wire N__9838;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9824;
    wire N__9823;
    wire N__9822;
    wire N__9819;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9793;
    wire N__9790;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9743;
    wire N__9740;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9715;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9698;
    wire N__9697;
    wire N__9696;
    wire N__9693;
    wire N__9690;
    wire N__9687;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9631;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9516;
    wire N__9515;
    wire N__9514;
    wire N__9513;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9502;
    wire N__9499;
    wire N__9498;
    wire N__9497;
    wire N__9496;
    wire N__9495;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9485;
    wire N__9484;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9442;
    wire N__9435;
    wire N__9428;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9070;
    wire N__9069;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9058;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9027;
    wire N__9024;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9010;
    wire N__9007;
    wire N__9002;
    wire N__9001;
    wire N__8992;
    wire N__8989;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire VCCG0;
    wire GNDG0;
    wire \transmit_module.Y_DELTA_PATTERN_37 ;
    wire \transmit_module.Y_DELTA_PATTERN_36 ;
    wire \transmit_module.Y_DELTA_PATTERN_31 ;
    wire \transmit_module.Y_DELTA_PATTERN_32 ;
    wire \transmit_module.Y_DELTA_PATTERN_33 ;
    wire \transmit_module.Y_DELTA_PATTERN_38 ;
    wire \transmit_module.Y_DELTA_PATTERN_35 ;
    wire \transmit_module.Y_DELTA_PATTERN_34 ;
    wire \transmit_module.Y_DELTA_PATTERN_9 ;
    wire \transmit_module.Y_DELTA_PATTERN_8 ;
    wire \transmit_module.Y_DELTA_PATTERN_22 ;
    wire \transmit_module.Y_DELTA_PATTERN_21 ;
    wire \transmit_module.Y_DELTA_PATTERN_20 ;
    wire \transmit_module.Y_DELTA_PATTERN_19 ;
    wire \transmit_module.Y_DELTA_PATTERN_18 ;
    wire \transmit_module.Y_DELTA_PATTERN_15 ;
    wire \transmit_module.Y_DELTA_PATTERN_23 ;
    wire \transmit_module.Y_DELTA_PATTERN_17 ;
    wire \transmit_module.Y_DELTA_PATTERN_16 ;
    wire \transmit_module.Y_DELTA_PATTERN_14 ;
    wire \transmit_module.Y_DELTA_PATTERN_39 ;
    wire \transmit_module.Y_DELTA_PATTERN_41 ;
    wire \transmit_module.Y_DELTA_PATTERN_40 ;
    wire \transmit_module.Y_DELTA_PATTERN_13 ;
    wire \transmit_module.Y_DELTA_PATTERN_12 ;
    wire \transmit_module.Y_DELTA_PATTERN_7 ;
    wire \transmit_module.Y_DELTA_PATTERN_6 ;
    wire \transmit_module.Y_DELTA_PATTERN_11 ;
    wire \transmit_module.Y_DELTA_PATTERN_10 ;
    wire \transmit_module.Y_DELTA_PATTERN_73 ;
    wire \transmit_module.Y_DELTA_PATTERN_72 ;
    wire \transmit_module.Y_DELTA_PATTERN_63 ;
    wire \transmit_module.Y_DELTA_PATTERN_71 ;
    wire \transmit_module.Y_DELTA_PATTERN_70 ;
    wire \transmit_module.Y_DELTA_PATTERN_66 ;
    wire \transmit_module.Y_DELTA_PATTERN_67 ;
    wire \transmit_module.Y_DELTA_PATTERN_65 ;
    wire \transmit_module.Y_DELTA_PATTERN_64 ;
    wire \transmit_module.Y_DELTA_PATTERN_69 ;
    wire \transmit_module.Y_DELTA_PATTERN_68 ;
    wire \transmit_module.Y_DELTA_PATTERN_24 ;
    wire \transmit_module.Y_DELTA_PATTERN_25 ;
    wire \transmit_module.Y_DELTA_PATTERN_43 ;
    wire \transmit_module.Y_DELTA_PATTERN_42 ;
    wire \transmit_module.Y_DELTA_PATTERN_44 ;
    wire \transmit_module.Y_DELTA_PATTERN_45 ;
    wire DEBUG_c_5_c;
    wire RX_DATA_3;
    wire \tvp_video_buffer.BUFFER_0_5 ;
    wire \tvp_video_buffer.BUFFER_1_5 ;
    wire n27;
    wire \line_buffer.n603 ;
    wire \line_buffer.n595 ;
    wire \line_buffer.n602 ;
    wire \line_buffer.n594 ;
    wire TVP_VIDEO_c_2;
    wire \transmit_module.Y_DELTA_PATTERN_74 ;
    wire \transmit_module.Y_DELTA_PATTERN_75 ;
    wire \transmit_module.Y_DELTA_PATTERN_78 ;
    wire \transmit_module.Y_DELTA_PATTERN_79 ;
    wire \transmit_module.Y_DELTA_PATTERN_77 ;
    wire \transmit_module.Y_DELTA_PATTERN_76 ;
    wire \transmit_module.Y_DELTA_PATTERN_62 ;
    wire \transmit_module.Y_DELTA_PATTERN_61 ;
    wire \transmit_module.Y_DELTA_PATTERN_80 ;
    wire \transmit_module.Y_DELTA_PATTERN_82 ;
    wire \transmit_module.Y_DELTA_PATTERN_81 ;
    wire \transmit_module.Y_DELTA_PATTERN_83 ;
    wire \transmit_module.Y_DELTA_PATTERN_85 ;
    wire \transmit_module.Y_DELTA_PATTERN_84 ;
    wire \transmit_module.Y_DELTA_PATTERN_26 ;
    wire \transmit_module.Y_DELTA_PATTERN_27 ;
    wire \transmit_module.Y_DELTA_PATTERN_28 ;
    wire \transmit_module.Y_DELTA_PATTERN_30 ;
    wire \transmit_module.Y_DELTA_PATTERN_29 ;
    wire \transmit_module.Y_DELTA_PATTERN_47 ;
    wire \transmit_module.Y_DELTA_PATTERN_46 ;
    wire \transmit_module.Y_DELTA_PATTERN_49 ;
    wire \transmit_module.Y_DELTA_PATTERN_48 ;
    wire \transmit_module.Y_DELTA_PATTERN_53 ;
    wire \transmit_module.Y_DELTA_PATTERN_52 ;
    wire \transmit_module.Y_DELTA_PATTERN_51 ;
    wire \transmit_module.Y_DELTA_PATTERN_50 ;
    wire \transmit_module.Y_DELTA_PATTERN_60 ;
    wire \transmit_module.Y_DELTA_PATTERN_59 ;
    wire \transmit_module.Y_DELTA_PATTERN_58 ;
    wire \transmit_module.Y_DELTA_PATTERN_54 ;
    wire \transmit_module.Y_DELTA_PATTERN_55 ;
    wire \transmit_module.Y_DELTA_PATTERN_57 ;
    wire \transmit_module.Y_DELTA_PATTERN_56 ;
    wire \transmit_module.Y_DELTA_PATTERN_86 ;
    wire \transmit_module.Y_DELTA_PATTERN_96 ;
    wire \transmit_module.Y_DELTA_PATTERN_99 ;
    wire \transmit_module.Y_DELTA_PATTERN_98 ;
    wire \transmit_module.Y_DELTA_PATTERN_97 ;
    wire \transmit_module.Y_DELTA_PATTERN_95 ;
    wire \transmit_module.n3683 ;
    wire \transmit_module.video_signal_controller.n6_cascade_ ;
    wire \transmit_module.ADDR_Y_COMPONENT_11 ;
    wire \transmit_module.ADDR_Y_COMPONENT_12 ;
    wire bfn_11_17_0_;
    wire \transmit_module.video_signal_controller.n3183 ;
    wire \transmit_module.video_signal_controller.n3184 ;
    wire \transmit_module.video_signal_controller.n3185 ;
    wire \transmit_module.video_signal_controller.n3186 ;
    wire \transmit_module.video_signal_controller.n3187 ;
    wire \transmit_module.video_signal_controller.n3188 ;
    wire \transmit_module.video_signal_controller.n3189 ;
    wire \transmit_module.video_signal_controller.n3190 ;
    wire bfn_11_18_0_;
    wire \transmit_module.video_signal_controller.n3191 ;
    wire \transmit_module.video_signal_controller.n3192 ;
    wire \transmit_module.video_signal_controller.n3193 ;
    wire \tvp_video_buffer.BUFFER_0_2 ;
    wire TVP_VIDEO_c_3;
    wire \tvp_video_buffer.BUFFER_0_3 ;
    wire \transmit_module.X_DELTA_PATTERN_15 ;
    wire \transmit_module.X_DELTA_PATTERN_14 ;
    wire \transmit_module.Y_DELTA_PATTERN_94 ;
    wire \transmit_module.Y_DELTA_PATTERN_93 ;
    wire \transmit_module.Y_DELTA_PATTERN_92 ;
    wire \transmit_module.Y_DELTA_PATTERN_87 ;
    wire \transmit_module.Y_DELTA_PATTERN_89 ;
    wire \transmit_module.Y_DELTA_PATTERN_88 ;
    wire \transmit_module.Y_DELTA_PATTERN_91 ;
    wire \transmit_module.Y_DELTA_PATTERN_90 ;
    wire \transmit_module.n2209 ;
    wire bfn_12_14_0_;
    wire \transmit_module.video_signal_controller.n3194 ;
    wire \transmit_module.video_signal_controller.n3195 ;
    wire \transmit_module.video_signal_controller.n3196 ;
    wire \transmit_module.video_signal_controller.n3197 ;
    wire \transmit_module.video_signal_controller.n3198 ;
    wire \transmit_module.video_signal_controller.n3199 ;
    wire \transmit_module.video_signal_controller.VGA_Y_7 ;
    wire \transmit_module.video_signal_controller.n3200 ;
    wire \transmit_module.video_signal_controller.n3201 ;
    wire \transmit_module.video_signal_controller.VGA_Y_8 ;
    wire bfn_12_15_0_;
    wire \transmit_module.video_signal_controller.n3202 ;
    wire \transmit_module.video_signal_controller.n3203 ;
    wire \transmit_module.video_signal_controller.n3204 ;
    wire \transmit_module.video_signal_controller.VGA_Y_11 ;
    wire \transmit_module.video_signal_controller.VGA_Y_10 ;
    wire \transmit_module.video_signal_controller.VGA_Y_5 ;
    wire \transmit_module.video_signal_controller.n3485_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_6 ;
    wire \transmit_module.video_signal_controller.n3676 ;
    wire \transmit_module.video_signal_controller.VGA_Y_9 ;
    wire \transmit_module.video_signal_controller.n3464_cascade_ ;
    wire \transmit_module.video_signal_controller.n3378 ;
    wire \transmit_module.ADDR_Y_COMPONENT_5 ;
    wire \transmit_module.video_signal_controller.VGA_Y_3 ;
    wire \transmit_module.video_signal_controller.n6_adj_622 ;
    wire \transmit_module.video_signal_controller.VGA_Y_4 ;
    wire \transmit_module.video_signal_controller.n2019 ;
    wire \transmit_module.video_signal_controller.n2050 ;
    wire \transmit_module.video_signal_controller.n2050_cascade_ ;
    wire \transmit_module.video_signal_controller.n2398 ;
    wire \transmit_module.video_signal_controller.VGA_X_3 ;
    wire \transmit_module.video_signal_controller.VGA_X_4 ;
    wire \transmit_module.video_signal_controller.VGA_X_6 ;
    wire \transmit_module.video_signal_controller.n3482_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_5 ;
    wire \transmit_module.video_signal_controller.n55 ;
    wire \transmit_module.video_signal_controller.n3478_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_7 ;
    wire \transmit_module.video_signal_controller.VGA_X_0 ;
    wire \transmit_module.ADDR_Y_COMPONENT_13 ;
    wire \transmit_module.n2073 ;
    wire n20;
    wire \tvp_video_buffer.BUFFER_1_2 ;
    wire RX_DATA_0;
    wire TVP_VIDEO_c_4;
    wire \tvp_video_buffer.BUFFER_0_4 ;
    wire TVP_VIDEO_c_8;
    wire \tvp_video_buffer.BUFFER_1_3 ;
    wire RX_DATA_1;
    wire \tvp_video_buffer.BUFFER_1_4 ;
    wire RX_DATA_2;
    wire \tvp_video_buffer.BUFFER_0_8 ;
    wire \tvp_video_buffer.BUFFER_1_8 ;
    wire bfn_13_9_0_;
    wire \receive_module.rx_counter.n3210 ;
    wire \receive_module.rx_counter.n3211 ;
    wire \receive_module.rx_counter.n3212 ;
    wire \receive_module.rx_counter.n3213 ;
    wire \receive_module.rx_counter.n3214 ;
    wire \receive_module.rx_counter.n3215 ;
    wire \receive_module.rx_counter.n3216 ;
    wire \receive_module.rx_counter.n3217 ;
    wire bfn_13_10_0_;
    wire \receive_module.rx_counter.n3218 ;
    wire bfn_13_11_0_;
    wire \receive_module.rx_counter.n3175 ;
    wire \receive_module.rx_counter.n3176 ;
    wire \receive_module.rx_counter.n3177 ;
    wire \receive_module.rx_counter.n3178 ;
    wire \receive_module.rx_counter.n3179 ;
    wire \receive_module.rx_counter.n3180 ;
    wire \receive_module.rx_counter.n3181 ;
    wire \receive_module.rx_counter.n3182 ;
    wire bfn_13_12_0_;
    wire \receive_module.rx_counter.n10 ;
    wire \receive_module.rx_counter.n14_cascade_ ;
    wire \line_buffer.n539 ;
    wire \line_buffer.n531 ;
    wire \transmit_module.old_VGA_HS ;
    wire \transmit_module.ADDR_Y_COMPONENT_7 ;
    wire \transmit_module.video_signal_controller.n7 ;
    wire ADV_HSYNC_c;
    wire \transmit_module.n141_cascade_ ;
    wire n22;
    wire \transmit_module.VGA_VISIBLE_Y ;
    wire \transmit_module.n140 ;
    wire \transmit_module.n140_cascade_ ;
    wire \transmit_module.n109 ;
    wire n21;
    wire \transmit_module.video_signal_controller.VGA_Y_1 ;
    wire \transmit_module.video_signal_controller.n3520 ;
    wire \transmit_module.video_signal_controller.VGA_Y_0 ;
    wire \transmit_module.video_signal_controller.VGA_Y_2 ;
    wire \transmit_module.video_signal_controller.n2958 ;
    wire \transmit_module.video_signal_controller.n2975 ;
    wire \transmit_module.n142 ;
    wire \transmit_module.n142_cascade_ ;
    wire \transmit_module.n111 ;
    wire n23;
    wire \transmit_module.video_signal_controller.n3366 ;
    wire \transmit_module.video_signal_controller.VGA_X_8 ;
    wire \transmit_module.video_signal_controller.n2017 ;
    wire \transmit_module.video_signal_controller.n3007_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_VISIBLE_N_588 ;
    wire \transmit_module.n143 ;
    wire \transmit_module.n143_cascade_ ;
    wire n24;
    wire \transmit_module.video_signal_controller.VGA_X_10 ;
    wire \transmit_module.video_signal_controller.n3007 ;
    wire \transmit_module.video_signal_controller.VGA_X_2 ;
    wire \transmit_module.video_signal_controller.VGA_X_1 ;
    wire \transmit_module.video_signal_controller.n3679 ;
    wire \transmit_module.n108 ;
    wire \transmit_module.video_signal_controller.VGA_X_9 ;
    wire \transmit_module.video_signal_controller.n6_adj_623 ;
    wire \transmit_module.n139 ;
    wire \transmit_module.n138_cascade_ ;
    wire n19;
    wire \line_buffer.n3531 ;
    wire \line_buffer.n3530 ;
    wire \line_buffer.n3620 ;
    wire \line_buffer.n571 ;
    wire \line_buffer.n563 ;
    wire \line_buffer.n3534 ;
    wire TX_DATA_7;
    wire ADV_B_c;
    wire \line_buffer.n474 ;
    wire \line_buffer.n466 ;
    wire \line_buffer.n3533 ;
    wire \line_buffer.n542 ;
    wire \receive_module.rx_counter.X_1 ;
    wire \receive_module.rx_counter.X_0 ;
    wire \receive_module.rx_counter.X_2 ;
    wire \receive_module.rx_counter.n3225_cascade_ ;
    wire \receive_module.rx_counter.n3458_cascade_ ;
    wire \receive_module.rx_counter.X_4 ;
    wire \receive_module.rx_counter.X_6 ;
    wire \receive_module.rx_counter.n3 ;
    wire \receive_module.rx_counter.X_3 ;
    wire \receive_module.rx_counter.X_5 ;
    wire \receive_module.rx_counter.X_7 ;
    wire \receive_module.rx_counter.n6 ;
    wire \receive_module.rx_counter.n7_cascade_ ;
    wire \receive_module.rx_counter.n3225 ;
    wire \receive_module.rx_counter.old_HS ;
    wire \receive_module.rx_counter.n2081 ;
    wire \line_buffer.n573 ;
    wire \receive_module.rx_counter.n3429 ;
    wire \receive_module.rx_counter.X_8 ;
    wire \receive_module.rx_counter.X_9 ;
    wire \receive_module.rx_counter.n39 ;
    wire \receive_module.rx_counter.Y_6 ;
    wire \receive_module.rx_counter.Y_5 ;
    wire \receive_module.rx_counter.n5_cascade_ ;
    wire \receive_module.rx_counter.Y_7 ;
    wire \receive_module.rx_counter.n3455_cascade_ ;
    wire \receive_module.rx_counter.n3680 ;
    wire \receive_module.rx_counter.Y_8 ;
    wire \receive_module.rx_counter.n3481 ;
    wire \receive_module.rx_counter.n4_adj_612_cascade_ ;
    wire \receive_module.rx_counter.n54 ;
    wire \receive_module.rx_counter.Y_1 ;
    wire \receive_module.rx_counter.Y_0 ;
    wire \receive_module.rx_counter.Y_2 ;
    wire \receive_module.rx_counter.n3453 ;
    wire \receive_module.rx_counter.Y_3 ;
    wire \receive_module.rx_counter.Y_4 ;
    wire \receive_module.rx_counter.n4 ;
    wire RX_TX_SYNC;
    wire \line_buffer.n477 ;
    wire \line_buffer.n541 ;
    wire \line_buffer.n605 ;
    wire \line_buffer.n568 ;
    wire \line_buffer.n560 ;
    wire \sync_buffer.BUFFER_0_0 ;
    wire \transmit_module.ADDR_Y_COMPONENT_6 ;
    wire bfn_14_15_0_;
    wire \transmit_module.n131 ;
    wire \transmit_module.n3162 ;
    wire \transmit_module.n3163 ;
    wire \transmit_module.n3164 ;
    wire \transmit_module.n128 ;
    wire \transmit_module.n3165 ;
    wire \transmit_module.TX_ADDR_5 ;
    wire \transmit_module.n127 ;
    wire \transmit_module.n3166 ;
    wire \transmit_module.n126 ;
    wire \transmit_module.n3167 ;
    wire \transmit_module.TX_ADDR_7 ;
    wire \transmit_module.n125 ;
    wire \transmit_module.n3168 ;
    wire \transmit_module.n3169 ;
    wire \transmit_module.n124 ;
    wire bfn_14_16_0_;
    wire \transmit_module.n123 ;
    wire \transmit_module.n3170 ;
    wire \transmit_module.n3171 ;
    wire \transmit_module.n121 ;
    wire \transmit_module.n3172 ;
    wire \transmit_module.n120 ;
    wire \transmit_module.n3173 ;
    wire \transmit_module.n3174 ;
    wire \transmit_module.n119 ;
    wire \transmit_module.n112 ;
    wire \transmit_module.n146 ;
    wire \sync_buffer.BUFFER_1_0 ;
    wire RX_TX_SYNC_BUFF;
    wire \transmit_module.n122 ;
    wire \transmit_module.n137_cascade_ ;
    wire \transmit_module.n138 ;
    wire \transmit_module.video_signal_controller.n3382 ;
    wire \transmit_module.video_signal_controller.n3017 ;
    wire \transmit_module.video_signal_controller.VGA_X_11 ;
    wire \transmit_module.video_signal_controller.n7_adj_624 ;
    wire \transmit_module.n132 ;
    wire \transmit_module.ADDR_Y_COMPONENT_9 ;
    wire \transmit_module.TX_ADDR_9 ;
    wire \transmit_module.n107 ;
    wire \transmit_module.n115 ;
    wire \transmit_module.n116 ;
    wire \transmit_module.n116_cascade_ ;
    wire \transmit_module.n147 ;
    wire n28;
    wire \transmit_module.n106 ;
    wire \transmit_module.n137 ;
    wire n18;
    wire \transmit_module.TX_ADDR_10 ;
    wire \transmit_module.ADDR_Y_COMPONENT_10 ;
    wire \transmit_module.TX_ADDR_8 ;
    wire \transmit_module.ADDR_Y_COMPONENT_8 ;
    wire \transmit_module.TX_ADDR_1 ;
    wire \transmit_module.ADDR_Y_COMPONENT_1 ;
    wire \transmit_module.TX_ADDR_0 ;
    wire \transmit_module.ADDR_Y_COMPONENT_0 ;
    wire DEBUG_c_1_c;
    wire DEBUG_c_6_c;
    wire \tvp_vs_buffer.BUFFER_0_0 ;
    wire \tvp_video_buffer.BUFFER_0_6 ;
    wire TVP_HSYNC_buff;
    wire \transmit_module.X_DELTA_PATTERN_10 ;
    wire \transmit_module.X_DELTA_PATTERN_9 ;
    wire \transmit_module.X_DELTA_PATTERN_11 ;
    wire \transmit_module.X_DELTA_PATTERN_13 ;
    wire \transmit_module.X_DELTA_PATTERN_12 ;
    wire bfn_15_11_0_;
    wire \receive_module.n3149 ;
    wire \receive_module.n3150 ;
    wire \receive_module.n3151 ;
    wire \receive_module.n3152 ;
    wire \receive_module.n3153 ;
    wire \receive_module.n3154 ;
    wire \receive_module.n3155 ;
    wire \receive_module.n3156 ;
    wire bfn_15_12_0_;
    wire \receive_module.n3157 ;
    wire \receive_module.n3158 ;
    wire \receive_module.n3159 ;
    wire \receive_module.n3160 ;
    wire \receive_module.n3161 ;
    wire \line_buffer.n606 ;
    wire \line_buffer.n476 ;
    wire \receive_module.n3674 ;
    wire RX_ADDR_11;
    wire RX_ADDR_12;
    wire RX_ADDR_13;
    wire \line_buffer.n574 ;
    wire \tvp_vs_buffer.BUFFER_1_0 ;
    wire \tvp_vs_buffer.BUFFER_2_0 ;
    wire \transmit_module.X_DELTA_PATTERN_0 ;
    wire \transmit_module.X_DELTA_PATTERN_1 ;
    wire \transmit_module.X_DELTA_PATTERN_8 ;
    wire \transmit_module.X_DELTA_PATTERN_2 ;
    wire \transmit_module.X_DELTA_PATTERN_3 ;
    wire \transmit_module.X_DELTA_PATTERN_7 ;
    wire \transmit_module.X_DELTA_PATTERN_4 ;
    wire \transmit_module.n129 ;
    wire \transmit_module.n110 ;
    wire \transmit_module.n141 ;
    wire \transmit_module.TX_ADDR_6 ;
    wire \transmit_module.VGA_VISIBLE ;
    wire \transmit_module.n130 ;
    wire \transmit_module.n145_cascade_ ;
    wire \transmit_module.Y_DELTA_PATTERN_2 ;
    wire \transmit_module.Y_DELTA_PATTERN_5 ;
    wire \transmit_module.Y_DELTA_PATTERN_4 ;
    wire \transmit_module.Y_DELTA_PATTERN_3 ;
    wire \transmit_module.Y_DELTA_PATTERN_1 ;
    wire \receive_module.n136 ;
    wire RX_ADDR_1;
    wire \receive_module.n135 ;
    wire RX_ADDR_2;
    wire \receive_module.n133 ;
    wire RX_ADDR_4;
    wire \receive_module.n132 ;
    wire RX_ADDR_5;
    wire \receive_module.n131 ;
    wire RX_ADDR_6;
    wire \receive_module.n130 ;
    wire RX_ADDR_7;
    wire \transmit_module.ADDR_Y_COMPONENT_3 ;
    wire \transmit_module.TX_ADDR_3 ;
    wire \receive_module.n128 ;
    wire RX_ADDR_9;
    wire GB_BUFFER_DEBUG_c_3_c_THRU_CO;
    wire n1821;
    wire \receive_module.n129 ;
    wire RX_ADDR_8;
    wire \receive_module.n137 ;
    wire RX_ADDR_0;
    wire \receive_module.n134 ;
    wire RX_ADDR_3;
    wire \receive_module.n127 ;
    wire RX_ADDR_10;
    wire \receive_module.n3677 ;
    wire LED_c;
    wire PULSE_1HZ;
    wire \receive_module.rx_counter.old_VS ;
    wire \receive_module.rx_counter.n3522_cascade_ ;
    wire \receive_module.rx_counter.n7_adj_619 ;
    wire \receive_module.rx_counter.n11 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_0 ;
    wire bfn_16_10_0_;
    wire \receive_module.rx_counter.FRAME_COUNTER_1 ;
    wire \receive_module.rx_counter.n3205 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_2 ;
    wire \receive_module.rx_counter.n3206 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_3 ;
    wire \receive_module.rx_counter.n3207 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_4 ;
    wire \receive_module.rx_counter.n3208 ;
    wire \receive_module.rx_counter.n3209 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_5 ;
    wire \receive_module.rx_counter.n3675 ;
    wire \receive_module.rx_counter.n2550 ;
    wire \tvp_video_buffer.BUFFER_1_6 ;
    wire RX_DATA_6;
    wire RX_DATA_4;
    wire \receive_module.sync_wd.n6_cascade_ ;
    wire \receive_module.sync_wd.n4_cascade_ ;
    wire TVP_VSYNC_buff;
    wire DEBUG_c_0;
    wire DEBUG_c_4;
    wire \receive_module.sync_wd.old_visible ;
    wire RX_DATA_7;
    wire \line_buffer.n569 ;
    wire \line_buffer.n561 ;
    wire \line_buffer.n567 ;
    wire \line_buffer.n559 ;
    wire \transmit_module.TX_ADDR_4 ;
    wire \transmit_module.ADDR_Y_COMPONENT_4 ;
    wire \transmit_module.n2313 ;
    wire \transmit_module.ADDR_Y_COMPONENT_2 ;
    wire \transmit_module.Y_DELTA_PATTERN_0 ;
    wire \transmit_module.TX_ADDR_2 ;
    wire \transmit_module.n114 ;
    wire \transmit_module.n145 ;
    wire n26;
    wire \line_buffer.n535 ;
    wire \line_buffer.n527 ;
    wire \transmit_module.n3678 ;
    wire ADV_VSYNC_c;
    wire \transmit_module.n113 ;
    wire \transmit_module.n144 ;
    wire n25;
    wire n1818;
    wire \line_buffer.n470 ;
    wire \line_buffer.n462 ;
    wire \line_buffer.n3590 ;
    wire \line_buffer.n3593_cascade_ ;
    wire \line_buffer.n3629 ;
    wire TX_DATA_3;
    wire \line_buffer.n471 ;
    wire \line_buffer.n463 ;
    wire \line_buffer.n3552 ;
    wire \line_buffer.n3551_cascade_ ;
    wire \line_buffer.n600 ;
    wire \line_buffer.n592 ;
    wire TX_DATA_4;
    wire n1817;
    wire TX_DATA_1;
    wire n1820;
    wire \tvp_hs_buffer.BUFFER_1_0 ;
    wire \line_buffer.n536 ;
    wire \line_buffer.n528 ;
    wire \line_buffer.n534 ;
    wire \line_buffer.n526 ;
    wire \transmit_module.X_DELTA_PATTERN_6 ;
    wire \transmit_module.X_DELTA_PATTERN_5 ;
    wire \transmit_module.n2087 ;
    wire \transmit_module.n3682 ;
    wire \line_buffer.n533 ;
    wire \line_buffer.n525 ;
    wire \line_buffer.n3653 ;
    wire \line_buffer.n468 ;
    wire \line_buffer.n460 ;
    wire \line_buffer.n3635 ;
    wire \line_buffer.n566 ;
    wire \line_buffer.n558 ;
    wire \line_buffer.n557 ;
    wire \line_buffer.n565 ;
    wire \line_buffer.n3632 ;
    wire \line_buffer.n3572 ;
    wire \line_buffer.n3602_cascade_ ;
    wire \line_buffer.n3570 ;
    wire \line_buffer.n472 ;
    wire \line_buffer.n464 ;
    wire \line_buffer.n3656 ;
    wire \line_buffer.n599 ;
    wire \line_buffer.n591 ;
    wire \line_buffer.n3626 ;
    wire TX_DATA_2;
    wire n1819;
    wire \line_buffer.n3537 ;
    wire \line_buffer.n3536 ;
    wire \line_buffer.n3614 ;
    wire \line_buffer.n469 ;
    wire \line_buffer.n461 ;
    wire \line_buffer.n3569 ;
    wire DEBUG_c_2_c;
    wire \tvp_hs_buffer.BUFFER_0_0 ;
    wire \line_buffer.n598 ;
    wire \line_buffer.n590 ;
    wire \line_buffer.n3573 ;
    wire \line_buffer.n3659 ;
    wire \line_buffer.n564 ;
    wire \line_buffer.n556 ;
    wire \line_buffer.n467 ;
    wire \line_buffer.n459 ;
    wire \line_buffer.n3638 ;
    wire \line_buffer.n3641 ;
    wire TX_DATA_0;
    wire \line_buffer.n532 ;
    wire \line_buffer.n524 ;
    wire \line_buffer.n3647 ;
    wire TX_DATA_5;
    wire n1816;
    wire \line_buffer.n537 ;
    wire \line_buffer.n529 ;
    wire \line_buffer.n3599 ;
    wire \line_buffer.n597 ;
    wire \line_buffer.n589 ;
    wire \line_buffer.n3650 ;
    wire \line_buffer.n570 ;
    wire \line_buffer.n562 ;
    wire \line_buffer.n3543 ;
    wire TX_ADDR_13;
    wire \line_buffer.n3608_cascade_ ;
    wire \line_buffer.n3576 ;
    wire TX_DATA_6;
    wire n1815;
    wire ADV_CLK_c;
    wire \transmit_module.n2388 ;
    wire \line_buffer.n596 ;
    wire \line_buffer.n588 ;
    wire \line_buffer.n3644 ;
    wire \line_buffer.n473 ;
    wire \line_buffer.n465 ;
    wire \line_buffer.n3575 ;
    wire \tvp_video_buffer.BUFFER_1_9 ;
    wire RX_DATA_5;
    wire \line_buffer.n601 ;
    wire TX_ADDR_12;
    wire \line_buffer.n593 ;
    wire \line_buffer.n3596 ;
    wire DEBUG_c_7_c;
    wire \tvp_video_buffer.BUFFER_0_7 ;
    wire \tvp_video_buffer.BUFFER_1_7 ;
    wire TX_ADDR_11;
    wire \line_buffer.n538 ;
    wire \line_buffer.n530 ;
    wire \line_buffer.n3542 ;
    wire CONSTANT_ONE_NET;
    wire TVP_VIDEO_c_9;
    wire \tvp_video_buffer.BUFFER_0_9 ;
    wire DEBUG_c_3_c;
    wire _gnd_net_;

    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \tx_pll.TX_PLL_inst .TEST_MODE=1'b0;
    defparam \tx_pll.TX_PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \tx_pll.TX_PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \tx_pll.TX_PLL_inst .FILTER_RANGE=3'b010;
    defparam \tx_pll.TX_PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \tx_pll.TX_PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \tx_pll.TX_PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \tx_pll.TX_PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \tx_pll.TX_PLL_inst .DIVR=4'b0000;
    defparam \tx_pll.TX_PLL_inst .DIVQ=3'b100;
    defparam \tx_pll.TX_PLL_inst .DIVF=7'b0100110;
    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \tx_pll.TX_PLL_inst  (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(ADV_CLK_c),
            .REFERENCECLK(N__16120),
            .RESETB(N__24513),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .PLLOUTGLOBAL());
    defparam \line_buffer.mem2_physical .WRITE_MODE=3;
    defparam \line_buffer.mem2_physical .READ_MODE=3;
    defparam \line_buffer.mem2_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem2_physical  (
            .RDATA({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,\line_buffer.n474 ,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,\line_buffer.n473 ,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .RADDR({N__13726,N__12214,N__10075,N__11095,N__11380,N__11947,N__11635,N__19339,N__20383,N__8833,N__13969}),
            .WADDR({N__17671,N__16225,N__15880,N__16516,N__16777,N__17032,N__17293,N__17902,N__15340,N__15592,N__18151}),
            .MASK({dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37}),
            .WDATA({dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,N__18580,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,N__19135,dangling_wire_49,dangling_wire_50,dangling_wire_51}),
            .RCLKE(),
            .RCLK(N__23413),
            .RE(N__24378),
            .WCLKE(),
            .WCLK(N__24162),
            .WE(N__13076));
    defparam \line_buffer.mem14_physical .WRITE_MODE=3;
    defparam \line_buffer.mem14_physical .READ_MODE=3;
    defparam \line_buffer.mem14_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem14_physical  (
            .RDATA({dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,\line_buffer.n561 ,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,\line_buffer.n560 ,dangling_wire_63,dangling_wire_64,dangling_wire_65}),
            .RADDR({N__13798,N__12286,N__10147,N__11167,N__11452,N__12019,N__11707,N__19411,N__20455,N__8905,N__14041}),
            .WADDR({N__17743,N__16297,N__15952,N__16588,N__16849,N__17104,N__17365,N__17974,N__15412,N__15664,N__18223}),
            .MASK({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .WDATA({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,N__22506,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,N__19002,dangling_wire_93,dangling_wire_94,dangling_wire_95}),
            .RCLKE(),
            .RCLK(N__23510),
            .RE(N__24363),
            .WCLKE(),
            .WCLK(N__24142),
            .WE(N__12890));
    defparam \line_buffer.mem5_physical .WRITE_MODE=3;
    defparam \line_buffer.mem5_physical .READ_MODE=3;
    defparam \line_buffer.mem5_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem5_physical  (
            .RDATA({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,\line_buffer.n571 ,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\line_buffer.n570 ,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .RADDR({N__13747,N__12223,N__10090,N__11116,N__11371,N__11968,N__11650,N__19348,N__20398,N__8836,N__13984}),
            .WADDR({N__17674,N__16222,N__15889,N__16525,N__16786,N__17047,N__17308,N__17911,N__15349,N__15601,N__18148}),
            .MASK({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .WDATA({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,N__18591,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,N__19146,dangling_wire_137,dangling_wire_138,dangling_wire_139}),
            .RCLKE(),
            .RCLK(N__22912),
            .RE(N__24409),
            .WCLKE(),
            .WCLK(N__24160),
            .WE(N__14753));
    defparam \line_buffer.mem11_physical .WRITE_MODE=3;
    defparam \line_buffer.mem11_physical .READ_MODE=3;
    defparam \line_buffer.mem11_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem11_physical  (
            .RDATA({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,\line_buffer.n529 ,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,\line_buffer.n528 ,dangling_wire_151,dangling_wire_152,dangling_wire_153}),
            .RADDR({N__13834,N__12322,N__10183,N__11203,N__11488,N__12055,N__11743,N__19447,N__20491,N__8941,N__14077}),
            .WADDR({N__17779,N__16333,N__15988,N__16624,N__16885,N__17140,N__17401,N__18010,N__15448,N__15700,N__18259}),
            .MASK({dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169}),
            .WDATA({dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,N__22518,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,N__19034,dangling_wire_181,dangling_wire_182,dangling_wire_183}),
            .RCLKE(),
            .RCLK(N__23688),
            .RE(N__24454),
            .WCLKE(),
            .WCLK(N__24130),
            .WE(N__13024));
    defparam \line_buffer.mem21_physical .WRITE_MODE=3;
    defparam \line_buffer.mem21_physical .READ_MODE=3;
    defparam \line_buffer.mem21_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem21_physical  (
            .RDATA({dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,\line_buffer.n591 ,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,\line_buffer.n590 ,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .RADDR({N__13702,N__12190,N__10051,N__11071,N__11356,N__11923,N__11611,N__19315,N__20359,N__8809,N__13945}),
            .WADDR({N__17647,N__16201,N__15856,N__16492,N__16753,N__17008,N__17269,N__17878,N__15316,N__15568,N__18127}),
            .MASK({dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213}),
            .WDATA({dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,N__9068,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,N__10513,dangling_wire_225,dangling_wire_226,dangling_wire_227}),
            .RCLKE(),
            .RCLK(N__23249),
            .RE(N__24425),
            .WCLKE(),
            .WCLK(N__24166),
            .WE(N__13414));
    defparam \line_buffer.mem12_physical .WRITE_MODE=3;
    defparam \line_buffer.mem12_physical .READ_MODE=3;
    defparam \line_buffer.mem12_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem12_physical  (
            .RDATA({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,\line_buffer.n527 ,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,\line_buffer.n526 ,dangling_wire_239,dangling_wire_240,dangling_wire_241}),
            .RADDR({N__13822,N__12310,N__10171,N__11191,N__11476,N__12043,N__11731,N__19435,N__20479,N__8929,N__14065}),
            .WADDR({N__17767,N__16321,N__15976,N__16612,N__16873,N__17128,N__17389,N__17998,N__15436,N__15688,N__18247}),
            .MASK({dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .WDATA({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,N__9074,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,N__10475,dangling_wire_269,dangling_wire_270,dangling_wire_271}),
            .RCLKE(),
            .RCLK(N__23621),
            .RE(N__24412),
            .WCLKE(),
            .WCLK(N__24136),
            .WE(N__13017));
    defparam \line_buffer.mem24_physical .WRITE_MODE=3;
    defparam \line_buffer.mem24_physical .READ_MODE=3;
    defparam \line_buffer.mem24_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem24_physical  (
            .RDATA({dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,\line_buffer.n535 ,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,\line_buffer.n534 ,dangling_wire_283,dangling_wire_284,dangling_wire_285}),
            .RADDR({N__13867,N__12343,N__10210,N__11236,N__11491,N__12088,N__11770,N__19468,N__20518,N__8956,N__14104}),
            .WADDR({N__17794,N__16342,N__16009,N__16645,N__16906,N__17167,N__17428,N__18031,N__15469,N__15721,N__18268}),
            .MASK({dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301}),
            .WDATA({dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,N__9057,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,N__10489,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .RCLKE(),
            .RCLK(N__23734),
            .RE(N__24523),
            .WCLKE(),
            .WCLK(N__24117),
            .WE(N__12639));
    defparam \line_buffer.mem1_physical .WRITE_MODE=3;
    defparam \line_buffer.mem1_physical .READ_MODE=3;
    defparam \line_buffer.mem1_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem1_physical  (
            .RDATA({dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,\line_buffer.n563 ,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,\line_buffer.n562 ,dangling_wire_327,dangling_wire_328,dangling_wire_329}),
            .RADDR({N__13858,N__12346,N__10207,N__11227,N__11507,N__12079,N__11767,N__19471,N__20515,N__8965,N__14101}),
            .WADDR({N__17803,N__16355,N__16012,N__16648,N__16909,N__17164,N__17425,N__18034,N__15472,N__15724,N__18281}),
            .MASK({dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345}),
            .WDATA({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,N__18557,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,N__19119,dangling_wire_357,dangling_wire_358,dangling_wire_359}),
            .RCLKE(),
            .RCLK(N__23722),
            .RE(N__24488),
            .WCLKE(),
            .WCLK(N__24113),
            .WE(N__12902));
    defparam \line_buffer.mem15_physical .WRITE_MODE=3;
    defparam \line_buffer.mem15_physical .READ_MODE=3;
    defparam \line_buffer.mem15_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem15_physical  (
            .RDATA({dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,\line_buffer.n559 ,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,\line_buffer.n558 ,dangling_wire_371,dangling_wire_372,dangling_wire_373}),
            .RADDR({N__13786,N__12274,N__10135,N__11155,N__11440,N__12007,N__11695,N__19399,N__20443,N__8893,N__14029}),
            .WADDR({N__17731,N__16285,N__15940,N__16576,N__16837,N__17092,N__17353,N__17962,N__15400,N__15652,N__18211}),
            .MASK({dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389}),
            .WDATA({dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,N__9069,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,N__10476,dangling_wire_401,dangling_wire_402,dangling_wire_403}),
            .RCLKE(),
            .RCLK(N__23509),
            .RE(N__24342),
            .WCLKE(),
            .WCLK(N__24144),
            .WE(N__12900));
    defparam \line_buffer.mem27_physical .WRITE_MODE=3;
    defparam \line_buffer.mem27_physical .READ_MODE=3;
    defparam \line_buffer.mem27_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem27_physical  (
            .RDATA({dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,\line_buffer.n567 ,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,\line_buffer.n566 ,dangling_wire_415,dangling_wire_416,dangling_wire_417}),
            .RADDR({N__13831,N__12307,N__10174,N__11200,N__11455,N__12052,N__11734,N__19432,N__20482,N__8920,N__14068}),
            .WADDR({N__17758,N__16306,N__15973,N__16609,N__16870,N__17131,N__17392,N__17995,N__15433,N__15685,N__18232}),
            .MASK({dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .WDATA({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,N__9038,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,N__10482,dangling_wire_445,dangling_wire_446,dangling_wire_447}),
            .RCLKE(),
            .RCLK(N__23696),
            .RE(N__24496),
            .WCLKE(),
            .WCLK(N__24137),
            .WE(N__14748));
    defparam \line_buffer.mem4_physical .WRITE_MODE=3;
    defparam \line_buffer.mem4_physical .READ_MODE=3;
    defparam \line_buffer.mem4_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem4_physical  (
            .RDATA({dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,\line_buffer.n539 ,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,\line_buffer.n538 ,dangling_wire_459,dangling_wire_460,dangling_wire_461}),
            .RADDR({N__13759,N__12235,N__10102,N__11128,N__11383,N__11980,N__11662,N__19360,N__20410,N__8848,N__13996}),
            .WADDR({N__17686,N__16234,N__15901,N__16537,N__16798,N__17059,N__17320,N__17923,N__15361,N__15613,N__18160}),
            .MASK({dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477}),
            .WDATA({dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,N__18581,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,N__19136,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .RCLKE(),
            .RCLK(N__23403),
            .RE(N__24468),
            .WCLKE(),
            .WCLK(N__24158),
            .WE(N__12640));
    defparam \line_buffer.mem16_physical .WRITE_MODE=3;
    defparam \line_buffer.mem16_physical .READ_MODE=3;
    defparam \line_buffer.mem16_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem16_physical  (
            .RDATA({dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,\line_buffer.n557 ,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,\line_buffer.n556 ,dangling_wire_503,dangling_wire_504,dangling_wire_505}),
            .RADDR({N__13774,N__12262,N__10123,N__11143,N__11428,N__11995,N__11683,N__19387,N__20431,N__8881,N__14017}),
            .WADDR({N__17719,N__16273,N__15928,N__16564,N__16825,N__17080,N__17341,N__17950,N__15388,N__15640,N__18199}),
            .MASK({dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521}),
            .WDATA({dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,N__10601,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,N__10717,dangling_wire_533,dangling_wire_534,dangling_wire_535}),
            .RCLKE(),
            .RCLK(N__23358),
            .RE(N__24322),
            .WCLKE(),
            .WCLK(N__24147),
            .WE(N__12901));
    defparam \line_buffer.mem30_physical .WRITE_MODE=3;
    defparam \line_buffer.mem30_physical .READ_MODE=3;
    defparam \line_buffer.mem30_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem30_physical  (
            .RDATA({dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,\line_buffer.n599 ,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,\line_buffer.n598 ,dangling_wire_547,dangling_wire_548,dangling_wire_549}),
            .RADDR({N__13783,N__12259,N__10126,N__11152,N__11407,N__12004,N__11686,N__19384,N__20434,N__8872,N__14020}),
            .WADDR({N__17710,N__16258,N__15925,N__16561,N__16822,N__17083,N__17344,N__17947,N__15385,N__15637,N__18184}),
            .MASK({dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565}),
            .WDATA({dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,N__9001,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,N__10496,dangling_wire_577,dangling_wire_578,dangling_wire_579}),
            .RCLKE(),
            .RCLK(N__23527),
            .RE(N__24435),
            .WCLKE(),
            .WCLK(N__24152),
            .WE(N__15024));
    defparam \line_buffer.mem7_physical .WRITE_MODE=3;
    defparam \line_buffer.mem7_physical .READ_MODE=3;
    defparam \line_buffer.mem7_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem7_physical  (
            .RDATA({dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,\line_buffer.n466 ,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,\line_buffer.n465 ,dangling_wire_591,dangling_wire_592,dangling_wire_593}),
            .RADDR({N__13723,N__12199,N__10066,N__11092,N__11347,N__11944,N__11626,N__19324,N__20374,N__8812,N__13960}),
            .WADDR({N__17650,N__16198,N__15865,N__16501,N__16762,N__17023,N__17284,N__17887,N__15325,N__15577,N__18124}),
            .MASK({dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609}),
            .WDATA({dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,N__18596,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,N__19148,dangling_wire_621,dangling_wire_622,dangling_wire_623}),
            .RCLKE(),
            .RCLK(N__23298),
            .RE(N__24521),
            .WCLKE(),
            .WCLK(N__24165),
            .WE(N__14987));
    defparam \line_buffer.mem20_physical .WRITE_MODE=3;
    defparam \line_buffer.mem20_physical .READ_MODE=3;
    defparam \line_buffer.mem20_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem20_physical  (
            .RDATA({dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,\line_buffer.n593 ,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,\line_buffer.n592 ,dangling_wire_635,dangling_wire_636,dangling_wire_637}),
            .RADDR({N__13714,N__12202,N__10063,N__11083,N__11368,N__11935,N__11623,N__19327,N__20371,N__8821,N__13957}),
            .WADDR({N__17659,N__16213,N__15868,N__16504,N__16765,N__17020,N__17281,N__17890,N__15328,N__15580,N__18139}),
            .MASK({dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653}),
            .WDATA({dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,N__22517,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,N__19043,dangling_wire_665,dangling_wire_666,dangling_wire_667}),
            .RCLKE(),
            .RCLK(N__23552),
            .RE(N__24424),
            .WCLKE(),
            .WCLK(N__24164),
            .WE(N__13413));
    defparam \line_buffer.mem13_physical .WRITE_MODE=3;
    defparam \line_buffer.mem13_physical .READ_MODE=3;
    defparam \line_buffer.mem13_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem13_physical  (
            .RDATA({dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,\line_buffer.n525 ,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,\line_buffer.n524 ,dangling_wire_679,dangling_wire_680,dangling_wire_681}),
            .RADDR({N__13810,N__12298,N__10159,N__11179,N__11464,N__12031,N__11719,N__19423,N__20467,N__8917,N__14053}),
            .WADDR({N__17755,N__16309,N__15964,N__16600,N__16861,N__17116,N__17377,N__17986,N__15424,N__15676,N__18235}),
            .MASK({dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697}),
            .WDATA({dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,N__10600,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,N__10716,dangling_wire_709,dangling_wire_710,dangling_wire_711}),
            .RCLKE(),
            .RCLK(N__23620),
            .RE(N__24411),
            .WCLKE(),
            .WCLK(N__24138),
            .WE(N__13016));
    defparam \line_buffer.mem19_physical .WRITE_MODE=3;
    defparam \line_buffer.mem19_physical .READ_MODE=3;
    defparam \line_buffer.mem19_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem19_physical  (
            .RDATA({dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,\line_buffer.n468 ,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,\line_buffer.n467 ,dangling_wire_723,dangling_wire_724,dangling_wire_725}),
            .RADDR({N__13738,N__12226,N__10087,N__11107,N__11392,N__11959,N__11647,N__19351,N__20395,N__8845,N__13981}),
            .WADDR({N__17683,N__16237,N__15892,N__16528,N__16789,N__17044,N__17305,N__17914,N__15352,N__15604,N__18163}),
            .MASK({dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741}),
            .WDATA({dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,N__10602,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,N__10728,dangling_wire_753,dangling_wire_754,dangling_wire_755}),
            .RCLKE(),
            .RCLK(N__23023),
            .RE(N__24377),
            .WCLKE(),
            .WCLK(N__24159),
            .WE(N__13072));
    defparam \line_buffer.mem23_physical .WRITE_MODE=3;
    defparam \line_buffer.mem23_physical .READ_MODE=3;
    defparam \line_buffer.mem23_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem23_physical  (
            .RDATA({dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,\line_buffer.n537 ,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,\line_buffer.n536 ,dangling_wire_767,dangling_wire_768,dangling_wire_769}),
            .RADDR({N__13874,N__12355,N__10220,N__11243,N__11503,N__12095,N__11780,N__19480,N__20528,N__8968,N__14114}),
            .WADDR({N__17806,N__16354,N__16021,N__16657,N__16918,N__17177,N__17438,N__18043,N__15481,N__15733,N__18280}),
            .MASK({dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785}),
            .WDATA({dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,N__22523,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,N__19006,dangling_wire_797,dangling_wire_798,dangling_wire_799}),
            .RCLKE(),
            .RCLK(N__23735),
            .RE(N__24524),
            .WCLKE(),
            .WCLK(N__24109),
            .WE(N__12641));
    defparam \line_buffer.mem0_physical .WRITE_MODE=3;
    defparam \line_buffer.mem0_physical .READ_MODE=3;
    defparam \line_buffer.mem0_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem0_physical  (
            .RDATA({dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,\line_buffer.n531 ,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,\line_buffer.n530 ,dangling_wire_811,dangling_wire_812,dangling_wire_813}),
            .RADDR({N__13870,N__12356,N__10219,N__11239,N__11513,N__12091,N__11779,N__19481,N__20527,N__8972,N__14113}),
            .WADDR({N__17810,N__16361,N__16022,N__16658,N__16919,N__17176,N__17437,N__18044,N__15482,N__15734,N__18287}),
            .MASK({dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829}),
            .WDATA({dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,N__18579,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,N__19120,dangling_wire_841,dangling_wire_842,dangling_wire_843}),
            .RCLKE(),
            .RCLK(N__23723),
            .RE(N__24489),
            .WCLKE(),
            .WCLK(N__24104),
            .WE(N__13028));
    defparam \line_buffer.mem26_physical .WRITE_MODE=3;
    defparam \line_buffer.mem26_physical .READ_MODE=3;
    defparam \line_buffer.mem26_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem26_physical  (
            .RDATA({dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,\line_buffer.n569 ,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,\line_buffer.n568 ,dangling_wire_855,dangling_wire_856,dangling_wire_857}),
            .RADDR({N__13843,N__12319,N__10186,N__11212,N__11467,N__12064,N__11746,N__19444,N__20494,N__8932,N__14080}),
            .WADDR({N__17770,N__16318,N__15985,N__16621,N__16882,N__17143,N__17404,N__18007,N__15445,N__15697,N__18244}),
            .MASK({dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873}),
            .WDATA({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,N__22513,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,N__19021,dangling_wire_885,dangling_wire_886,dangling_wire_887}),
            .RCLKE(),
            .RCLK(N__23724),
            .RE(N__24408),
            .WCLKE(),
            .WCLK(N__24134),
            .WE(N__14749));
    defparam \line_buffer.mem3_physical .WRITE_MODE=3;
    defparam \line_buffer.mem3_physical .READ_MODE=3;
    defparam \line_buffer.mem3_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem3_physical  (
            .RDATA({dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,\line_buffer.n595 ,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,\line_buffer.n594 ,dangling_wire_899,dangling_wire_900,dangling_wire_901}),
            .RADDR({N__13795,N__12271,N__10138,N__11164,N__11419,N__12016,N__11698,N__19396,N__20446,N__8884,N__14032}),
            .WADDR({N__17722,N__16270,N__15937,N__16573,N__16834,N__17095,N__17356,N__17959,N__15397,N__15649,N__18196}),
            .MASK({dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917}),
            .WDATA({dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,N__18556,dangling_wire_922,dangling_wire_923,dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,dangling_wire_928,N__19111,dangling_wire_929,dangling_wire_930,dangling_wire_931}),
            .RCLKE(),
            .RCLK(N__23478),
            .RE(N__24469),
            .WCLKE(),
            .WCLK(N__24145),
            .WE(N__13403));
    defparam \line_buffer.mem17_physical .WRITE_MODE=3;
    defparam \line_buffer.mem17_physical .READ_MODE=3;
    defparam \line_buffer.mem17_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem17_physical  (
            .RDATA({dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,\line_buffer.n472 ,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,\line_buffer.n471 ,dangling_wire_943,dangling_wire_944,dangling_wire_945}),
            .RADDR({N__13762,N__12250,N__10111,N__11131,N__11416,N__11983,N__11671,N__19375,N__20419,N__8869,N__14005}),
            .WADDR({N__17707,N__16261,N__15916,N__16552,N__16813,N__17068,N__17329,N__17938,N__15376,N__15628,N__18187}),
            .MASK({dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961}),
            .WDATA({dangling_wire_962,dangling_wire_963,dangling_wire_964,dangling_wire_965,N__22483,dangling_wire_966,dangling_wire_967,dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,dangling_wire_972,N__19036,dangling_wire_973,dangling_wire_974,dangling_wire_975}),
            .RCLKE(),
            .RCLK(N__23357),
            .RE(N__24269),
            .WCLKE(),
            .WCLK(N__24153),
            .WE(N__13061));
    defparam \line_buffer.mem31_physical .WRITE_MODE=3;
    defparam \line_buffer.mem31_physical .READ_MODE=3;
    defparam \line_buffer.mem31_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem31_physical  (
            .RDATA({dangling_wire_976,dangling_wire_977,dangling_wire_978,dangling_wire_979,\line_buffer.n597 ,dangling_wire_980,dangling_wire_981,dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,\line_buffer.n596 ,dangling_wire_987,dangling_wire_988,dangling_wire_989}),
            .RADDR({N__13771,N__12247,N__10114,N__11140,N__11395,N__11992,N__11674,N__19372,N__20422,N__8860,N__14008}),
            .WADDR({N__17698,N__16246,N__15913,N__16549,N__16810,N__17071,N__17332,N__17935,N__15373,N__15625,N__18172}),
            .MASK({dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997,dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005}),
            .WDATA({dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,dangling_wire_1009,N__10610,dangling_wire_1010,dangling_wire_1011,dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,dangling_wire_1016,N__10736,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019}),
            .RCLKE(),
            .RCLK(N__23331),
            .RE(N__24343),
            .WCLKE(),
            .WCLK(N__24154),
            .WE(N__15031));
    defparam \line_buffer.mem9_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .WRITE_MODE=3;
    defparam \line_buffer.mem9_physical .READ_MODE=3;
    defparam \line_buffer.mem9_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem9_physical  (
            .RDATA({dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,dangling_wire_1023,\line_buffer.n462 ,dangling_wire_1024,dangling_wire_1025,dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,\line_buffer.n461 ,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033}),
            .RADDR({N__13699,N__12175,N__10042,N__11068,N__11323,N__11920,N__11602,N__19300,N__20350,N__8788,N__13936}),
            .WADDR({N__17626,N__16174,N__15841,N__16477,N__16738,N__16999,N__17260,N__17863,N__15301,N__15553,N__18100}),
            .MASK({dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041,dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049}),
            .WDATA({dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,dangling_wire_1053,N__9058,dangling_wire_1054,dangling_wire_1055,dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,dangling_wire_1060,N__10517,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063}),
            .RCLKE(),
            .RCLK(N__22955),
            .RE(N__24407),
            .WCLKE(),
            .WCLK(N__24169),
            .WE(N__14993));
    defparam \line_buffer.mem29_physical .WRITE_MODE=3;
    defparam \line_buffer.mem29_physical .READ_MODE=3;
    defparam \line_buffer.mem29_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem29_physical  (
            .RDATA({dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,dangling_wire_1067,\line_buffer.n601 ,dangling_wire_1068,dangling_wire_1069,dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,\line_buffer.n600 ,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077}),
            .RADDR({N__13807,N__12283,N__10150,N__11176,N__11431,N__12028,N__11710,N__19408,N__20458,N__8896,N__14044}),
            .WADDR({N__17734,N__16282,N__15949,N__16585,N__16846,N__17107,N__17368,N__17971,N__15409,N__15661,N__18208}),
            .MASK({dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085,dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093}),
            .WDATA({dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,dangling_wire_1097,N__22519,dangling_wire_1098,dangling_wire_1099,dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,dangling_wire_1104,N__19001,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107}),
            .RCLKE(),
            .RCLK(N__23636),
            .RE(N__24470),
            .WCLKE(),
            .WCLK(N__24143),
            .WE(N__15015));
    defparam \line_buffer.mem6_physical .WRITE_MODE=3;
    defparam \line_buffer.mem6_physical .READ_MODE=3;
    defparam \line_buffer.mem6_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem6_physical  (
            .RDATA({dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,dangling_wire_1111,\line_buffer.n603 ,dangling_wire_1112,dangling_wire_1113,dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,\line_buffer.n602 ,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121}),
            .RADDR({N__13735,N__12211,N__10078,N__11104,N__11359,N__11956,N__11638,N__19336,N__20386,N__8824,N__13972}),
            .WADDR({N__17662,N__16210,N__15877,N__16513,N__16774,N__17035,N__17296,N__17899,N__15337,N__15589,N__18136}),
            .MASK({dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129,dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137}),
            .WDATA({dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,dangling_wire_1141,N__18592,dangling_wire_1142,dangling_wire_1143,dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,dangling_wire_1148,N__19147,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151}),
            .RCLKE(),
            .RCLK(N__23466),
            .RE(N__24505),
            .WCLKE(),
            .WCLK(N__24163),
            .WE(N__15035));
    defparam \line_buffer.mem10_physical .WRITE_MODE=3;
    defparam \line_buffer.mem10_physical .READ_MODE=3;
    defparam \line_buffer.mem10_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem10_physical  (
            .RDATA({dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,dangling_wire_1155,\line_buffer.n460 ,dangling_wire_1156,dangling_wire_1157,dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,\line_buffer.n459 ,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165}),
            .RADDR({N__13846,N__12334,N__10195,N__11215,N__11500,N__12067,N__11755,N__19459,N__20503,N__8953,N__14089}),
            .WADDR({N__17791,N__16345,N__16000,N__16636,N__16897,N__17152,N__17413,N__18022,N__15460,N__15712,N__18271}),
            .MASK({dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173,dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181}),
            .WDATA({dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,dangling_wire_1185,N__10599,dangling_wire_1186,dangling_wire_1187,dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,dangling_wire_1192,N__10715,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195}),
            .RCLKE(),
            .RCLK(N__23689),
            .RE(N__24455),
            .WCLKE(),
            .WCLK(N__24120),
            .WE(N__14992));
    defparam \line_buffer.mem22_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .WRITE_MODE=3;
    defparam \line_buffer.mem22_physical .READ_MODE=3;
    defparam \line_buffer.mem22_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem22_physical  (
            .RDATA({dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,dangling_wire_1199,\line_buffer.n589 ,dangling_wire_1200,dangling_wire_1201,dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,\line_buffer.n588 ,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209}),
            .RADDR({N__13690,N__12178,N__10039,N__11059,N__11344,N__11911,N__11599,N__19303,N__20347,N__8797,N__13933}),
            .WADDR({N__17635,N__16189,N__15844,N__16480,N__16741,N__16996,N__17257,N__17866,N__15304,N__15556,N__18115}),
            .MASK({dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217,dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225}),
            .WDATA({dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,dangling_wire_1229,N__10609,dangling_wire_1230,dangling_wire_1231,dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,dangling_wire_1236,N__10735,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239}),
            .RCLKE(),
            .RCLK(N__23253),
            .RE(N__24462),
            .WCLKE(),
            .WCLK(N__24168),
            .WE(N__13418));
    defparam \line_buffer.mem25_physical .WRITE_MODE=3;
    defparam \line_buffer.mem25_physical .READ_MODE=3;
    defparam \line_buffer.mem25_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem25_physical  (
            .RDATA({dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,dangling_wire_1243,\line_buffer.n533 ,dangling_wire_1244,dangling_wire_1245,dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,\line_buffer.n532 ,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253}),
            .RADDR({N__13855,N__12331,N__10198,N__11224,N__11479,N__12076,N__11758,N__19456,N__20506,N__8944,N__14092}),
            .WADDR({N__17782,N__16330,N__15997,N__16633,N__16894,N__17155,N__17416,N__18019,N__15457,N__15709,N__18256}),
            .MASK({dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261,dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269}),
            .WDATA({dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,dangling_wire_1273,N__10594,dangling_wire_1274,dangling_wire_1275,dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,dangling_wire_1280,N__10708,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283}),
            .RCLKE(),
            .RCLK(N__23730),
            .RE(N__24514),
            .WCLKE(),
            .WCLK(N__24126),
            .WE(N__12626));
    defparam \line_buffer.mem8_physical .WRITE_MODE=3;
    defparam \line_buffer.mem8_physical .READ_MODE=3;
    defparam \line_buffer.mem8_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem8_physical  (
            .RDATA({dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,dangling_wire_1287,\line_buffer.n464 ,dangling_wire_1288,dangling_wire_1289,dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,\line_buffer.n463 ,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297}),
            .RADDR({N__13711,N__12187,N__10054,N__11080,N__11335,N__11932,N__11614,N__19312,N__20362,N__8800,N__13948}),
            .WADDR({N__17638,N__16186,N__15853,N__16489,N__16750,N__17011,N__17272,N__17875,N__15313,N__15565,N__18112}),
            .MASK({dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305,dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313}),
            .WDATA({dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,dangling_wire_1317,N__22496,dangling_wire_1318,dangling_wire_1319,dangling_wire_1320,dangling_wire_1321,dangling_wire_1322,dangling_wire_1323,dangling_wire_1324,N__19035,dangling_wire_1325,dangling_wire_1326,dangling_wire_1327}),
            .RCLKE(),
            .RCLK(N__23083),
            .RE(N__24522),
            .WCLKE(),
            .WCLK(N__24167),
            .WE(N__14988));
    defparam \line_buffer.mem28_physical .WRITE_MODE=3;
    defparam \line_buffer.mem28_physical .READ_MODE=3;
    defparam \line_buffer.mem28_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem28_physical  (
            .RDATA({dangling_wire_1328,dangling_wire_1329,dangling_wire_1330,dangling_wire_1331,\line_buffer.n565 ,dangling_wire_1332,dangling_wire_1333,dangling_wire_1334,dangling_wire_1335,dangling_wire_1336,dangling_wire_1337,dangling_wire_1338,\line_buffer.n564 ,dangling_wire_1339,dangling_wire_1340,dangling_wire_1341}),
            .RADDR({N__13819,N__12295,N__10162,N__11188,N__11443,N__12040,N__11722,N__19420,N__20470,N__8908,N__14056}),
            .WADDR({N__17746,N__16294,N__15961,N__16597,N__16858,N__17119,N__17380,N__17983,N__15421,N__15673,N__18220}),
            .MASK({dangling_wire_1342,dangling_wire_1343,dangling_wire_1344,dangling_wire_1345,dangling_wire_1346,dangling_wire_1347,dangling_wire_1348,dangling_wire_1349,dangling_wire_1350,dangling_wire_1351,dangling_wire_1352,dangling_wire_1353,dangling_wire_1354,dangling_wire_1355,dangling_wire_1356,dangling_wire_1357}),
            .WDATA({dangling_wire_1358,dangling_wire_1359,dangling_wire_1360,dangling_wire_1361,N__10595,dangling_wire_1362,dangling_wire_1363,dangling_wire_1364,dangling_wire_1365,dangling_wire_1366,dangling_wire_1367,dangling_wire_1368,N__10724,dangling_wire_1369,dangling_wire_1370,dangling_wire_1371}),
            .RCLKE(),
            .RCLK(N__23037),
            .RE(N__24410),
            .WCLKE(),
            .WCLK(N__24140),
            .WE(N__14741));
    defparam \line_buffer.mem18_physical .WRITE_MODE=3;
    defparam \line_buffer.mem18_physical .READ_MODE=3;
    defparam \line_buffer.mem18_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem18_physical  (
            .RDATA({dangling_wire_1372,dangling_wire_1373,dangling_wire_1374,dangling_wire_1375,\line_buffer.n470 ,dangling_wire_1376,dangling_wire_1377,dangling_wire_1378,dangling_wire_1379,dangling_wire_1380,dangling_wire_1381,dangling_wire_1382,\line_buffer.n469 ,dangling_wire_1383,dangling_wire_1384,dangling_wire_1385}),
            .RADDR({N__13750,N__12238,N__10099,N__11119,N__11404,N__11971,N__11659,N__19363,N__20407,N__8857,N__13993}),
            .WADDR({N__17695,N__16249,N__15904,N__16540,N__16801,N__17056,N__17317,N__17926,N__15364,N__15616,N__18175}),
            .MASK({dangling_wire_1386,dangling_wire_1387,dangling_wire_1388,dangling_wire_1389,dangling_wire_1390,dangling_wire_1391,dangling_wire_1392,dangling_wire_1393,dangling_wire_1394,dangling_wire_1395,dangling_wire_1396,dangling_wire_1397,dangling_wire_1398,dangling_wire_1399,dangling_wire_1400,dangling_wire_1401}),
            .WDATA({dangling_wire_1402,dangling_wire_1403,dangling_wire_1404,dangling_wire_1405,N__9070,dangling_wire_1406,dangling_wire_1407,dangling_wire_1408,dangling_wire_1409,dangling_wire_1410,dangling_wire_1411,dangling_wire_1412,N__10500,dangling_wire_1413,dangling_wire_1414,dangling_wire_1415}),
            .RCLKE(),
            .RCLK(N__23184),
            .RE(N__24323),
            .WCLKE(),
            .WCLK(N__24156),
            .WE(N__13071));
    PRE_IO_GBUF DEBUG_c_3_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__25263),
            .GLOBALBUFFEROUTPUT(DEBUG_c_3_c));
    defparam DEBUG_c_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_3_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_3_pad_iopad (
            .OE(N__25265),
            .DIN(N__25264),
            .DOUT(N__25263),
            .PACKAGEPIN(TVP_CLK));
    defparam DEBUG_c_3_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_3_pad_preio (
            .PADOEN(N__25265),
            .PADOUT(N__25264),
            .PADIN(N__25263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_CLK_pad_iopad (
            .OE(N__25254),
            .DIN(N__25253),
            .DOUT(N__25252),
            .PACKAGEPIN(ADV_CLK));
    defparam ADV_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_CLK_pad_preio (
            .PADOEN(N__25254),
            .PADOUT(N__25253),
            .PADIN(N__25252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23278),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_2_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_2_pad_iopad (
            .OE(N__25245),
            .DIN(N__25244),
            .DOUT(N__25243),
            .PACKAGEPIN(TVP_HSYNC));
    defparam DEBUG_c_2_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_2_pad_preio (
            .PADOEN(N__25245),
            .PADOUT(N__25244),
            .PADIN(N__25243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_3_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_3_iopad (
            .OE(N__25236),
            .DIN(N__25235),
            .DOUT(N__25234),
            .PACKAGEPIN(DEBUG[3]));
    defparam DEBUG_pad_3_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_3_preio (
            .PADOEN(N__25236),
            .PADOUT(N__25235),
            .PADIN(N__25234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16121),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_2_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_2_iopad (
            .OE(N__25227),
            .DIN(N__25226),
            .DOUT(N__25225),
            .PACKAGEPIN(TVP_VIDEO[2]));
    defparam TVP_VIDEO_pad_2_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_2_preio (
            .PADOEN(N__25227),
            .PADOUT(N__25226),
            .PADIN(N__25225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_5_iopad (
            .OE(N__25218),
            .DIN(N__25217),
            .DOUT(N__25216),
            .PACKAGEPIN(ADV_G[5]));
    defparam ADV_G_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_5_preio (
            .PADOEN(N__25218),
            .PADOUT(N__25217),
            .PADIN(N__25216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21994),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_3_iopad (
            .OE(N__25209),
            .DIN(N__25208),
            .DOUT(N__25207),
            .PACKAGEPIN(ADV_R[3]));
    defparam ADV_R_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_3_preio (
            .PADOEN(N__25209),
            .PADOUT(N__25208),
            .PADIN(N__25207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19263),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_0_iopad (
            .OE(N__25200),
            .DIN(N__25199),
            .DOUT(N__25198),
            .PACKAGEPIN(ADV_R[0]));
    defparam ADV_R_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_0_preio (
            .PADOEN(N__25200),
            .PADOUT(N__25199),
            .PADIN(N__25198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16084),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_2_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_2_iopad (
            .OE(N__25191),
            .DIN(N__25190),
            .DOUT(N__25189),
            .PACKAGEPIN(DEBUG[2]));
    defparam DEBUG_pad_2_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_2_preio (
            .PADOEN(N__25191),
            .PADOUT(N__25190),
            .PADIN(N__25189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21644),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_3_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_3_iopad (
            .OE(N__25182),
            .DIN(N__25181),
            .DOUT(N__25180),
            .PACKAGEPIN(TVP_VIDEO[3]));
    defparam TVP_VIDEO_pad_3_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_3_preio (
            .PADOEN(N__25182),
            .PADOUT(N__25181),
            .PADIN(N__25180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_4_iopad (
            .OE(N__25173),
            .DIN(N__25172),
            .DOUT(N__25171),
            .PACKAGEPIN(ADV_G[4]));
    defparam ADV_G_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_4_preio (
            .PADOEN(N__25173),
            .PADOUT(N__25172),
            .PADIN(N__25171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20969),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_5_iopad (
            .OE(N__25164),
            .DIN(N__25163),
            .DOUT(N__25162),
            .PACKAGEPIN(ADV_R[5]));
    defparam ADV_R_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_5_preio (
            .PADOEN(N__25164),
            .PADOUT(N__25163),
            .PADIN(N__25162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21984),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_9_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_9_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_9_iopad (
            .OE(N__25155),
            .DIN(N__25154),
            .DOUT(N__25153),
            .PACKAGEPIN(TVP_VIDEO[9]));
    defparam TVP_VIDEO_pad_9_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_9_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_9_preio (
            .PADOEN(N__25155),
            .PADOUT(N__25154),
            .PADIN(N__25153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_1_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_1_iopad (
            .OE(N__25146),
            .DIN(N__25145),
            .DOUT(N__25144),
            .PACKAGEPIN(DEBUG[1]));
    defparam DEBUG_pad_1_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_1_preio (
            .PADOEN(N__25146),
            .PADOUT(N__25145),
            .PADIN(N__25144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14426),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_6_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_6_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_6_pad_iopad (
            .OE(N__25137),
            .DIN(N__25136),
            .DOUT(N__25135),
            .PACKAGEPIN(TVP_VIDEO[6]));
    defparam DEBUG_c_6_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_6_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_6_pad_preio (
            .PADOEN(N__25137),
            .PADOUT(N__25136),
            .PADIN(N__25135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_6_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_1_iopad (
            .OE(N__25128),
            .DIN(N__25127),
            .DOUT(N__25126),
            .PACKAGEPIN(ADV_B[1]));
    defparam ADV_B_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_1_preio (
            .PADOEN(N__25128),
            .PADOUT(N__25127),
            .PADIN(N__25126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20875),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_SYNC_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_SYNC_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_SYNC_N_pad_iopad (
            .OE(N__25119),
            .DIN(N__25118),
            .DOUT(N__25117),
            .PACKAGEPIN(ADV_SYNC_N));
    defparam ADV_SYNC_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_SYNC_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_SYNC_N_pad_preio (
            .PADOEN(N__25119),
            .PADOUT(N__25118),
            .PADIN(N__25117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_6_iopad (
            .OE(N__25110),
            .DIN(N__25109),
            .DOUT(N__25108),
            .PACKAGEPIN(ADV_B[6]));
    defparam ADV_B_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_6_preio (
            .PADOEN(N__25110),
            .PADOUT(N__25109),
            .PADIN(N__25108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23791),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_6_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_6_iopad (
            .OE(N__25101),
            .DIN(N__25100),
            .DOUT(N__25099),
            .PACKAGEPIN(DEBUG[6]));
    defparam DEBUG_pad_6_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_6_preio (
            .PADOEN(N__25101),
            .PADOUT(N__25100),
            .PADIN(N__25099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14399),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_0_iopad (
            .OE(N__25092),
            .DIN(N__25091),
            .DOUT(N__25090),
            .PACKAGEPIN(ADV_G[0]));
    defparam ADV_G_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_0_preio (
            .PADOEN(N__25092),
            .PADOUT(N__25091),
            .PADIN(N__25090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16085),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_1_iopad (
            .OE(N__25083),
            .DIN(N__25082),
            .DOUT(N__25081),
            .PACKAGEPIN(ADV_R[1]));
    defparam ADV_R_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_1_preio (
            .PADOEN(N__25083),
            .PADOUT(N__25082),
            .PADIN(N__25081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20890),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_5_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_5_iopad (
            .OE(N__25074),
            .DIN(N__25073),
            .DOUT(N__25072),
            .PACKAGEPIN(DEBUG[5]));
    defparam DEBUG_pad_5_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_5_preio (
            .PADOEN(N__25074),
            .PADOUT(N__25073),
            .PADIN(N__25072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9107),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_7_iopad (
            .OE(N__25065),
            .DIN(N__25064),
            .DOUT(N__25063),
            .PACKAGEPIN(ADV_G[7]));
    defparam ADV_G_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_7_preio (
            .PADOEN(N__25065),
            .PADOUT(N__25064),
            .PADIN(N__25063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12727),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_6_iopad (
            .OE(N__25056),
            .DIN(N__25055),
            .DOUT(N__25054),
            .PACKAGEPIN(ADV_R[6]));
    defparam ADV_R_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_6_preio (
            .PADOEN(N__25056),
            .PADOUT(N__25055),
            .PADIN(N__25054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23795),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_BLANK_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_BLANK_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_BLANK_N_pad_iopad (
            .OE(N__25047),
            .DIN(N__25046),
            .DOUT(N__25045),
            .PACKAGEPIN(ADV_BLANK_N));
    defparam ADV_BLANK_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_BLANK_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_BLANK_N_pad_preio (
            .PADOEN(N__25047),
            .PADOUT(N__25046),
            .PADIN(N__25045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24512),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_0_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_0_iopad (
            .OE(N__25038),
            .DIN(N__25037),
            .DOUT(N__25036),
            .PACKAGEPIN(DEBUG[0]));
    defparam DEBUG_pad_0_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_0_preio (
            .PADOEN(N__25038),
            .PADOUT(N__25037),
            .PADIN(N__25036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18818),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_2_iopad (
            .OE(N__25029),
            .DIN(N__25028),
            .DOUT(N__25027),
            .PACKAGEPIN(ADV_B[2]));
    defparam ADV_B_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_2_preio (
            .PADOEN(N__25029),
            .PADOUT(N__25028),
            .PADIN(N__25027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21747),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_7_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_7_pad_iopad (
            .OE(N__25020),
            .DIN(N__25019),
            .DOUT(N__25018),
            .PACKAGEPIN(TVP_VIDEO[7]));
    defparam DEBUG_c_7_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_7_pad_preio (
            .PADOEN(N__25020),
            .PADOUT(N__25019),
            .PADIN(N__25018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_7_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_1_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_1_pad_iopad (
            .OE(N__25011),
            .DIN(N__25010),
            .DOUT(N__25009),
            .PACKAGEPIN(TVP_VSYNC));
    defparam DEBUG_c_1_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_1_pad_preio (
            .PADOEN(N__25011),
            .PADOUT(N__25010),
            .PADIN(N__25009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_5_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_5_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_5_pad_iopad (
            .OE(N__25002),
            .DIN(N__25001),
            .DOUT(N__25000),
            .PACKAGEPIN(TVP_VIDEO[5]));
    defparam DEBUG_c_5_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_5_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_5_pad_preio (
            .PADOEN(N__25002),
            .PADOUT(N__25001),
            .PADIN(N__25000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_5_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_7_iopad (
            .OE(N__24993),
            .DIN(N__24992),
            .DOUT(N__24991),
            .PACKAGEPIN(ADV_B[7]));
    defparam ADV_B_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_7_preio (
            .PADOEN(N__24993),
            .PADOUT(N__24992),
            .PADIN(N__24991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12726),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b1;
    IO_PAD LED_pad_iopad (
            .OE(N__24984),
            .DIN(N__24983),
            .DOUT(N__24982),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__24984),
            .PADOUT(N__24983),
            .PADIN(N__24982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17495),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_4_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_4_iopad (
            .OE(N__24975),
            .DIN(N__24974),
            .DOUT(N__24973),
            .PACKAGEPIN(TVP_VIDEO[4]));
    defparam TVP_VIDEO_pad_4_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_4_preio (
            .PADOEN(N__24975),
            .PADOUT(N__24974),
            .PADIN(N__24973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_3_iopad (
            .OE(N__24966),
            .DIN(N__24965),
            .DOUT(N__24964),
            .PACKAGEPIN(ADV_G[3]));
    defparam ADV_G_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_3_preio (
            .PADOEN(N__24966),
            .PADOUT(N__24965),
            .PADIN(N__24964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19268),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_HSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_HSYNC_pad_iopad (
            .OE(N__24957),
            .DIN(N__24956),
            .DOUT(N__24955),
            .PACKAGEPIN(ADV_HSYNC));
    defparam ADV_HSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_HSYNC_pad_preio (
            .PADOEN(N__24957),
            .PADOUT(N__24956),
            .PADIN(N__24955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10829),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_2_iopad (
            .OE(N__24948),
            .DIN(N__24947),
            .DOUT(N__24946),
            .PACKAGEPIN(ADV_R[2]));
    defparam ADV_R_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_2_preio (
            .PADOEN(N__24948),
            .PADOUT(N__24947),
            .PADIN(N__24946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21760),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_4_iopad (
            .OE(N__24939),
            .DIN(N__24938),
            .DOUT(N__24937),
            .PACKAGEPIN(ADV_B[4]));
    defparam ADV_B_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_4_preio (
            .PADOEN(N__24939),
            .PADOUT(N__24938),
            .PADIN(N__24937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20964),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_4_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_4_iopad (
            .OE(N__24930),
            .DIN(N__24929),
            .DOUT(N__24928),
            .PACKAGEPIN(DEBUG[4]));
    defparam DEBUG_pad_4_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_4_preio (
            .PADOEN(N__24930),
            .PADOUT(N__24929),
            .PADIN(N__24928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18767),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_6_iopad (
            .OE(N__24921),
            .DIN(N__24920),
            .DOUT(N__24919),
            .PACKAGEPIN(ADV_G[6]));
    defparam ADV_G_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_6_preio (
            .PADOEN(N__24921),
            .PADOUT(N__24920),
            .PADIN(N__24919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23790),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_7_iopad (
            .OE(N__24912),
            .DIN(N__24911),
            .DOUT(N__24910),
            .PACKAGEPIN(ADV_R[7]));
    defparam ADV_R_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_7_preio (
            .PADOEN(N__24912),
            .PADOUT(N__24911),
            .PADIN(N__24910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12728),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_3_iopad (
            .OE(N__24903),
            .DIN(N__24902),
            .DOUT(N__24901),
            .PACKAGEPIN(ADV_B[3]));
    defparam ADV_B_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_3_preio (
            .PADOEN(N__24903),
            .PADOUT(N__24902),
            .PADIN(N__24901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19264),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_4_iopad (
            .OE(N__24894),
            .DIN(N__24893),
            .DOUT(N__24892),
            .PACKAGEPIN(ADV_R[4]));
    defparam ADV_R_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_4_preio (
            .PADOEN(N__24894),
            .PADOUT(N__24893),
            .PADIN(N__24892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20965),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_8_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_8_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_8_iopad (
            .OE(N__24885),
            .DIN(N__24884),
            .DOUT(N__24883),
            .PACKAGEPIN(TVP_VIDEO[8]));
    defparam TVP_VIDEO_pad_8_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_8_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_8_preio (
            .PADOEN(N__24885),
            .PADOUT(N__24884),
            .PADIN(N__24883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_0_iopad (
            .OE(N__24876),
            .DIN(N__24875),
            .DOUT(N__24874),
            .PACKAGEPIN(ADV_B[0]));
    defparam ADV_B_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_0_preio (
            .PADOEN(N__24876),
            .PADOUT(N__24875),
            .PADIN(N__24874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16074),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_2_iopad (
            .OE(N__24867),
            .DIN(N__24866),
            .DOUT(N__24865),
            .PACKAGEPIN(ADV_G[2]));
    defparam ADV_G_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_2_preio (
            .PADOEN(N__24867),
            .PADOUT(N__24866),
            .PADIN(N__24865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21764),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_VSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_VSYNC_pad_iopad (
            .OE(N__24858),
            .DIN(N__24857),
            .DOUT(N__24856),
            .PACKAGEPIN(ADV_VSYNC));
    defparam ADV_VSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_VSYNC_pad_preio (
            .PADOEN(N__24858),
            .PADOUT(N__24857),
            .PADIN(N__24856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19996),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_5_iopad (
            .OE(N__24849),
            .DIN(N__24848),
            .DOUT(N__24847),
            .PACKAGEPIN(ADV_B[5]));
    defparam ADV_B_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_5_preio (
            .PADOEN(N__24849),
            .PADOUT(N__24848),
            .PADIN(N__24847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21995),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_7_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_7_iopad (
            .OE(N__24840),
            .DIN(N__24839),
            .DOUT(N__24838),
            .PACKAGEPIN(DEBUG[7]));
    defparam DEBUG_pad_7_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_7_preio (
            .PADOEN(N__24840),
            .PADOUT(N__24839),
            .PADIN(N__24838),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22169),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_1_iopad (
            .OE(N__24831),
            .DIN(N__24830),
            .DOUT(N__24829),
            .PACKAGEPIN(ADV_G[1]));
    defparam ADV_G_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_1_preio (
            .PADOEN(N__24831),
            .PADOUT(N__24830),
            .PADIN(N__24829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__6001 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__6000 (
            .O(N__24809),
            .I(\tvp_video_buffer.BUFFER_0_7 ));
    InMux I__5999 (
            .O(N__24806),
            .I(N__24803));
    LocalMux I__5998 (
            .O(N__24803),
            .I(\tvp_video_buffer.BUFFER_1_7 ));
    InMux I__5997 (
            .O(N__24800),
            .I(N__24790));
    InMux I__5996 (
            .O(N__24799),
            .I(N__24787));
    InMux I__5995 (
            .O(N__24798),
            .I(N__24781));
    InMux I__5994 (
            .O(N__24797),
            .I(N__24776));
    InMux I__5993 (
            .O(N__24796),
            .I(N__24773));
    InMux I__5992 (
            .O(N__24795),
            .I(N__24769));
    InMux I__5991 (
            .O(N__24794),
            .I(N__24766));
    InMux I__5990 (
            .O(N__24793),
            .I(N__24760));
    LocalMux I__5989 (
            .O(N__24790),
            .I(N__24757));
    LocalMux I__5988 (
            .O(N__24787),
            .I(N__24754));
    InMux I__5987 (
            .O(N__24786),
            .I(N__24749));
    InMux I__5986 (
            .O(N__24785),
            .I(N__24749));
    InMux I__5985 (
            .O(N__24784),
            .I(N__24746));
    LocalMux I__5984 (
            .O(N__24781),
            .I(N__24740));
    InMux I__5983 (
            .O(N__24780),
            .I(N__24737));
    InMux I__5982 (
            .O(N__24779),
            .I(N__24734));
    LocalMux I__5981 (
            .O(N__24776),
            .I(N__24727));
    LocalMux I__5980 (
            .O(N__24773),
            .I(N__24727));
    InMux I__5979 (
            .O(N__24772),
            .I(N__24724));
    LocalMux I__5978 (
            .O(N__24769),
            .I(N__24719));
    LocalMux I__5977 (
            .O(N__24766),
            .I(N__24719));
    InMux I__5976 (
            .O(N__24765),
            .I(N__24716));
    InMux I__5975 (
            .O(N__24764),
            .I(N__24711));
    InMux I__5974 (
            .O(N__24763),
            .I(N__24708));
    LocalMux I__5973 (
            .O(N__24760),
            .I(N__24705));
    Span4Mux_h I__5972 (
            .O(N__24757),
            .I(N__24696));
    Span4Mux_v I__5971 (
            .O(N__24754),
            .I(N__24696));
    LocalMux I__5970 (
            .O(N__24749),
            .I(N__24696));
    LocalMux I__5969 (
            .O(N__24746),
            .I(N__24696));
    InMux I__5968 (
            .O(N__24745),
            .I(N__24693));
    InMux I__5967 (
            .O(N__24744),
            .I(N__24690));
    InMux I__5966 (
            .O(N__24743),
            .I(N__24687));
    Span4Mux_v I__5965 (
            .O(N__24740),
            .I(N__24681));
    LocalMux I__5964 (
            .O(N__24737),
            .I(N__24681));
    LocalMux I__5963 (
            .O(N__24734),
            .I(N__24678));
    InMux I__5962 (
            .O(N__24733),
            .I(N__24675));
    InMux I__5961 (
            .O(N__24732),
            .I(N__24672));
    Span4Mux_v I__5960 (
            .O(N__24727),
            .I(N__24669));
    LocalMux I__5959 (
            .O(N__24724),
            .I(N__24666));
    Span4Mux_v I__5958 (
            .O(N__24719),
            .I(N__24663));
    LocalMux I__5957 (
            .O(N__24716),
            .I(N__24660));
    InMux I__5956 (
            .O(N__24715),
            .I(N__24657));
    InMux I__5955 (
            .O(N__24714),
            .I(N__24654));
    LocalMux I__5954 (
            .O(N__24711),
            .I(N__24651));
    LocalMux I__5953 (
            .O(N__24708),
            .I(N__24642));
    Span4Mux_h I__5952 (
            .O(N__24705),
            .I(N__24642));
    Span4Mux_v I__5951 (
            .O(N__24696),
            .I(N__24642));
    LocalMux I__5950 (
            .O(N__24693),
            .I(N__24642));
    LocalMux I__5949 (
            .O(N__24690),
            .I(N__24636));
    LocalMux I__5948 (
            .O(N__24687),
            .I(N__24636));
    InMux I__5947 (
            .O(N__24686),
            .I(N__24633));
    Span4Mux_v I__5946 (
            .O(N__24681),
            .I(N__24630));
    Span4Mux_v I__5945 (
            .O(N__24678),
            .I(N__24625));
    LocalMux I__5944 (
            .O(N__24675),
            .I(N__24625));
    LocalMux I__5943 (
            .O(N__24672),
            .I(N__24618));
    Span4Mux_v I__5942 (
            .O(N__24669),
            .I(N__24618));
    Span4Mux_v I__5941 (
            .O(N__24666),
            .I(N__24618));
    Span4Mux_v I__5940 (
            .O(N__24663),
            .I(N__24613));
    Span4Mux_v I__5939 (
            .O(N__24660),
            .I(N__24613));
    LocalMux I__5938 (
            .O(N__24657),
            .I(N__24606));
    LocalMux I__5937 (
            .O(N__24654),
            .I(N__24606));
    Span4Mux_h I__5936 (
            .O(N__24651),
            .I(N__24606));
    Span4Mux_h I__5935 (
            .O(N__24642),
            .I(N__24603));
    InMux I__5934 (
            .O(N__24641),
            .I(N__24600));
    Span12Mux_h I__5933 (
            .O(N__24636),
            .I(N__24597));
    LocalMux I__5932 (
            .O(N__24633),
            .I(N__24594));
    Span4Mux_v I__5931 (
            .O(N__24630),
            .I(N__24585));
    Span4Mux_v I__5930 (
            .O(N__24625),
            .I(N__24585));
    Span4Mux_h I__5929 (
            .O(N__24618),
            .I(N__24585));
    Span4Mux_h I__5928 (
            .O(N__24613),
            .I(N__24585));
    Span4Mux_h I__5927 (
            .O(N__24606),
            .I(N__24582));
    Span4Mux_h I__5926 (
            .O(N__24603),
            .I(N__24579));
    LocalMux I__5925 (
            .O(N__24600),
            .I(TX_ADDR_11));
    Odrv12 I__5924 (
            .O(N__24597),
            .I(TX_ADDR_11));
    Odrv12 I__5923 (
            .O(N__24594),
            .I(TX_ADDR_11));
    Odrv4 I__5922 (
            .O(N__24585),
            .I(TX_ADDR_11));
    Odrv4 I__5921 (
            .O(N__24582),
            .I(TX_ADDR_11));
    Odrv4 I__5920 (
            .O(N__24579),
            .I(TX_ADDR_11));
    InMux I__5919 (
            .O(N__24566),
            .I(N__24563));
    LocalMux I__5918 (
            .O(N__24563),
            .I(N__24560));
    Span4Mux_v I__5917 (
            .O(N__24560),
            .I(N__24557));
    Sp12to4 I__5916 (
            .O(N__24557),
            .I(N__24554));
    Odrv12 I__5915 (
            .O(N__24554),
            .I(\line_buffer.n538 ));
    InMux I__5914 (
            .O(N__24551),
            .I(N__24548));
    LocalMux I__5913 (
            .O(N__24548),
            .I(N__24545));
    Span4Mux_v I__5912 (
            .O(N__24545),
            .I(N__24542));
    Span4Mux_h I__5911 (
            .O(N__24542),
            .I(N__24539));
    Sp12to4 I__5910 (
            .O(N__24539),
            .I(N__24536));
    Span12Mux_v I__5909 (
            .O(N__24536),
            .I(N__24533));
    Odrv12 I__5908 (
            .O(N__24533),
            .I(\line_buffer.n530 ));
    InMux I__5907 (
            .O(N__24530),
            .I(N__24527));
    LocalMux I__5906 (
            .O(N__24527),
            .I(\line_buffer.n3542 ));
    SRMux I__5905 (
            .O(N__24524),
            .I(N__24518));
    SRMux I__5904 (
            .O(N__24523),
            .I(N__24515));
    SRMux I__5903 (
            .O(N__24522),
            .I(N__24509));
    SRMux I__5902 (
            .O(N__24521),
            .I(N__24506));
    LocalMux I__5901 (
            .O(N__24518),
            .I(N__24500));
    LocalMux I__5900 (
            .O(N__24515),
            .I(N__24500));
    SRMux I__5899 (
            .O(N__24514),
            .I(N__24497));
    IoInMux I__5898 (
            .O(N__24513),
            .I(N__24493));
    IoInMux I__5897 (
            .O(N__24512),
            .I(N__24490));
    LocalMux I__5896 (
            .O(N__24509),
            .I(N__24485));
    LocalMux I__5895 (
            .O(N__24506),
            .I(N__24482));
    SRMux I__5894 (
            .O(N__24505),
            .I(N__24479));
    Span4Mux_s2_v I__5893 (
            .O(N__24500),
            .I(N__24474));
    LocalMux I__5892 (
            .O(N__24497),
            .I(N__24474));
    SRMux I__5891 (
            .O(N__24496),
            .I(N__24471));
    LocalMux I__5890 (
            .O(N__24493),
            .I(N__24463));
    LocalMux I__5889 (
            .O(N__24490),
            .I(N__24463));
    SRMux I__5888 (
            .O(N__24489),
            .I(N__24459));
    SRMux I__5887 (
            .O(N__24488),
            .I(N__24456));
    Span4Mux_v I__5886 (
            .O(N__24485),
            .I(N__24447));
    Span4Mux_h I__5885 (
            .O(N__24482),
            .I(N__24447));
    LocalMux I__5884 (
            .O(N__24479),
            .I(N__24447));
    Span4Mux_v I__5883 (
            .O(N__24474),
            .I(N__24442));
    LocalMux I__5882 (
            .O(N__24471),
            .I(N__24442));
    SRMux I__5881 (
            .O(N__24470),
            .I(N__24439));
    SRMux I__5880 (
            .O(N__24469),
            .I(N__24436));
    SRMux I__5879 (
            .O(N__24468),
            .I(N__24432));
    IoSpan4Mux I__5878 (
            .O(N__24463),
            .I(N__24429));
    SRMux I__5877 (
            .O(N__24462),
            .I(N__24426));
    LocalMux I__5876 (
            .O(N__24459),
            .I(N__24419));
    LocalMux I__5875 (
            .O(N__24456),
            .I(N__24419));
    SRMux I__5874 (
            .O(N__24455),
            .I(N__24416));
    SRMux I__5873 (
            .O(N__24454),
            .I(N__24413));
    Span4Mux_v I__5872 (
            .O(N__24447),
            .I(N__24404));
    Span4Mux_v I__5871 (
            .O(N__24442),
            .I(N__24397));
    LocalMux I__5870 (
            .O(N__24439),
            .I(N__24397));
    LocalMux I__5869 (
            .O(N__24436),
            .I(N__24397));
    SRMux I__5868 (
            .O(N__24435),
            .I(N__24394));
    LocalMux I__5867 (
            .O(N__24432),
            .I(N__24391));
    IoSpan4Mux I__5866 (
            .O(N__24429),
            .I(N__24388));
    LocalMux I__5865 (
            .O(N__24426),
            .I(N__24385));
    SRMux I__5864 (
            .O(N__24425),
            .I(N__24382));
    SRMux I__5863 (
            .O(N__24424),
            .I(N__24379));
    Span4Mux_s2_v I__5862 (
            .O(N__24419),
            .I(N__24370));
    LocalMux I__5861 (
            .O(N__24416),
            .I(N__24370));
    LocalMux I__5860 (
            .O(N__24413),
            .I(N__24370));
    SRMux I__5859 (
            .O(N__24412),
            .I(N__24367));
    SRMux I__5858 (
            .O(N__24411),
            .I(N__24364));
    SRMux I__5857 (
            .O(N__24410),
            .I(N__24360));
    SRMux I__5856 (
            .O(N__24409),
            .I(N__24357));
    SRMux I__5855 (
            .O(N__24408),
            .I(N__24354));
    SRMux I__5854 (
            .O(N__24407),
            .I(N__24351));
    Span4Mux_v I__5853 (
            .O(N__24404),
            .I(N__24344));
    Span4Mux_v I__5852 (
            .O(N__24397),
            .I(N__24344));
    LocalMux I__5851 (
            .O(N__24394),
            .I(N__24344));
    Span4Mux_h I__5850 (
            .O(N__24391),
            .I(N__24339));
    Span4Mux_s3_v I__5849 (
            .O(N__24388),
            .I(N__24330));
    Span4Mux_s3_v I__5848 (
            .O(N__24385),
            .I(N__24330));
    LocalMux I__5847 (
            .O(N__24382),
            .I(N__24330));
    LocalMux I__5846 (
            .O(N__24379),
            .I(N__24330));
    SRMux I__5845 (
            .O(N__24378),
            .I(N__24327));
    SRMux I__5844 (
            .O(N__24377),
            .I(N__24324));
    Span4Mux_v I__5843 (
            .O(N__24370),
            .I(N__24315));
    LocalMux I__5842 (
            .O(N__24367),
            .I(N__24315));
    LocalMux I__5841 (
            .O(N__24364),
            .I(N__24315));
    SRMux I__5840 (
            .O(N__24363),
            .I(N__24312));
    LocalMux I__5839 (
            .O(N__24360),
            .I(N__24309));
    LocalMux I__5838 (
            .O(N__24357),
            .I(N__24306));
    LocalMux I__5837 (
            .O(N__24354),
            .I(N__24303));
    LocalMux I__5836 (
            .O(N__24351),
            .I(N__24300));
    Span4Mux_v I__5835 (
            .O(N__24344),
            .I(N__24297));
    SRMux I__5834 (
            .O(N__24343),
            .I(N__24294));
    SRMux I__5833 (
            .O(N__24342),
            .I(N__24291));
    Span4Mux_h I__5832 (
            .O(N__24339),
            .I(N__24288));
    Span4Mux_v I__5831 (
            .O(N__24330),
            .I(N__24281));
    LocalMux I__5830 (
            .O(N__24327),
            .I(N__24281));
    LocalMux I__5829 (
            .O(N__24324),
            .I(N__24281));
    SRMux I__5828 (
            .O(N__24323),
            .I(N__24278));
    SRMux I__5827 (
            .O(N__24322),
            .I(N__24275));
    Span4Mux_v I__5826 (
            .O(N__24315),
            .I(N__24270));
    LocalMux I__5825 (
            .O(N__24312),
            .I(N__24270));
    Span12Mux_s9_h I__5824 (
            .O(N__24309),
            .I(N__24266));
    Span12Mux_s9_h I__5823 (
            .O(N__24306),
            .I(N__24263));
    Span12Mux_h I__5822 (
            .O(N__24303),
            .I(N__24260));
    Span12Mux_h I__5821 (
            .O(N__24300),
            .I(N__24257));
    Sp12to4 I__5820 (
            .O(N__24297),
            .I(N__24252));
    LocalMux I__5819 (
            .O(N__24294),
            .I(N__24252));
    LocalMux I__5818 (
            .O(N__24291),
            .I(N__24249));
    Span4Mux_h I__5817 (
            .O(N__24288),
            .I(N__24246));
    Span4Mux_v I__5816 (
            .O(N__24281),
            .I(N__24241));
    LocalMux I__5815 (
            .O(N__24278),
            .I(N__24241));
    LocalMux I__5814 (
            .O(N__24275),
            .I(N__24238));
    Span4Mux_v I__5813 (
            .O(N__24270),
            .I(N__24235));
    SRMux I__5812 (
            .O(N__24269),
            .I(N__24232));
    Span12Mux_h I__5811 (
            .O(N__24266),
            .I(N__24227));
    Span12Mux_h I__5810 (
            .O(N__24263),
            .I(N__24227));
    Span12Mux_v I__5809 (
            .O(N__24260),
            .I(N__24220));
    Span12Mux_v I__5808 (
            .O(N__24257),
            .I(N__24220));
    Span12Mux_h I__5807 (
            .O(N__24252),
            .I(N__24220));
    Span4Mux_h I__5806 (
            .O(N__24249),
            .I(N__24217));
    Span4Mux_h I__5805 (
            .O(N__24246),
            .I(N__24210));
    Span4Mux_h I__5804 (
            .O(N__24241),
            .I(N__24210));
    Span4Mux_h I__5803 (
            .O(N__24238),
            .I(N__24210));
    Span4Mux_v I__5802 (
            .O(N__24235),
            .I(N__24205));
    LocalMux I__5801 (
            .O(N__24232),
            .I(N__24205));
    Odrv12 I__5800 (
            .O(N__24227),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__5799 (
            .O(N__24220),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5798 (
            .O(N__24217),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5797 (
            .O(N__24210),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5796 (
            .O(N__24205),
            .I(CONSTANT_ONE_NET));
    InMux I__5795 (
            .O(N__24194),
            .I(N__24191));
    LocalMux I__5794 (
            .O(N__24191),
            .I(N__24188));
    Odrv12 I__5793 (
            .O(N__24188),
            .I(TVP_VIDEO_c_9));
    InMux I__5792 (
            .O(N__24185),
            .I(N__24182));
    LocalMux I__5791 (
            .O(N__24182),
            .I(N__24179));
    Span4Mux_v I__5790 (
            .O(N__24179),
            .I(N__24176));
    Odrv4 I__5789 (
            .O(N__24176),
            .I(\tvp_video_buffer.BUFFER_0_9 ));
    InMux I__5788 (
            .O(N__24173),
            .I(N__24170));
    LocalMux I__5787 (
            .O(N__24170),
            .I(N__24149));
    ClkMux I__5786 (
            .O(N__24169),
            .I(N__23957));
    ClkMux I__5785 (
            .O(N__24168),
            .I(N__23957));
    ClkMux I__5784 (
            .O(N__24167),
            .I(N__23957));
    ClkMux I__5783 (
            .O(N__24166),
            .I(N__23957));
    ClkMux I__5782 (
            .O(N__24165),
            .I(N__23957));
    ClkMux I__5781 (
            .O(N__24164),
            .I(N__23957));
    ClkMux I__5780 (
            .O(N__24163),
            .I(N__23957));
    ClkMux I__5779 (
            .O(N__24162),
            .I(N__23957));
    ClkMux I__5778 (
            .O(N__24161),
            .I(N__23957));
    ClkMux I__5777 (
            .O(N__24160),
            .I(N__23957));
    ClkMux I__5776 (
            .O(N__24159),
            .I(N__23957));
    ClkMux I__5775 (
            .O(N__24158),
            .I(N__23957));
    ClkMux I__5774 (
            .O(N__24157),
            .I(N__23957));
    ClkMux I__5773 (
            .O(N__24156),
            .I(N__23957));
    ClkMux I__5772 (
            .O(N__24155),
            .I(N__23957));
    ClkMux I__5771 (
            .O(N__24154),
            .I(N__23957));
    ClkMux I__5770 (
            .O(N__24153),
            .I(N__23957));
    ClkMux I__5769 (
            .O(N__24152),
            .I(N__23957));
    Glb2LocalMux I__5768 (
            .O(N__24149),
            .I(N__23957));
    ClkMux I__5767 (
            .O(N__24148),
            .I(N__23957));
    ClkMux I__5766 (
            .O(N__24147),
            .I(N__23957));
    ClkMux I__5765 (
            .O(N__24146),
            .I(N__23957));
    ClkMux I__5764 (
            .O(N__24145),
            .I(N__23957));
    ClkMux I__5763 (
            .O(N__24144),
            .I(N__23957));
    ClkMux I__5762 (
            .O(N__24143),
            .I(N__23957));
    ClkMux I__5761 (
            .O(N__24142),
            .I(N__23957));
    ClkMux I__5760 (
            .O(N__24141),
            .I(N__23957));
    ClkMux I__5759 (
            .O(N__24140),
            .I(N__23957));
    ClkMux I__5758 (
            .O(N__24139),
            .I(N__23957));
    ClkMux I__5757 (
            .O(N__24138),
            .I(N__23957));
    ClkMux I__5756 (
            .O(N__24137),
            .I(N__23957));
    ClkMux I__5755 (
            .O(N__24136),
            .I(N__23957));
    ClkMux I__5754 (
            .O(N__24135),
            .I(N__23957));
    ClkMux I__5753 (
            .O(N__24134),
            .I(N__23957));
    ClkMux I__5752 (
            .O(N__24133),
            .I(N__23957));
    ClkMux I__5751 (
            .O(N__24132),
            .I(N__23957));
    ClkMux I__5750 (
            .O(N__24131),
            .I(N__23957));
    ClkMux I__5749 (
            .O(N__24130),
            .I(N__23957));
    ClkMux I__5748 (
            .O(N__24129),
            .I(N__23957));
    ClkMux I__5747 (
            .O(N__24128),
            .I(N__23957));
    ClkMux I__5746 (
            .O(N__24127),
            .I(N__23957));
    ClkMux I__5745 (
            .O(N__24126),
            .I(N__23957));
    ClkMux I__5744 (
            .O(N__24125),
            .I(N__23957));
    ClkMux I__5743 (
            .O(N__24124),
            .I(N__23957));
    ClkMux I__5742 (
            .O(N__24123),
            .I(N__23957));
    ClkMux I__5741 (
            .O(N__24122),
            .I(N__23957));
    ClkMux I__5740 (
            .O(N__24121),
            .I(N__23957));
    ClkMux I__5739 (
            .O(N__24120),
            .I(N__23957));
    ClkMux I__5738 (
            .O(N__24119),
            .I(N__23957));
    ClkMux I__5737 (
            .O(N__24118),
            .I(N__23957));
    ClkMux I__5736 (
            .O(N__24117),
            .I(N__23957));
    ClkMux I__5735 (
            .O(N__24116),
            .I(N__23957));
    ClkMux I__5734 (
            .O(N__24115),
            .I(N__23957));
    ClkMux I__5733 (
            .O(N__24114),
            .I(N__23957));
    ClkMux I__5732 (
            .O(N__24113),
            .I(N__23957));
    ClkMux I__5731 (
            .O(N__24112),
            .I(N__23957));
    ClkMux I__5730 (
            .O(N__24111),
            .I(N__23957));
    ClkMux I__5729 (
            .O(N__24110),
            .I(N__23957));
    ClkMux I__5728 (
            .O(N__24109),
            .I(N__23957));
    ClkMux I__5727 (
            .O(N__24108),
            .I(N__23957));
    ClkMux I__5726 (
            .O(N__24107),
            .I(N__23957));
    ClkMux I__5725 (
            .O(N__24106),
            .I(N__23957));
    ClkMux I__5724 (
            .O(N__24105),
            .I(N__23957));
    ClkMux I__5723 (
            .O(N__24104),
            .I(N__23957));
    ClkMux I__5722 (
            .O(N__24103),
            .I(N__23957));
    ClkMux I__5721 (
            .O(N__24102),
            .I(N__23957));
    ClkMux I__5720 (
            .O(N__24101),
            .I(N__23957));
    ClkMux I__5719 (
            .O(N__24100),
            .I(N__23957));
    ClkMux I__5718 (
            .O(N__24099),
            .I(N__23957));
    ClkMux I__5717 (
            .O(N__24098),
            .I(N__23957));
    GlobalMux I__5716 (
            .O(N__23957),
            .I(N__23954));
    gio2CtrlBuf I__5715 (
            .O(N__23954),
            .I(DEBUG_c_3_c));
    CascadeMux I__5714 (
            .O(N__23951),
            .I(N__23945));
    CascadeMux I__5713 (
            .O(N__23950),
            .I(N__23941));
    CascadeMux I__5712 (
            .O(N__23949),
            .I(N__23934));
    InMux I__5711 (
            .O(N__23948),
            .I(N__23929));
    InMux I__5710 (
            .O(N__23945),
            .I(N__23926));
    InMux I__5709 (
            .O(N__23944),
            .I(N__23923));
    InMux I__5708 (
            .O(N__23941),
            .I(N__23920));
    InMux I__5707 (
            .O(N__23940),
            .I(N__23914));
    InMux I__5706 (
            .O(N__23939),
            .I(N__23911));
    InMux I__5705 (
            .O(N__23938),
            .I(N__23908));
    InMux I__5704 (
            .O(N__23937),
            .I(N__23905));
    InMux I__5703 (
            .O(N__23934),
            .I(N__23902));
    CascadeMux I__5702 (
            .O(N__23933),
            .I(N__23899));
    InMux I__5701 (
            .O(N__23932),
            .I(N__23896));
    LocalMux I__5700 (
            .O(N__23929),
            .I(N__23891));
    LocalMux I__5699 (
            .O(N__23926),
            .I(N__23891));
    LocalMux I__5698 (
            .O(N__23923),
            .I(N__23886));
    LocalMux I__5697 (
            .O(N__23920),
            .I(N__23886));
    CascadeMux I__5696 (
            .O(N__23919),
            .I(N__23883));
    InMux I__5695 (
            .O(N__23918),
            .I(N__23880));
    InMux I__5694 (
            .O(N__23917),
            .I(N__23877));
    LocalMux I__5693 (
            .O(N__23914),
            .I(N__23874));
    LocalMux I__5692 (
            .O(N__23911),
            .I(N__23871));
    LocalMux I__5691 (
            .O(N__23908),
            .I(N__23864));
    LocalMux I__5690 (
            .O(N__23905),
            .I(N__23864));
    LocalMux I__5689 (
            .O(N__23902),
            .I(N__23864));
    InMux I__5688 (
            .O(N__23899),
            .I(N__23861));
    LocalMux I__5687 (
            .O(N__23896),
            .I(N__23856));
    Span4Mux_h I__5686 (
            .O(N__23891),
            .I(N__23856));
    Span4Mux_h I__5685 (
            .O(N__23886),
            .I(N__23853));
    InMux I__5684 (
            .O(N__23883),
            .I(N__23850));
    LocalMux I__5683 (
            .O(N__23880),
            .I(N__23847));
    LocalMux I__5682 (
            .O(N__23877),
            .I(N__23844));
    Span4Mux_v I__5681 (
            .O(N__23874),
            .I(N__23839));
    Span4Mux_h I__5680 (
            .O(N__23871),
            .I(N__23839));
    Span12Mux_h I__5679 (
            .O(N__23864),
            .I(N__23836));
    LocalMux I__5678 (
            .O(N__23861),
            .I(N__23827));
    Span4Mux_h I__5677 (
            .O(N__23856),
            .I(N__23827));
    Span4Mux_h I__5676 (
            .O(N__23853),
            .I(N__23827));
    LocalMux I__5675 (
            .O(N__23850),
            .I(N__23827));
    Span4Mux_h I__5674 (
            .O(N__23847),
            .I(N__23822));
    Span4Mux_h I__5673 (
            .O(N__23844),
            .I(N__23822));
    Odrv4 I__5672 (
            .O(N__23839),
            .I(TX_ADDR_13));
    Odrv12 I__5671 (
            .O(N__23836),
            .I(TX_ADDR_13));
    Odrv4 I__5670 (
            .O(N__23827),
            .I(TX_ADDR_13));
    Odrv4 I__5669 (
            .O(N__23822),
            .I(TX_ADDR_13));
    CascadeMux I__5668 (
            .O(N__23813),
            .I(\line_buffer.n3608_cascade_ ));
    InMux I__5667 (
            .O(N__23810),
            .I(N__23807));
    LocalMux I__5666 (
            .O(N__23807),
            .I(N__23804));
    Odrv4 I__5665 (
            .O(N__23804),
            .I(\line_buffer.n3576 ));
    InMux I__5664 (
            .O(N__23801),
            .I(N__23798));
    LocalMux I__5663 (
            .O(N__23798),
            .I(TX_DATA_6));
    IoInMux I__5662 (
            .O(N__23795),
            .I(N__23792));
    LocalMux I__5661 (
            .O(N__23792),
            .I(N__23787));
    IoInMux I__5660 (
            .O(N__23791),
            .I(N__23784));
    IoInMux I__5659 (
            .O(N__23790),
            .I(N__23781));
    Span4Mux_s3_h I__5658 (
            .O(N__23787),
            .I(N__23778));
    LocalMux I__5657 (
            .O(N__23784),
            .I(N__23775));
    LocalMux I__5656 (
            .O(N__23781),
            .I(N__23772));
    Span4Mux_v I__5655 (
            .O(N__23778),
            .I(N__23769));
    Span4Mux_s3_v I__5654 (
            .O(N__23775),
            .I(N__23766));
    IoSpan4Mux I__5653 (
            .O(N__23772),
            .I(N__23763));
    Span4Mux_v I__5652 (
            .O(N__23769),
            .I(N__23760));
    Span4Mux_h I__5651 (
            .O(N__23766),
            .I(N__23757));
    Span4Mux_s3_v I__5650 (
            .O(N__23763),
            .I(N__23754));
    Sp12to4 I__5649 (
            .O(N__23760),
            .I(N__23751));
    Sp12to4 I__5648 (
            .O(N__23757),
            .I(N__23748));
    Sp12to4 I__5647 (
            .O(N__23754),
            .I(N__23745));
    Span12Mux_h I__5646 (
            .O(N__23751),
            .I(N__23738));
    Span12Mux_s10_v I__5645 (
            .O(N__23748),
            .I(N__23738));
    Span12Mux_s10_v I__5644 (
            .O(N__23745),
            .I(N__23738));
    Odrv12 I__5643 (
            .O(N__23738),
            .I(n1815));
    ClkMux I__5642 (
            .O(N__23735),
            .I(N__23731));
    ClkMux I__5641 (
            .O(N__23734),
            .I(N__23725));
    LocalMux I__5640 (
            .O(N__23731),
            .I(N__23719));
    ClkMux I__5639 (
            .O(N__23730),
            .I(N__23716));
    ClkMux I__5638 (
            .O(N__23729),
            .I(N__23711));
    ClkMux I__5637 (
            .O(N__23728),
            .I(N__23705));
    LocalMux I__5636 (
            .O(N__23725),
            .I(N__23700));
    ClkMux I__5635 (
            .O(N__23724),
            .I(N__23697));
    ClkMux I__5634 (
            .O(N__23723),
            .I(N__23693));
    ClkMux I__5633 (
            .O(N__23722),
            .I(N__23690));
    Span4Mux_s2_v I__5632 (
            .O(N__23719),
            .I(N__23681));
    LocalMux I__5631 (
            .O(N__23716),
            .I(N__23681));
    ClkMux I__5630 (
            .O(N__23715),
            .I(N__23678));
    ClkMux I__5629 (
            .O(N__23714),
            .I(N__23674));
    LocalMux I__5628 (
            .O(N__23711),
            .I(N__23671));
    ClkMux I__5627 (
            .O(N__23710),
            .I(N__23668));
    ClkMux I__5626 (
            .O(N__23709),
            .I(N__23663));
    ClkMux I__5625 (
            .O(N__23708),
            .I(N__23660));
    LocalMux I__5624 (
            .O(N__23705),
            .I(N__23657));
    ClkMux I__5623 (
            .O(N__23704),
            .I(N__23653));
    ClkMux I__5622 (
            .O(N__23703),
            .I(N__23650));
    Span4Mux_v I__5621 (
            .O(N__23700),
            .I(N__23641));
    LocalMux I__5620 (
            .O(N__23697),
            .I(N__23641));
    ClkMux I__5619 (
            .O(N__23696),
            .I(N__23638));
    LocalMux I__5618 (
            .O(N__23693),
            .I(N__23631));
    LocalMux I__5617 (
            .O(N__23690),
            .I(N__23628));
    ClkMux I__5616 (
            .O(N__23689),
            .I(N__23625));
    ClkMux I__5615 (
            .O(N__23688),
            .I(N__23622));
    ClkMux I__5614 (
            .O(N__23687),
            .I(N__23617));
    ClkMux I__5613 (
            .O(N__23686),
            .I(N__23614));
    Span4Mux_v I__5612 (
            .O(N__23681),
            .I(N__23608));
    LocalMux I__5611 (
            .O(N__23678),
            .I(N__23608));
    ClkMux I__5610 (
            .O(N__23677),
            .I(N__23605));
    LocalMux I__5609 (
            .O(N__23674),
            .I(N__23595));
    Span4Mux_h I__5608 (
            .O(N__23671),
            .I(N__23590));
    LocalMux I__5607 (
            .O(N__23668),
            .I(N__23590));
    ClkMux I__5606 (
            .O(N__23667),
            .I(N__23587));
    ClkMux I__5605 (
            .O(N__23666),
            .I(N__23584));
    LocalMux I__5604 (
            .O(N__23663),
            .I(N__23581));
    LocalMux I__5603 (
            .O(N__23660),
            .I(N__23578));
    Span4Mux_h I__5602 (
            .O(N__23657),
            .I(N__23575));
    ClkMux I__5601 (
            .O(N__23656),
            .I(N__23572));
    LocalMux I__5600 (
            .O(N__23653),
            .I(N__23567));
    LocalMux I__5599 (
            .O(N__23650),
            .I(N__23564));
    ClkMux I__5598 (
            .O(N__23649),
            .I(N__23561));
    ClkMux I__5597 (
            .O(N__23648),
            .I(N__23557));
    ClkMux I__5596 (
            .O(N__23647),
            .I(N__23554));
    ClkMux I__5595 (
            .O(N__23646),
            .I(N__23547));
    Span4Mux_v I__5594 (
            .O(N__23641),
            .I(N__23542));
    LocalMux I__5593 (
            .O(N__23638),
            .I(N__23542));
    ClkMux I__5592 (
            .O(N__23637),
            .I(N__23539));
    ClkMux I__5591 (
            .O(N__23636),
            .I(N__23536));
    ClkMux I__5590 (
            .O(N__23635),
            .I(N__23533));
    ClkMux I__5589 (
            .O(N__23634),
            .I(N__23528));
    Span4Mux_s2_v I__5588 (
            .O(N__23631),
            .I(N__23520));
    Span4Mux_h I__5587 (
            .O(N__23628),
            .I(N__23520));
    LocalMux I__5586 (
            .O(N__23625),
            .I(N__23520));
    LocalMux I__5585 (
            .O(N__23622),
            .I(N__23517));
    ClkMux I__5584 (
            .O(N__23621),
            .I(N__23514));
    ClkMux I__5583 (
            .O(N__23620),
            .I(N__23511));
    LocalMux I__5582 (
            .O(N__23617),
            .I(N__23506));
    LocalMux I__5581 (
            .O(N__23614),
            .I(N__23503));
    ClkMux I__5580 (
            .O(N__23613),
            .I(N__23500));
    Span4Mux_v I__5579 (
            .O(N__23608),
            .I(N__23495));
    LocalMux I__5578 (
            .O(N__23605),
            .I(N__23495));
    ClkMux I__5577 (
            .O(N__23604),
            .I(N__23492));
    ClkMux I__5576 (
            .O(N__23603),
            .I(N__23489));
    ClkMux I__5575 (
            .O(N__23602),
            .I(N__23483));
    ClkMux I__5574 (
            .O(N__23601),
            .I(N__23479));
    ClkMux I__5573 (
            .O(N__23600),
            .I(N__23475));
    ClkMux I__5572 (
            .O(N__23599),
            .I(N__23471));
    ClkMux I__5571 (
            .O(N__23598),
            .I(N__23468));
    Span4Mux_h I__5570 (
            .O(N__23595),
            .I(N__23457));
    Span4Mux_h I__5569 (
            .O(N__23590),
            .I(N__23457));
    LocalMux I__5568 (
            .O(N__23587),
            .I(N__23457));
    LocalMux I__5567 (
            .O(N__23584),
            .I(N__23457));
    Span4Mux_v I__5566 (
            .O(N__23581),
            .I(N__23452));
    Span4Mux_h I__5565 (
            .O(N__23578),
            .I(N__23452));
    Span4Mux_v I__5564 (
            .O(N__23575),
            .I(N__23447));
    LocalMux I__5563 (
            .O(N__23572),
            .I(N__23447));
    ClkMux I__5562 (
            .O(N__23571),
            .I(N__23444));
    ClkMux I__5561 (
            .O(N__23570),
            .I(N__23441));
    Span4Mux_h I__5560 (
            .O(N__23567),
            .I(N__23436));
    Span4Mux_v I__5559 (
            .O(N__23564),
            .I(N__23431));
    LocalMux I__5558 (
            .O(N__23561),
            .I(N__23431));
    ClkMux I__5557 (
            .O(N__23560),
            .I(N__23428));
    LocalMux I__5556 (
            .O(N__23557),
            .I(N__23425));
    LocalMux I__5555 (
            .O(N__23554),
            .I(N__23422));
    ClkMux I__5554 (
            .O(N__23553),
            .I(N__23419));
    ClkMux I__5553 (
            .O(N__23552),
            .I(N__23414));
    ClkMux I__5552 (
            .O(N__23551),
            .I(N__23410));
    ClkMux I__5551 (
            .O(N__23550),
            .I(N__23406));
    LocalMux I__5550 (
            .O(N__23547),
            .I(N__23400));
    Span4Mux_h I__5549 (
            .O(N__23542),
            .I(N__23395));
    LocalMux I__5548 (
            .O(N__23539),
            .I(N__23395));
    LocalMux I__5547 (
            .O(N__23536),
            .I(N__23390));
    LocalMux I__5546 (
            .O(N__23533),
            .I(N__23390));
    ClkMux I__5545 (
            .O(N__23532),
            .I(N__23387));
    ClkMux I__5544 (
            .O(N__23531),
            .I(N__23384));
    LocalMux I__5543 (
            .O(N__23528),
            .I(N__23380));
    ClkMux I__5542 (
            .O(N__23527),
            .I(N__23377));
    Span4Mux_v I__5541 (
            .O(N__23520),
            .I(N__23368));
    Span4Mux_h I__5540 (
            .O(N__23517),
            .I(N__23368));
    LocalMux I__5539 (
            .O(N__23514),
            .I(N__23368));
    LocalMux I__5538 (
            .O(N__23511),
            .I(N__23365));
    ClkMux I__5537 (
            .O(N__23510),
            .I(N__23362));
    ClkMux I__5536 (
            .O(N__23509),
            .I(N__23359));
    Span4Mux_v I__5535 (
            .O(N__23506),
            .I(N__23350));
    Span4Mux_h I__5534 (
            .O(N__23503),
            .I(N__23350));
    LocalMux I__5533 (
            .O(N__23500),
            .I(N__23350));
    Span4Mux_h I__5532 (
            .O(N__23495),
            .I(N__23343));
    LocalMux I__5531 (
            .O(N__23492),
            .I(N__23343));
    LocalMux I__5530 (
            .O(N__23489),
            .I(N__23343));
    ClkMux I__5529 (
            .O(N__23488),
            .I(N__23340));
    ClkMux I__5528 (
            .O(N__23487),
            .I(N__23337));
    ClkMux I__5527 (
            .O(N__23486),
            .I(N__23332));
    LocalMux I__5526 (
            .O(N__23483),
            .I(N__23328));
    ClkMux I__5525 (
            .O(N__23482),
            .I(N__23325));
    LocalMux I__5524 (
            .O(N__23479),
            .I(N__23321));
    ClkMux I__5523 (
            .O(N__23478),
            .I(N__23318));
    LocalMux I__5522 (
            .O(N__23475),
            .I(N__23315));
    ClkMux I__5521 (
            .O(N__23474),
            .I(N__23312));
    LocalMux I__5520 (
            .O(N__23471),
            .I(N__23309));
    LocalMux I__5519 (
            .O(N__23468),
            .I(N__23306));
    ClkMux I__5518 (
            .O(N__23467),
            .I(N__23303));
    ClkMux I__5517 (
            .O(N__23466),
            .I(N__23299));
    Span4Mux_h I__5516 (
            .O(N__23457),
            .I(N__23295));
    Span4Mux_h I__5515 (
            .O(N__23452),
            .I(N__23288));
    Span4Mux_v I__5514 (
            .O(N__23447),
            .I(N__23288));
    LocalMux I__5513 (
            .O(N__23444),
            .I(N__23288));
    LocalMux I__5512 (
            .O(N__23441),
            .I(N__23285));
    ClkMux I__5511 (
            .O(N__23440),
            .I(N__23282));
    ClkMux I__5510 (
            .O(N__23439),
            .I(N__23279));
    Span4Mux_v I__5509 (
            .O(N__23436),
            .I(N__23271));
    Span4Mux_h I__5508 (
            .O(N__23431),
            .I(N__23271));
    LocalMux I__5507 (
            .O(N__23428),
            .I(N__23271));
    Span4Mux_v I__5506 (
            .O(N__23425),
            .I(N__23264));
    Span4Mux_v I__5505 (
            .O(N__23422),
            .I(N__23264));
    LocalMux I__5504 (
            .O(N__23419),
            .I(N__23264));
    ClkMux I__5503 (
            .O(N__23418),
            .I(N__23261));
    ClkMux I__5502 (
            .O(N__23417),
            .I(N__23258));
    LocalMux I__5501 (
            .O(N__23414),
            .I(N__23254));
    ClkMux I__5500 (
            .O(N__23413),
            .I(N__23250));
    LocalMux I__5499 (
            .O(N__23410),
            .I(N__23245));
    ClkMux I__5498 (
            .O(N__23409),
            .I(N__23242));
    LocalMux I__5497 (
            .O(N__23406),
            .I(N__23239));
    ClkMux I__5496 (
            .O(N__23405),
            .I(N__23236));
    ClkMux I__5495 (
            .O(N__23404),
            .I(N__23233));
    ClkMux I__5494 (
            .O(N__23403),
            .I(N__23229));
    Span4Mux_h I__5493 (
            .O(N__23400),
            .I(N__23216));
    Span4Mux_v I__5492 (
            .O(N__23395),
            .I(N__23216));
    Span4Mux_h I__5491 (
            .O(N__23390),
            .I(N__23216));
    LocalMux I__5490 (
            .O(N__23387),
            .I(N__23216));
    LocalMux I__5489 (
            .O(N__23384),
            .I(N__23216));
    ClkMux I__5488 (
            .O(N__23383),
            .I(N__23213));
    Span4Mux_v I__5487 (
            .O(N__23380),
            .I(N__23208));
    LocalMux I__5486 (
            .O(N__23377),
            .I(N__23208));
    ClkMux I__5485 (
            .O(N__23376),
            .I(N__23205));
    ClkMux I__5484 (
            .O(N__23375),
            .I(N__23202));
    Span4Mux_v I__5483 (
            .O(N__23368),
            .I(N__23194));
    Span4Mux_h I__5482 (
            .O(N__23365),
            .I(N__23194));
    LocalMux I__5481 (
            .O(N__23362),
            .I(N__23194));
    LocalMux I__5480 (
            .O(N__23359),
            .I(N__23191));
    ClkMux I__5479 (
            .O(N__23358),
            .I(N__23188));
    ClkMux I__5478 (
            .O(N__23357),
            .I(N__23185));
    Span4Mux_h I__5477 (
            .O(N__23350),
            .I(N__23177));
    Span4Mux_v I__5476 (
            .O(N__23343),
            .I(N__23177));
    LocalMux I__5475 (
            .O(N__23340),
            .I(N__23177));
    LocalMux I__5474 (
            .O(N__23337),
            .I(N__23174));
    ClkMux I__5473 (
            .O(N__23336),
            .I(N__23171));
    ClkMux I__5472 (
            .O(N__23335),
            .I(N__23168));
    LocalMux I__5471 (
            .O(N__23332),
            .I(N__23165));
    ClkMux I__5470 (
            .O(N__23331),
            .I(N__23162));
    Span4Mux_v I__5469 (
            .O(N__23328),
            .I(N__23157));
    LocalMux I__5468 (
            .O(N__23325),
            .I(N__23157));
    ClkMux I__5467 (
            .O(N__23324),
            .I(N__23154));
    Span4Mux_v I__5466 (
            .O(N__23321),
            .I(N__23149));
    LocalMux I__5465 (
            .O(N__23318),
            .I(N__23149));
    Span4Mux_h I__5464 (
            .O(N__23315),
            .I(N__23144));
    LocalMux I__5463 (
            .O(N__23312),
            .I(N__23144));
    Span4Mux_v I__5462 (
            .O(N__23309),
            .I(N__23137));
    Span4Mux_h I__5461 (
            .O(N__23306),
            .I(N__23137));
    LocalMux I__5460 (
            .O(N__23303),
            .I(N__23137));
    ClkMux I__5459 (
            .O(N__23302),
            .I(N__23134));
    LocalMux I__5458 (
            .O(N__23299),
            .I(N__23129));
    ClkMux I__5457 (
            .O(N__23298),
            .I(N__23126));
    Span4Mux_v I__5456 (
            .O(N__23295),
            .I(N__23118));
    Span4Mux_h I__5455 (
            .O(N__23288),
            .I(N__23118));
    Span4Mux_h I__5454 (
            .O(N__23285),
            .I(N__23118));
    LocalMux I__5453 (
            .O(N__23282),
            .I(N__23115));
    LocalMux I__5452 (
            .O(N__23279),
            .I(N__23112));
    IoInMux I__5451 (
            .O(N__23278),
            .I(N__23109));
    Span4Mux_h I__5450 (
            .O(N__23271),
            .I(N__23106));
    Span4Mux_h I__5449 (
            .O(N__23264),
            .I(N__23099));
    LocalMux I__5448 (
            .O(N__23261),
            .I(N__23099));
    LocalMux I__5447 (
            .O(N__23258),
            .I(N__23099));
    ClkMux I__5446 (
            .O(N__23257),
            .I(N__23096));
    Span4Mux_h I__5445 (
            .O(N__23254),
            .I(N__23093));
    ClkMux I__5444 (
            .O(N__23253),
            .I(N__23090));
    LocalMux I__5443 (
            .O(N__23250),
            .I(N__23087));
    ClkMux I__5442 (
            .O(N__23249),
            .I(N__23084));
    ClkMux I__5441 (
            .O(N__23248),
            .I(N__23080));
    Span4Mux_v I__5440 (
            .O(N__23245),
            .I(N__23075));
    LocalMux I__5439 (
            .O(N__23242),
            .I(N__23075));
    Span4Mux_v I__5438 (
            .O(N__23239),
            .I(N__23068));
    LocalMux I__5437 (
            .O(N__23236),
            .I(N__23068));
    LocalMux I__5436 (
            .O(N__23233),
            .I(N__23068));
    ClkMux I__5435 (
            .O(N__23232),
            .I(N__23065));
    LocalMux I__5434 (
            .O(N__23229),
            .I(N__23062));
    ClkMux I__5433 (
            .O(N__23228),
            .I(N__23059));
    ClkMux I__5432 (
            .O(N__23227),
            .I(N__23056));
    Span4Mux_h I__5431 (
            .O(N__23216),
            .I(N__23051));
    LocalMux I__5430 (
            .O(N__23213),
            .I(N__23051));
    Span4Mux_h I__5429 (
            .O(N__23208),
            .I(N__23046));
    LocalMux I__5428 (
            .O(N__23205),
            .I(N__23046));
    LocalMux I__5427 (
            .O(N__23202),
            .I(N__23043));
    ClkMux I__5426 (
            .O(N__23201),
            .I(N__23040));
    Span4Mux_v I__5425 (
            .O(N__23194),
            .I(N__23030));
    Span4Mux_h I__5424 (
            .O(N__23191),
            .I(N__23030));
    LocalMux I__5423 (
            .O(N__23188),
            .I(N__23030));
    LocalMux I__5422 (
            .O(N__23185),
            .I(N__23027));
    ClkMux I__5421 (
            .O(N__23184),
            .I(N__23024));
    Span4Mux_v I__5420 (
            .O(N__23177),
            .I(N__23020));
    Span4Mux_v I__5419 (
            .O(N__23174),
            .I(N__23015));
    LocalMux I__5418 (
            .O(N__23171),
            .I(N__23015));
    LocalMux I__5417 (
            .O(N__23168),
            .I(N__23012));
    Span4Mux_v I__5416 (
            .O(N__23165),
            .I(N__23003));
    LocalMux I__5415 (
            .O(N__23162),
            .I(N__23003));
    Span4Mux_v I__5414 (
            .O(N__23157),
            .I(N__23003));
    LocalMux I__5413 (
            .O(N__23154),
            .I(N__23003));
    Span4Mux_h I__5412 (
            .O(N__23149),
            .I(N__22994));
    Span4Mux_v I__5411 (
            .O(N__23144),
            .I(N__22994));
    Span4Mux_h I__5410 (
            .O(N__23137),
            .I(N__22994));
    LocalMux I__5409 (
            .O(N__23134),
            .I(N__22994));
    ClkMux I__5408 (
            .O(N__23133),
            .I(N__22991));
    ClkMux I__5407 (
            .O(N__23132),
            .I(N__22988));
    Span4Mux_v I__5406 (
            .O(N__23129),
            .I(N__22982));
    LocalMux I__5405 (
            .O(N__23126),
            .I(N__22982));
    ClkMux I__5404 (
            .O(N__23125),
            .I(N__22979));
    Span4Mux_v I__5403 (
            .O(N__23118),
            .I(N__22972));
    Span4Mux_h I__5402 (
            .O(N__23115),
            .I(N__22972));
    Span4Mux_h I__5401 (
            .O(N__23112),
            .I(N__22972));
    LocalMux I__5400 (
            .O(N__23109),
            .I(N__22969));
    Span4Mux_v I__5399 (
            .O(N__23106),
            .I(N__22964));
    Span4Mux_h I__5398 (
            .O(N__23099),
            .I(N__22964));
    LocalMux I__5397 (
            .O(N__23096),
            .I(N__22961));
    Span4Mux_v I__5396 (
            .O(N__23093),
            .I(N__22956));
    LocalMux I__5395 (
            .O(N__23090),
            .I(N__22956));
    Span4Mux_h I__5394 (
            .O(N__23087),
            .I(N__22952));
    LocalMux I__5393 (
            .O(N__23084),
            .I(N__22949));
    ClkMux I__5392 (
            .O(N__23083),
            .I(N__22946));
    LocalMux I__5391 (
            .O(N__23080),
            .I(N__22943));
    Span4Mux_v I__5390 (
            .O(N__23075),
            .I(N__22936));
    Span4Mux_h I__5389 (
            .O(N__23068),
            .I(N__22936));
    LocalMux I__5388 (
            .O(N__23065),
            .I(N__22936));
    Span4Mux_h I__5387 (
            .O(N__23062),
            .I(N__22931));
    LocalMux I__5386 (
            .O(N__23059),
            .I(N__22931));
    LocalMux I__5385 (
            .O(N__23056),
            .I(N__22928));
    Span4Mux_v I__5384 (
            .O(N__23051),
            .I(N__22919));
    Span4Mux_h I__5383 (
            .O(N__23046),
            .I(N__22919));
    Span4Mux_h I__5382 (
            .O(N__23043),
            .I(N__22919));
    LocalMux I__5381 (
            .O(N__23040),
            .I(N__22919));
    ClkMux I__5380 (
            .O(N__23039),
            .I(N__22916));
    ClkMux I__5379 (
            .O(N__23038),
            .I(N__22913));
    ClkMux I__5378 (
            .O(N__23037),
            .I(N__22909));
    Span4Mux_v I__5377 (
            .O(N__23030),
            .I(N__22901));
    Span4Mux_h I__5376 (
            .O(N__23027),
            .I(N__22901));
    LocalMux I__5375 (
            .O(N__23024),
            .I(N__22901));
    ClkMux I__5374 (
            .O(N__23023),
            .I(N__22898));
    Span4Mux_v I__5373 (
            .O(N__23020),
            .I(N__22895));
    Span4Mux_v I__5372 (
            .O(N__23015),
            .I(N__22892));
    Span4Mux_v I__5371 (
            .O(N__23012),
            .I(N__22887));
    Span4Mux_h I__5370 (
            .O(N__23003),
            .I(N__22887));
    Span4Mux_h I__5369 (
            .O(N__22994),
            .I(N__22880));
    LocalMux I__5368 (
            .O(N__22991),
            .I(N__22880));
    LocalMux I__5367 (
            .O(N__22988),
            .I(N__22880));
    ClkMux I__5366 (
            .O(N__22987),
            .I(N__22877));
    Span4Mux_h I__5365 (
            .O(N__22982),
            .I(N__22873));
    LocalMux I__5364 (
            .O(N__22979),
            .I(N__22870));
    Span4Mux_v I__5363 (
            .O(N__22972),
            .I(N__22866));
    IoSpan4Mux I__5362 (
            .O(N__22969),
            .I(N__22863));
    Span4Mux_v I__5361 (
            .O(N__22964),
            .I(N__22858));
    Span4Mux_h I__5360 (
            .O(N__22961),
            .I(N__22858));
    Span4Mux_h I__5359 (
            .O(N__22956),
            .I(N__22855));
    ClkMux I__5358 (
            .O(N__22955),
            .I(N__22852));
    Span4Mux_v I__5357 (
            .O(N__22952),
            .I(N__22847));
    Span4Mux_h I__5356 (
            .O(N__22949),
            .I(N__22847));
    LocalMux I__5355 (
            .O(N__22946),
            .I(N__22844));
    Span4Mux_h I__5354 (
            .O(N__22943),
            .I(N__22841));
    Span4Mux_v I__5353 (
            .O(N__22936),
            .I(N__22830));
    Span4Mux_h I__5352 (
            .O(N__22931),
            .I(N__22830));
    Span4Mux_h I__5351 (
            .O(N__22928),
            .I(N__22830));
    Span4Mux_v I__5350 (
            .O(N__22919),
            .I(N__22830));
    LocalMux I__5349 (
            .O(N__22916),
            .I(N__22830));
    LocalMux I__5348 (
            .O(N__22913),
            .I(N__22827));
    ClkMux I__5347 (
            .O(N__22912),
            .I(N__22824));
    LocalMux I__5346 (
            .O(N__22909),
            .I(N__22821));
    ClkMux I__5345 (
            .O(N__22908),
            .I(N__22818));
    Span4Mux_v I__5344 (
            .O(N__22901),
            .I(N__22815));
    LocalMux I__5343 (
            .O(N__22898),
            .I(N__22812));
    Span4Mux_h I__5342 (
            .O(N__22895),
            .I(N__22807));
    Span4Mux_v I__5341 (
            .O(N__22892),
            .I(N__22807));
    Span4Mux_h I__5340 (
            .O(N__22887),
            .I(N__22800));
    Span4Mux_v I__5339 (
            .O(N__22880),
            .I(N__22800));
    LocalMux I__5338 (
            .O(N__22877),
            .I(N__22800));
    ClkMux I__5337 (
            .O(N__22876),
            .I(N__22797));
    Span4Mux_h I__5336 (
            .O(N__22873),
            .I(N__22792));
    Span4Mux_v I__5335 (
            .O(N__22870),
            .I(N__22792));
    ClkMux I__5334 (
            .O(N__22869),
            .I(N__22789));
    Span4Mux_v I__5333 (
            .O(N__22866),
            .I(N__22786));
    IoSpan4Mux I__5332 (
            .O(N__22863),
            .I(N__22783));
    Span4Mux_v I__5331 (
            .O(N__22858),
            .I(N__22780));
    Span4Mux_h I__5330 (
            .O(N__22855),
            .I(N__22777));
    LocalMux I__5329 (
            .O(N__22852),
            .I(N__22774));
    Span4Mux_h I__5328 (
            .O(N__22847),
            .I(N__22771));
    Span4Mux_h I__5327 (
            .O(N__22844),
            .I(N__22768));
    Span4Mux_v I__5326 (
            .O(N__22841),
            .I(N__22761));
    Span4Mux_v I__5325 (
            .O(N__22830),
            .I(N__22761));
    Span4Mux_h I__5324 (
            .O(N__22827),
            .I(N__22761));
    LocalMux I__5323 (
            .O(N__22824),
            .I(N__22758));
    Span12Mux_h I__5322 (
            .O(N__22821),
            .I(N__22753));
    LocalMux I__5321 (
            .O(N__22818),
            .I(N__22753));
    Sp12to4 I__5320 (
            .O(N__22815),
            .I(N__22746));
    Sp12to4 I__5319 (
            .O(N__22812),
            .I(N__22746));
    Sp12to4 I__5318 (
            .O(N__22807),
            .I(N__22746));
    Span4Mux_v I__5317 (
            .O(N__22800),
            .I(N__22737));
    LocalMux I__5316 (
            .O(N__22797),
            .I(N__22737));
    Span4Mux_v I__5315 (
            .O(N__22792),
            .I(N__22737));
    LocalMux I__5314 (
            .O(N__22789),
            .I(N__22737));
    IoSpan4Mux I__5313 (
            .O(N__22786),
            .I(N__22732));
    IoSpan4Mux I__5312 (
            .O(N__22783),
            .I(N__22732));
    Span4Mux_v I__5311 (
            .O(N__22780),
            .I(N__22729));
    Span4Mux_h I__5310 (
            .O(N__22777),
            .I(N__22726));
    Span12Mux_h I__5309 (
            .O(N__22774),
            .I(N__22723));
    Span4Mux_h I__5308 (
            .O(N__22771),
            .I(N__22716));
    Span4Mux_h I__5307 (
            .O(N__22768),
            .I(N__22716));
    Span4Mux_v I__5306 (
            .O(N__22761),
            .I(N__22716));
    Span12Mux_h I__5305 (
            .O(N__22758),
            .I(N__22707));
    Span12Mux_v I__5304 (
            .O(N__22753),
            .I(N__22707));
    Span12Mux_h I__5303 (
            .O(N__22746),
            .I(N__22707));
    Sp12to4 I__5302 (
            .O(N__22737),
            .I(N__22707));
    Odrv4 I__5301 (
            .O(N__22732),
            .I(ADV_CLK_c));
    Odrv4 I__5300 (
            .O(N__22729),
            .I(ADV_CLK_c));
    Odrv4 I__5299 (
            .O(N__22726),
            .I(ADV_CLK_c));
    Odrv12 I__5298 (
            .O(N__22723),
            .I(ADV_CLK_c));
    Odrv4 I__5297 (
            .O(N__22716),
            .I(ADV_CLK_c));
    Odrv12 I__5296 (
            .O(N__22707),
            .I(ADV_CLK_c));
    SRMux I__5295 (
            .O(N__22694),
            .I(N__22689));
    SRMux I__5294 (
            .O(N__22693),
            .I(N__22684));
    SRMux I__5293 (
            .O(N__22692),
            .I(N__22681));
    LocalMux I__5292 (
            .O(N__22689),
            .I(N__22677));
    SRMux I__5291 (
            .O(N__22688),
            .I(N__22674));
    SRMux I__5290 (
            .O(N__22687),
            .I(N__22671));
    LocalMux I__5289 (
            .O(N__22684),
            .I(N__22667));
    LocalMux I__5288 (
            .O(N__22681),
            .I(N__22664));
    SRMux I__5287 (
            .O(N__22680),
            .I(N__22661));
    Span4Mux_h I__5286 (
            .O(N__22677),
            .I(N__22656));
    LocalMux I__5285 (
            .O(N__22674),
            .I(N__22656));
    LocalMux I__5284 (
            .O(N__22671),
            .I(N__22653));
    SRMux I__5283 (
            .O(N__22670),
            .I(N__22650));
    Span4Mux_v I__5282 (
            .O(N__22667),
            .I(N__22646));
    Span4Mux_v I__5281 (
            .O(N__22664),
            .I(N__22641));
    LocalMux I__5280 (
            .O(N__22661),
            .I(N__22641));
    Span4Mux_h I__5279 (
            .O(N__22656),
            .I(N__22634));
    Span4Mux_h I__5278 (
            .O(N__22653),
            .I(N__22634));
    LocalMux I__5277 (
            .O(N__22650),
            .I(N__22634));
    SRMux I__5276 (
            .O(N__22649),
            .I(N__22631));
    Span4Mux_h I__5275 (
            .O(N__22646),
            .I(N__22626));
    Span4Mux_v I__5274 (
            .O(N__22641),
            .I(N__22626));
    Span4Mux_v I__5273 (
            .O(N__22634),
            .I(N__22623));
    LocalMux I__5272 (
            .O(N__22631),
            .I(N__22620));
    Odrv4 I__5271 (
            .O(N__22626),
            .I(\transmit_module.n2388 ));
    Odrv4 I__5270 (
            .O(N__22623),
            .I(\transmit_module.n2388 ));
    Odrv12 I__5269 (
            .O(N__22620),
            .I(\transmit_module.n2388 ));
    InMux I__5268 (
            .O(N__22613),
            .I(N__22610));
    LocalMux I__5267 (
            .O(N__22610),
            .I(N__22607));
    Span4Mux_v I__5266 (
            .O(N__22607),
            .I(N__22604));
    Sp12to4 I__5265 (
            .O(N__22604),
            .I(N__22601));
    Odrv12 I__5264 (
            .O(N__22601),
            .I(\line_buffer.n596 ));
    InMux I__5263 (
            .O(N__22598),
            .I(N__22595));
    LocalMux I__5262 (
            .O(N__22595),
            .I(N__22592));
    Span4Mux_h I__5261 (
            .O(N__22592),
            .I(N__22589));
    Span4Mux_v I__5260 (
            .O(N__22589),
            .I(N__22586));
    Span4Mux_v I__5259 (
            .O(N__22586),
            .I(N__22583));
    Span4Mux_h I__5258 (
            .O(N__22583),
            .I(N__22580));
    Odrv4 I__5257 (
            .O(N__22580),
            .I(\line_buffer.n588 ));
    InMux I__5256 (
            .O(N__22577),
            .I(N__22574));
    LocalMux I__5255 (
            .O(N__22574),
            .I(\line_buffer.n3644 ));
    InMux I__5254 (
            .O(N__22571),
            .I(N__22568));
    LocalMux I__5253 (
            .O(N__22568),
            .I(N__22565));
    Span4Mux_h I__5252 (
            .O(N__22565),
            .I(N__22562));
    Span4Mux_h I__5251 (
            .O(N__22562),
            .I(N__22559));
    Odrv4 I__5250 (
            .O(N__22559),
            .I(\line_buffer.n473 ));
    InMux I__5249 (
            .O(N__22556),
            .I(N__22553));
    LocalMux I__5248 (
            .O(N__22553),
            .I(N__22550));
    Span4Mux_v I__5247 (
            .O(N__22550),
            .I(N__22547));
    Sp12to4 I__5246 (
            .O(N__22547),
            .I(N__22544));
    Odrv12 I__5245 (
            .O(N__22544),
            .I(\line_buffer.n465 ));
    InMux I__5244 (
            .O(N__22541),
            .I(N__22538));
    LocalMux I__5243 (
            .O(N__22538),
            .I(N__22535));
    Odrv12 I__5242 (
            .O(N__22535),
            .I(\line_buffer.n3575 ));
    InMux I__5241 (
            .O(N__22532),
            .I(N__22529));
    LocalMux I__5240 (
            .O(N__22529),
            .I(N__22526));
    Odrv12 I__5239 (
            .O(N__22526),
            .I(\tvp_video_buffer.BUFFER_1_9 ));
    InMux I__5238 (
            .O(N__22523),
            .I(N__22520));
    LocalMux I__5237 (
            .O(N__22520),
            .I(N__22514));
    InMux I__5236 (
            .O(N__22519),
            .I(N__22510));
    InMux I__5235 (
            .O(N__22518),
            .I(N__22507));
    InMux I__5234 (
            .O(N__22517),
            .I(N__22503));
    Span4Mux_s2_v I__5233 (
            .O(N__22514),
            .I(N__22500));
    InMux I__5232 (
            .O(N__22513),
            .I(N__22497));
    LocalMux I__5231 (
            .O(N__22510),
            .I(N__22493));
    LocalMux I__5230 (
            .O(N__22507),
            .I(N__22490));
    InMux I__5229 (
            .O(N__22506),
            .I(N__22487));
    LocalMux I__5228 (
            .O(N__22503),
            .I(N__22484));
    Span4Mux_v I__5227 (
            .O(N__22500),
            .I(N__22478));
    LocalMux I__5226 (
            .O(N__22497),
            .I(N__22478));
    InMux I__5225 (
            .O(N__22496),
            .I(N__22475));
    Span4Mux_h I__5224 (
            .O(N__22493),
            .I(N__22472));
    Span4Mux_v I__5223 (
            .O(N__22490),
            .I(N__22469));
    LocalMux I__5222 (
            .O(N__22487),
            .I(N__22466));
    Span4Mux_v I__5221 (
            .O(N__22484),
            .I(N__22463));
    InMux I__5220 (
            .O(N__22483),
            .I(N__22460));
    Span4Mux_h I__5219 (
            .O(N__22478),
            .I(N__22457));
    LocalMux I__5218 (
            .O(N__22475),
            .I(N__22453));
    Span4Mux_v I__5217 (
            .O(N__22472),
            .I(N__22450));
    Span4Mux_v I__5216 (
            .O(N__22469),
            .I(N__22445));
    Span4Mux_h I__5215 (
            .O(N__22466),
            .I(N__22445));
    Span4Mux_v I__5214 (
            .O(N__22463),
            .I(N__22440));
    LocalMux I__5213 (
            .O(N__22460),
            .I(N__22440));
    Span4Mux_h I__5212 (
            .O(N__22457),
            .I(N__22437));
    InMux I__5211 (
            .O(N__22456),
            .I(N__22434));
    Span12Mux_h I__5210 (
            .O(N__22453),
            .I(N__22431));
    Sp12to4 I__5209 (
            .O(N__22450),
            .I(N__22428));
    Span4Mux_v I__5208 (
            .O(N__22445),
            .I(N__22423));
    Span4Mux_v I__5207 (
            .O(N__22440),
            .I(N__22423));
    Sp12to4 I__5206 (
            .O(N__22437),
            .I(N__22418));
    LocalMux I__5205 (
            .O(N__22434),
            .I(N__22418));
    Span12Mux_v I__5204 (
            .O(N__22431),
            .I(N__22409));
    Span12Mux_h I__5203 (
            .O(N__22428),
            .I(N__22409));
    Sp12to4 I__5202 (
            .O(N__22423),
            .I(N__22409));
    Span12Mux_v I__5201 (
            .O(N__22418),
            .I(N__22409));
    Odrv12 I__5200 (
            .O(N__22409),
            .I(RX_DATA_5));
    InMux I__5199 (
            .O(N__22406),
            .I(N__22403));
    LocalMux I__5198 (
            .O(N__22403),
            .I(N__22400));
    Span12Mux_v I__5197 (
            .O(N__22400),
            .I(N__22397));
    Odrv12 I__5196 (
            .O(N__22397),
            .I(\line_buffer.n601 ));
    CascadeMux I__5195 (
            .O(N__22394),
            .I(N__22385));
    CascadeMux I__5194 (
            .O(N__22393),
            .I(N__22382));
    CascadeMux I__5193 (
            .O(N__22392),
            .I(N__22378));
    InMux I__5192 (
            .O(N__22391),
            .I(N__22369));
    InMux I__5191 (
            .O(N__22390),
            .I(N__22366));
    InMux I__5190 (
            .O(N__22389),
            .I(N__22363));
    InMux I__5189 (
            .O(N__22388),
            .I(N__22360));
    InMux I__5188 (
            .O(N__22385),
            .I(N__22357));
    InMux I__5187 (
            .O(N__22382),
            .I(N__22354));
    CascadeMux I__5186 (
            .O(N__22381),
            .I(N__22351));
    InMux I__5185 (
            .O(N__22378),
            .I(N__22347));
    CascadeMux I__5184 (
            .O(N__22377),
            .I(N__22343));
    CascadeMux I__5183 (
            .O(N__22376),
            .I(N__22340));
    InMux I__5182 (
            .O(N__22375),
            .I(N__22334));
    InMux I__5181 (
            .O(N__22374),
            .I(N__22331));
    CascadeMux I__5180 (
            .O(N__22373),
            .I(N__22328));
    CascadeMux I__5179 (
            .O(N__22372),
            .I(N__22325));
    LocalMux I__5178 (
            .O(N__22369),
            .I(N__22322));
    LocalMux I__5177 (
            .O(N__22366),
            .I(N__22313));
    LocalMux I__5176 (
            .O(N__22363),
            .I(N__22313));
    LocalMux I__5175 (
            .O(N__22360),
            .I(N__22313));
    LocalMux I__5174 (
            .O(N__22357),
            .I(N__22313));
    LocalMux I__5173 (
            .O(N__22354),
            .I(N__22310));
    InMux I__5172 (
            .O(N__22351),
            .I(N__22307));
    InMux I__5171 (
            .O(N__22350),
            .I(N__22302));
    LocalMux I__5170 (
            .O(N__22347),
            .I(N__22299));
    InMux I__5169 (
            .O(N__22346),
            .I(N__22296));
    InMux I__5168 (
            .O(N__22343),
            .I(N__22293));
    InMux I__5167 (
            .O(N__22340),
            .I(N__22290));
    InMux I__5166 (
            .O(N__22339),
            .I(N__22287));
    InMux I__5165 (
            .O(N__22338),
            .I(N__22284));
    InMux I__5164 (
            .O(N__22337),
            .I(N__22281));
    LocalMux I__5163 (
            .O(N__22334),
            .I(N__22276));
    LocalMux I__5162 (
            .O(N__22331),
            .I(N__22276));
    InMux I__5161 (
            .O(N__22328),
            .I(N__22273));
    InMux I__5160 (
            .O(N__22325),
            .I(N__22270));
    Span4Mux_v I__5159 (
            .O(N__22322),
            .I(N__22260));
    Span4Mux_v I__5158 (
            .O(N__22313),
            .I(N__22260));
    Span4Mux_h I__5157 (
            .O(N__22310),
            .I(N__22260));
    LocalMux I__5156 (
            .O(N__22307),
            .I(N__22260));
    InMux I__5155 (
            .O(N__22306),
            .I(N__22257));
    InMux I__5154 (
            .O(N__22305),
            .I(N__22254));
    LocalMux I__5153 (
            .O(N__22302),
            .I(N__22249));
    Span4Mux_v I__5152 (
            .O(N__22299),
            .I(N__22249));
    LocalMux I__5151 (
            .O(N__22296),
            .I(N__22242));
    LocalMux I__5150 (
            .O(N__22293),
            .I(N__22242));
    LocalMux I__5149 (
            .O(N__22290),
            .I(N__22242));
    LocalMux I__5148 (
            .O(N__22287),
            .I(N__22229));
    LocalMux I__5147 (
            .O(N__22284),
            .I(N__22229));
    LocalMux I__5146 (
            .O(N__22281),
            .I(N__22229));
    Span4Mux_v I__5145 (
            .O(N__22276),
            .I(N__22229));
    LocalMux I__5144 (
            .O(N__22273),
            .I(N__22229));
    LocalMux I__5143 (
            .O(N__22270),
            .I(N__22229));
    InMux I__5142 (
            .O(N__22269),
            .I(N__22226));
    Span4Mux_h I__5141 (
            .O(N__22260),
            .I(N__22223));
    LocalMux I__5140 (
            .O(N__22257),
            .I(N__22220));
    LocalMux I__5139 (
            .O(N__22254),
            .I(N__22211));
    Span4Mux_h I__5138 (
            .O(N__22249),
            .I(N__22211));
    Span4Mux_v I__5137 (
            .O(N__22242),
            .I(N__22211));
    Span4Mux_v I__5136 (
            .O(N__22229),
            .I(N__22211));
    LocalMux I__5135 (
            .O(N__22226),
            .I(N__22208));
    Span4Mux_h I__5134 (
            .O(N__22223),
            .I(N__22205));
    Span4Mux_v I__5133 (
            .O(N__22220),
            .I(N__22200));
    Span4Mux_h I__5132 (
            .O(N__22211),
            .I(N__22200));
    Odrv4 I__5131 (
            .O(N__22208),
            .I(TX_ADDR_12));
    Odrv4 I__5130 (
            .O(N__22205),
            .I(TX_ADDR_12));
    Odrv4 I__5129 (
            .O(N__22200),
            .I(TX_ADDR_12));
    InMux I__5128 (
            .O(N__22193),
            .I(N__22190));
    LocalMux I__5127 (
            .O(N__22190),
            .I(N__22187));
    Span4Mux_v I__5126 (
            .O(N__22187),
            .I(N__22184));
    Span4Mux_v I__5125 (
            .O(N__22184),
            .I(N__22181));
    Span4Mux_h I__5124 (
            .O(N__22181),
            .I(N__22178));
    Odrv4 I__5123 (
            .O(N__22178),
            .I(\line_buffer.n593 ));
    InMux I__5122 (
            .O(N__22175),
            .I(N__22172));
    LocalMux I__5121 (
            .O(N__22172),
            .I(\line_buffer.n3596 ));
    IoInMux I__5120 (
            .O(N__22169),
            .I(N__22166));
    LocalMux I__5119 (
            .O(N__22166),
            .I(N__22162));
    InMux I__5118 (
            .O(N__22165),
            .I(N__22159));
    IoSpan4Mux I__5117 (
            .O(N__22162),
            .I(N__22156));
    LocalMux I__5116 (
            .O(N__22159),
            .I(N__22153));
    Span4Mux_s2_h I__5115 (
            .O(N__22156),
            .I(N__22150));
    Span4Mux_v I__5114 (
            .O(N__22153),
            .I(N__22147));
    Sp12to4 I__5113 (
            .O(N__22150),
            .I(N__22144));
    Sp12to4 I__5112 (
            .O(N__22147),
            .I(N__22141));
    Span12Mux_v I__5111 (
            .O(N__22144),
            .I(N__22138));
    Span12Mux_h I__5110 (
            .O(N__22141),
            .I(N__22135));
    Span12Mux_h I__5109 (
            .O(N__22138),
            .I(N__22132));
    Span12Mux_v I__5108 (
            .O(N__22135),
            .I(N__22129));
    Odrv12 I__5107 (
            .O(N__22132),
            .I(DEBUG_c_7_c));
    Odrv12 I__5106 (
            .O(N__22129),
            .I(DEBUG_c_7_c));
    InMux I__5105 (
            .O(N__22124),
            .I(N__22121));
    LocalMux I__5104 (
            .O(N__22121),
            .I(N__22118));
    Span4Mux_v I__5103 (
            .O(N__22118),
            .I(N__22115));
    Span4Mux_h I__5102 (
            .O(N__22115),
            .I(N__22112));
    Odrv4 I__5101 (
            .O(N__22112),
            .I(\line_buffer.n467 ));
    CascadeMux I__5100 (
            .O(N__22109),
            .I(N__22106));
    InMux I__5099 (
            .O(N__22106),
            .I(N__22103));
    LocalMux I__5098 (
            .O(N__22103),
            .I(N__22100));
    Span4Mux_v I__5097 (
            .O(N__22100),
            .I(N__22097));
    Sp12to4 I__5096 (
            .O(N__22097),
            .I(N__22094));
    Span12Mux_h I__5095 (
            .O(N__22094),
            .I(N__22091));
    Span12Mux_v I__5094 (
            .O(N__22091),
            .I(N__22088));
    Odrv12 I__5093 (
            .O(N__22088),
            .I(\line_buffer.n459 ));
    InMux I__5092 (
            .O(N__22085),
            .I(N__22082));
    LocalMux I__5091 (
            .O(N__22082),
            .I(N__22079));
    Odrv4 I__5090 (
            .O(N__22079),
            .I(\line_buffer.n3638 ));
    InMux I__5089 (
            .O(N__22076),
            .I(N__22073));
    LocalMux I__5088 (
            .O(N__22073),
            .I(\line_buffer.n3641 ));
    InMux I__5087 (
            .O(N__22070),
            .I(N__22067));
    LocalMux I__5086 (
            .O(N__22067),
            .I(N__22064));
    Span4Mux_v I__5085 (
            .O(N__22064),
            .I(N__22061));
    Odrv4 I__5084 (
            .O(N__22061),
            .I(TX_DATA_0));
    InMux I__5083 (
            .O(N__22058),
            .I(N__22055));
    LocalMux I__5082 (
            .O(N__22055),
            .I(N__22052));
    Span4Mux_v I__5081 (
            .O(N__22052),
            .I(N__22049));
    Span4Mux_v I__5080 (
            .O(N__22049),
            .I(N__22046));
    Sp12to4 I__5079 (
            .O(N__22046),
            .I(N__22043));
    Span12Mux_h I__5078 (
            .O(N__22043),
            .I(N__22040));
    Span12Mux_v I__5077 (
            .O(N__22040),
            .I(N__22037));
    Odrv12 I__5076 (
            .O(N__22037),
            .I(\line_buffer.n532 ));
    CascadeMux I__5075 (
            .O(N__22034),
            .I(N__22031));
    InMux I__5074 (
            .O(N__22031),
            .I(N__22028));
    LocalMux I__5073 (
            .O(N__22028),
            .I(N__22025));
    Span4Mux_h I__5072 (
            .O(N__22025),
            .I(N__22022));
    Span4Mux_h I__5071 (
            .O(N__22022),
            .I(N__22019));
    Span4Mux_v I__5070 (
            .O(N__22019),
            .I(N__22016));
    Span4Mux_v I__5069 (
            .O(N__22016),
            .I(N__22013));
    Odrv4 I__5068 (
            .O(N__22013),
            .I(\line_buffer.n524 ));
    InMux I__5067 (
            .O(N__22010),
            .I(N__22007));
    LocalMux I__5066 (
            .O(N__22007),
            .I(\line_buffer.n3647 ));
    InMux I__5065 (
            .O(N__22004),
            .I(N__22001));
    LocalMux I__5064 (
            .O(N__22001),
            .I(N__21998));
    Odrv12 I__5063 (
            .O(N__21998),
            .I(TX_DATA_5));
    IoInMux I__5062 (
            .O(N__21995),
            .I(N__21991));
    IoInMux I__5061 (
            .O(N__21994),
            .I(N__21988));
    LocalMux I__5060 (
            .O(N__21991),
            .I(N__21985));
    LocalMux I__5059 (
            .O(N__21988),
            .I(N__21981));
    Span4Mux_s0_v I__5058 (
            .O(N__21985),
            .I(N__21978));
    IoInMux I__5057 (
            .O(N__21984),
            .I(N__21975));
    Span4Mux_s3_v I__5056 (
            .O(N__21981),
            .I(N__21972));
    Sp12to4 I__5055 (
            .O(N__21978),
            .I(N__21969));
    LocalMux I__5054 (
            .O(N__21975),
            .I(N__21966));
    Span4Mux_v I__5053 (
            .O(N__21972),
            .I(N__21963));
    Span12Mux_h I__5052 (
            .O(N__21969),
            .I(N__21960));
    Span12Mux_s6_h I__5051 (
            .O(N__21966),
            .I(N__21955));
    Sp12to4 I__5050 (
            .O(N__21963),
            .I(N__21955));
    Odrv12 I__5049 (
            .O(N__21960),
            .I(n1816));
    Odrv12 I__5048 (
            .O(N__21955),
            .I(n1816));
    InMux I__5047 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__5046 (
            .O(N__21947),
            .I(N__21944));
    Span4Mux_v I__5045 (
            .O(N__21944),
            .I(N__21941));
    Sp12to4 I__5044 (
            .O(N__21941),
            .I(N__21938));
    Span12Mux_v I__5043 (
            .O(N__21938),
            .I(N__21935));
    Odrv12 I__5042 (
            .O(N__21935),
            .I(\line_buffer.n537 ));
    CascadeMux I__5041 (
            .O(N__21932),
            .I(N__21929));
    InMux I__5040 (
            .O(N__21929),
            .I(N__21926));
    LocalMux I__5039 (
            .O(N__21926),
            .I(N__21923));
    Span4Mux_h I__5038 (
            .O(N__21923),
            .I(N__21920));
    Span4Mux_h I__5037 (
            .O(N__21920),
            .I(N__21917));
    Span4Mux_v I__5036 (
            .O(N__21917),
            .I(N__21914));
    Span4Mux_v I__5035 (
            .O(N__21914),
            .I(N__21911));
    Odrv4 I__5034 (
            .O(N__21911),
            .I(\line_buffer.n529 ));
    InMux I__5033 (
            .O(N__21908),
            .I(N__21905));
    LocalMux I__5032 (
            .O(N__21905),
            .I(\line_buffer.n3599 ));
    InMux I__5031 (
            .O(N__21902),
            .I(N__21899));
    LocalMux I__5030 (
            .O(N__21899),
            .I(N__21896));
    Odrv12 I__5029 (
            .O(N__21896),
            .I(\line_buffer.n597 ));
    InMux I__5028 (
            .O(N__21893),
            .I(N__21890));
    LocalMux I__5027 (
            .O(N__21890),
            .I(N__21887));
    Span12Mux_h I__5026 (
            .O(N__21887),
            .I(N__21884));
    Span12Mux_v I__5025 (
            .O(N__21884),
            .I(N__21881));
    Odrv12 I__5024 (
            .O(N__21881),
            .I(\line_buffer.n589 ));
    InMux I__5023 (
            .O(N__21878),
            .I(N__21875));
    LocalMux I__5022 (
            .O(N__21875),
            .I(N__21872));
    Span4Mux_h I__5021 (
            .O(N__21872),
            .I(N__21869));
    Odrv4 I__5020 (
            .O(N__21869),
            .I(\line_buffer.n3650 ));
    InMux I__5019 (
            .O(N__21866),
            .I(N__21863));
    LocalMux I__5018 (
            .O(N__21863),
            .I(N__21860));
    Span4Mux_v I__5017 (
            .O(N__21860),
            .I(N__21857));
    Span4Mux_v I__5016 (
            .O(N__21857),
            .I(N__21854));
    Sp12to4 I__5015 (
            .O(N__21854),
            .I(N__21851));
    Odrv12 I__5014 (
            .O(N__21851),
            .I(\line_buffer.n570 ));
    InMux I__5013 (
            .O(N__21848),
            .I(N__21845));
    LocalMux I__5012 (
            .O(N__21845),
            .I(N__21842));
    Span4Mux_v I__5011 (
            .O(N__21842),
            .I(N__21839));
    Sp12to4 I__5010 (
            .O(N__21839),
            .I(N__21836));
    Span12Mux_h I__5009 (
            .O(N__21836),
            .I(N__21833));
    Span12Mux_v I__5008 (
            .O(N__21833),
            .I(N__21830));
    Odrv12 I__5007 (
            .O(N__21830),
            .I(\line_buffer.n562 ));
    InMux I__5006 (
            .O(N__21827),
            .I(N__21824));
    LocalMux I__5005 (
            .O(N__21824),
            .I(N__21821));
    Odrv12 I__5004 (
            .O(N__21821),
            .I(\line_buffer.n3543 ));
    InMux I__5003 (
            .O(N__21818),
            .I(N__21815));
    LocalMux I__5002 (
            .O(N__21815),
            .I(N__21812));
    Span4Mux_v I__5001 (
            .O(N__21812),
            .I(N__21809));
    Odrv4 I__5000 (
            .O(N__21809),
            .I(\line_buffer.n3656 ));
    InMux I__4999 (
            .O(N__21806),
            .I(N__21803));
    LocalMux I__4998 (
            .O(N__21803),
            .I(N__21800));
    Span4Mux_v I__4997 (
            .O(N__21800),
            .I(N__21797));
    Sp12to4 I__4996 (
            .O(N__21797),
            .I(N__21794));
    Odrv12 I__4995 (
            .O(N__21794),
            .I(\line_buffer.n599 ));
    InMux I__4994 (
            .O(N__21791),
            .I(N__21788));
    LocalMux I__4993 (
            .O(N__21788),
            .I(N__21785));
    Span12Mux_v I__4992 (
            .O(N__21785),
            .I(N__21782));
    Odrv12 I__4991 (
            .O(N__21782),
            .I(\line_buffer.n591 ));
    InMux I__4990 (
            .O(N__21779),
            .I(N__21776));
    LocalMux I__4989 (
            .O(N__21776),
            .I(\line_buffer.n3626 ));
    InMux I__4988 (
            .O(N__21773),
            .I(N__21770));
    LocalMux I__4987 (
            .O(N__21770),
            .I(N__21767));
    Odrv12 I__4986 (
            .O(N__21767),
            .I(TX_DATA_2));
    IoInMux I__4985 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__4984 (
            .O(N__21761),
            .I(N__21757));
    IoInMux I__4983 (
            .O(N__21760),
            .I(N__21754));
    Span4Mux_s3_v I__4982 (
            .O(N__21757),
            .I(N__21751));
    LocalMux I__4981 (
            .O(N__21754),
            .I(N__21748));
    Span4Mux_v I__4980 (
            .O(N__21751),
            .I(N__21744));
    IoSpan4Mux I__4979 (
            .O(N__21748),
            .I(N__21741));
    IoInMux I__4978 (
            .O(N__21747),
            .I(N__21738));
    Span4Mux_v I__4977 (
            .O(N__21744),
            .I(N__21733));
    Span4Mux_s3_h I__4976 (
            .O(N__21741),
            .I(N__21733));
    LocalMux I__4975 (
            .O(N__21738),
            .I(N__21730));
    Span4Mux_h I__4974 (
            .O(N__21733),
            .I(N__21727));
    Span4Mux_s3_v I__4973 (
            .O(N__21730),
            .I(N__21724));
    Span4Mux_h I__4972 (
            .O(N__21727),
            .I(N__21721));
    Span4Mux_v I__4971 (
            .O(N__21724),
            .I(N__21718));
    Span4Mux_h I__4970 (
            .O(N__21721),
            .I(N__21713));
    Span4Mux_v I__4969 (
            .O(N__21718),
            .I(N__21713));
    Odrv4 I__4968 (
            .O(N__21713),
            .I(n1819));
    InMux I__4967 (
            .O(N__21710),
            .I(N__21707));
    LocalMux I__4966 (
            .O(N__21707),
            .I(\line_buffer.n3537 ));
    InMux I__4965 (
            .O(N__21704),
            .I(N__21701));
    LocalMux I__4964 (
            .O(N__21701),
            .I(N__21698));
    Span12Mux_v I__4963 (
            .O(N__21698),
            .I(N__21695));
    Odrv12 I__4962 (
            .O(N__21695),
            .I(\line_buffer.n3536 ));
    InMux I__4961 (
            .O(N__21692),
            .I(N__21689));
    LocalMux I__4960 (
            .O(N__21689),
            .I(\line_buffer.n3614 ));
    InMux I__4959 (
            .O(N__21686),
            .I(N__21683));
    LocalMux I__4958 (
            .O(N__21683),
            .I(N__21680));
    Span12Mux_s10_v I__4957 (
            .O(N__21680),
            .I(N__21677));
    Odrv12 I__4956 (
            .O(N__21677),
            .I(\line_buffer.n469 ));
    InMux I__4955 (
            .O(N__21674),
            .I(N__21671));
    LocalMux I__4954 (
            .O(N__21671),
            .I(N__21668));
    Span4Mux_v I__4953 (
            .O(N__21668),
            .I(N__21665));
    Span4Mux_h I__4952 (
            .O(N__21665),
            .I(N__21662));
    Span4Mux_h I__4951 (
            .O(N__21662),
            .I(N__21659));
    Odrv4 I__4950 (
            .O(N__21659),
            .I(\line_buffer.n461 ));
    InMux I__4949 (
            .O(N__21656),
            .I(N__21653));
    LocalMux I__4948 (
            .O(N__21653),
            .I(N__21650));
    Span12Mux_v I__4947 (
            .O(N__21650),
            .I(N__21647));
    Odrv12 I__4946 (
            .O(N__21647),
            .I(\line_buffer.n3569 ));
    IoInMux I__4945 (
            .O(N__21644),
            .I(N__21641));
    LocalMux I__4944 (
            .O(N__21641),
            .I(N__21638));
    IoSpan4Mux I__4943 (
            .O(N__21638),
            .I(N__21635));
    Span4Mux_s3_h I__4942 (
            .O(N__21635),
            .I(N__21632));
    Span4Mux_h I__4941 (
            .O(N__21632),
            .I(N__21629));
    Span4Mux_h I__4940 (
            .O(N__21629),
            .I(N__21625));
    InMux I__4939 (
            .O(N__21628),
            .I(N__21622));
    Span4Mux_h I__4938 (
            .O(N__21625),
            .I(N__21617));
    LocalMux I__4937 (
            .O(N__21622),
            .I(N__21617));
    Span4Mux_h I__4936 (
            .O(N__21617),
            .I(N__21614));
    Sp12to4 I__4935 (
            .O(N__21614),
            .I(N__21611));
    Odrv12 I__4934 (
            .O(N__21611),
            .I(DEBUG_c_2_c));
    InMux I__4933 (
            .O(N__21608),
            .I(N__21605));
    LocalMux I__4932 (
            .O(N__21605),
            .I(\tvp_hs_buffer.BUFFER_0_0 ));
    InMux I__4931 (
            .O(N__21602),
            .I(N__21599));
    LocalMux I__4930 (
            .O(N__21599),
            .I(N__21596));
    Span4Mux_v I__4929 (
            .O(N__21596),
            .I(N__21593));
    Sp12to4 I__4928 (
            .O(N__21593),
            .I(N__21590));
    Odrv12 I__4927 (
            .O(N__21590),
            .I(\line_buffer.n598 ));
    InMux I__4926 (
            .O(N__21587),
            .I(N__21584));
    LocalMux I__4925 (
            .O(N__21584),
            .I(N__21581));
    Span4Mux_v I__4924 (
            .O(N__21581),
            .I(N__21578));
    Sp12to4 I__4923 (
            .O(N__21578),
            .I(N__21575));
    Span12Mux_h I__4922 (
            .O(N__21575),
            .I(N__21572));
    Span12Mux_v I__4921 (
            .O(N__21572),
            .I(N__21569));
    Odrv12 I__4920 (
            .O(N__21569),
            .I(\line_buffer.n590 ));
    InMux I__4919 (
            .O(N__21566),
            .I(N__21563));
    LocalMux I__4918 (
            .O(N__21563),
            .I(\line_buffer.n3573 ));
    InMux I__4917 (
            .O(N__21560),
            .I(N__21557));
    LocalMux I__4916 (
            .O(N__21557),
            .I(\line_buffer.n3659 ));
    InMux I__4915 (
            .O(N__21554),
            .I(N__21551));
    LocalMux I__4914 (
            .O(N__21551),
            .I(N__21548));
    Span4Mux_v I__4913 (
            .O(N__21548),
            .I(N__21545));
    Span4Mux_v I__4912 (
            .O(N__21545),
            .I(N__21542));
    Sp12to4 I__4911 (
            .O(N__21542),
            .I(N__21539));
    Odrv12 I__4910 (
            .O(N__21539),
            .I(\line_buffer.n564 ));
    InMux I__4909 (
            .O(N__21536),
            .I(N__21533));
    LocalMux I__4908 (
            .O(N__21533),
            .I(N__21530));
    Span4Mux_v I__4907 (
            .O(N__21530),
            .I(N__21527));
    Span4Mux_h I__4906 (
            .O(N__21527),
            .I(N__21524));
    Odrv4 I__4905 (
            .O(N__21524),
            .I(\line_buffer.n556 ));
    InMux I__4904 (
            .O(N__21521),
            .I(N__21518));
    LocalMux I__4903 (
            .O(N__21518),
            .I(N__21515));
    Span4Mux_v I__4902 (
            .O(N__21515),
            .I(N__21512));
    Span4Mux_h I__4901 (
            .O(N__21512),
            .I(N__21509));
    Span4Mux_h I__4900 (
            .O(N__21509),
            .I(N__21506));
    Odrv4 I__4899 (
            .O(N__21506),
            .I(\line_buffer.n534 ));
    InMux I__4898 (
            .O(N__21503),
            .I(N__21500));
    LocalMux I__4897 (
            .O(N__21500),
            .I(N__21497));
    Odrv12 I__4896 (
            .O(N__21497),
            .I(\line_buffer.n526 ));
    InMux I__4895 (
            .O(N__21494),
            .I(N__21491));
    LocalMux I__4894 (
            .O(N__21491),
            .I(N__21488));
    Odrv4 I__4893 (
            .O(N__21488),
            .I(\transmit_module.X_DELTA_PATTERN_6 ));
    InMux I__4892 (
            .O(N__21485),
            .I(N__21482));
    LocalMux I__4891 (
            .O(N__21482),
            .I(N__21479));
    Odrv4 I__4890 (
            .O(N__21479),
            .I(\transmit_module.X_DELTA_PATTERN_5 ));
    CEMux I__4889 (
            .O(N__21476),
            .I(N__21471));
    CEMux I__4888 (
            .O(N__21475),
            .I(N__21468));
    CEMux I__4887 (
            .O(N__21474),
            .I(N__21465));
    LocalMux I__4886 (
            .O(N__21471),
            .I(N__21461));
    LocalMux I__4885 (
            .O(N__21468),
            .I(N__21458));
    LocalMux I__4884 (
            .O(N__21465),
            .I(N__21455));
    CEMux I__4883 (
            .O(N__21464),
            .I(N__21452));
    Span4Mux_v I__4882 (
            .O(N__21461),
            .I(N__21449));
    Span4Mux_h I__4881 (
            .O(N__21458),
            .I(N__21446));
    Span4Mux_h I__4880 (
            .O(N__21455),
            .I(N__21443));
    LocalMux I__4879 (
            .O(N__21452),
            .I(N__21440));
    Odrv4 I__4878 (
            .O(N__21449),
            .I(\transmit_module.n2087 ));
    Odrv4 I__4877 (
            .O(N__21446),
            .I(\transmit_module.n2087 ));
    Odrv4 I__4876 (
            .O(N__21443),
            .I(\transmit_module.n2087 ));
    Odrv12 I__4875 (
            .O(N__21440),
            .I(\transmit_module.n2087 ));
    CEMux I__4874 (
            .O(N__21431),
            .I(N__21423));
    CEMux I__4873 (
            .O(N__21430),
            .I(N__21420));
    CEMux I__4872 (
            .O(N__21429),
            .I(N__21417));
    CEMux I__4871 (
            .O(N__21428),
            .I(N__21414));
    CEMux I__4870 (
            .O(N__21427),
            .I(N__21411));
    CEMux I__4869 (
            .O(N__21426),
            .I(N__21408));
    LocalMux I__4868 (
            .O(N__21423),
            .I(N__21402));
    LocalMux I__4867 (
            .O(N__21420),
            .I(N__21399));
    LocalMux I__4866 (
            .O(N__21417),
            .I(N__21392));
    LocalMux I__4865 (
            .O(N__21414),
            .I(N__21392));
    LocalMux I__4864 (
            .O(N__21411),
            .I(N__21392));
    LocalMux I__4863 (
            .O(N__21408),
            .I(N__21389));
    CEMux I__4862 (
            .O(N__21407),
            .I(N__21386));
    CEMux I__4861 (
            .O(N__21406),
            .I(N__21383));
    CEMux I__4860 (
            .O(N__21405),
            .I(N__21378));
    Span4Mux_v I__4859 (
            .O(N__21402),
            .I(N__21373));
    Span4Mux_v I__4858 (
            .O(N__21399),
            .I(N__21373));
    Span4Mux_v I__4857 (
            .O(N__21392),
            .I(N__21366));
    Span4Mux_h I__4856 (
            .O(N__21389),
            .I(N__21366));
    LocalMux I__4855 (
            .O(N__21386),
            .I(N__21366));
    LocalMux I__4854 (
            .O(N__21383),
            .I(N__21363));
    CEMux I__4853 (
            .O(N__21382),
            .I(N__21359));
    CEMux I__4852 (
            .O(N__21381),
            .I(N__21356));
    LocalMux I__4851 (
            .O(N__21378),
            .I(N__21351));
    Span4Mux_h I__4850 (
            .O(N__21373),
            .I(N__21344));
    Span4Mux_h I__4849 (
            .O(N__21366),
            .I(N__21344));
    Span4Mux_v I__4848 (
            .O(N__21363),
            .I(N__21344));
    SRMux I__4847 (
            .O(N__21362),
            .I(N__21341));
    LocalMux I__4846 (
            .O(N__21359),
            .I(N__21338));
    LocalMux I__4845 (
            .O(N__21356),
            .I(N__21335));
    SRMux I__4844 (
            .O(N__21355),
            .I(N__21332));
    SRMux I__4843 (
            .O(N__21354),
            .I(N__21328));
    Span4Mux_v I__4842 (
            .O(N__21351),
            .I(N__21322));
    Span4Mux_h I__4841 (
            .O(N__21344),
            .I(N__21322));
    LocalMux I__4840 (
            .O(N__21341),
            .I(N__21319));
    Span4Mux_h I__4839 (
            .O(N__21338),
            .I(N__21312));
    Span4Mux_v I__4838 (
            .O(N__21335),
            .I(N__21312));
    LocalMux I__4837 (
            .O(N__21332),
            .I(N__21312));
    CEMux I__4836 (
            .O(N__21331),
            .I(N__21309));
    LocalMux I__4835 (
            .O(N__21328),
            .I(N__21306));
    SRMux I__4834 (
            .O(N__21327),
            .I(N__21303));
    Span4Mux_h I__4833 (
            .O(N__21322),
            .I(N__21300));
    Span4Mux_h I__4832 (
            .O(N__21319),
            .I(N__21297));
    Span4Mux_h I__4831 (
            .O(N__21312),
            .I(N__21294));
    LocalMux I__4830 (
            .O(N__21309),
            .I(N__21287));
    Sp12to4 I__4829 (
            .O(N__21306),
            .I(N__21287));
    LocalMux I__4828 (
            .O(N__21303),
            .I(N__21287));
    Odrv4 I__4827 (
            .O(N__21300),
            .I(\transmit_module.n3682 ));
    Odrv4 I__4826 (
            .O(N__21297),
            .I(\transmit_module.n3682 ));
    Odrv4 I__4825 (
            .O(N__21294),
            .I(\transmit_module.n3682 ));
    Odrv12 I__4824 (
            .O(N__21287),
            .I(\transmit_module.n3682 ));
    InMux I__4823 (
            .O(N__21278),
            .I(N__21275));
    LocalMux I__4822 (
            .O(N__21275),
            .I(N__21272));
    Span4Mux_h I__4821 (
            .O(N__21272),
            .I(N__21269));
    Sp12to4 I__4820 (
            .O(N__21269),
            .I(N__21266));
    Span12Mux_v I__4819 (
            .O(N__21266),
            .I(N__21263));
    Odrv12 I__4818 (
            .O(N__21263),
            .I(\line_buffer.n533 ));
    CascadeMux I__4817 (
            .O(N__21260),
            .I(N__21257));
    InMux I__4816 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__4815 (
            .O(N__21254),
            .I(N__21251));
    Span4Mux_v I__4814 (
            .O(N__21251),
            .I(N__21248));
    Span4Mux_h I__4813 (
            .O(N__21248),
            .I(N__21245));
    Odrv4 I__4812 (
            .O(N__21245),
            .I(\line_buffer.n525 ));
    InMux I__4811 (
            .O(N__21242),
            .I(N__21239));
    LocalMux I__4810 (
            .O(N__21239),
            .I(\line_buffer.n3653 ));
    InMux I__4809 (
            .O(N__21236),
            .I(N__21233));
    LocalMux I__4808 (
            .O(N__21233),
            .I(N__21230));
    Span12Mux_v I__4807 (
            .O(N__21230),
            .I(N__21227));
    Odrv12 I__4806 (
            .O(N__21227),
            .I(\line_buffer.n468 ));
    CascadeMux I__4805 (
            .O(N__21224),
            .I(N__21221));
    InMux I__4804 (
            .O(N__21221),
            .I(N__21218));
    LocalMux I__4803 (
            .O(N__21218),
            .I(N__21215));
    Span12Mux_v I__4802 (
            .O(N__21215),
            .I(N__21212));
    Odrv12 I__4801 (
            .O(N__21212),
            .I(\line_buffer.n460 ));
    InMux I__4800 (
            .O(N__21209),
            .I(N__21206));
    LocalMux I__4799 (
            .O(N__21206),
            .I(\line_buffer.n3635 ));
    InMux I__4798 (
            .O(N__21203),
            .I(N__21200));
    LocalMux I__4797 (
            .O(N__21200),
            .I(N__21197));
    Span4Mux_v I__4796 (
            .O(N__21197),
            .I(N__21194));
    Span4Mux_h I__4795 (
            .O(N__21194),
            .I(N__21191));
    Span4Mux_h I__4794 (
            .O(N__21191),
            .I(N__21188));
    Odrv4 I__4793 (
            .O(N__21188),
            .I(\line_buffer.n566 ));
    InMux I__4792 (
            .O(N__21185),
            .I(N__21182));
    LocalMux I__4791 (
            .O(N__21182),
            .I(N__21179));
    Odrv12 I__4790 (
            .O(N__21179),
            .I(\line_buffer.n558 ));
    InMux I__4789 (
            .O(N__21176),
            .I(N__21173));
    LocalMux I__4788 (
            .O(N__21173),
            .I(N__21170));
    Odrv12 I__4787 (
            .O(N__21170),
            .I(\line_buffer.n557 ));
    InMux I__4786 (
            .O(N__21167),
            .I(N__21164));
    LocalMux I__4785 (
            .O(N__21164),
            .I(N__21161));
    Span4Mux_v I__4784 (
            .O(N__21161),
            .I(N__21158));
    Span4Mux_h I__4783 (
            .O(N__21158),
            .I(N__21155));
    Span4Mux_h I__4782 (
            .O(N__21155),
            .I(N__21152));
    Odrv4 I__4781 (
            .O(N__21152),
            .I(\line_buffer.n565 ));
    InMux I__4780 (
            .O(N__21149),
            .I(N__21146));
    LocalMux I__4779 (
            .O(N__21146),
            .I(\line_buffer.n3632 ));
    InMux I__4778 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__4777 (
            .O(N__21140),
            .I(N__21137));
    Span4Mux_v I__4776 (
            .O(N__21137),
            .I(N__21134));
    Odrv4 I__4775 (
            .O(N__21134),
            .I(\line_buffer.n3572 ));
    CascadeMux I__4774 (
            .O(N__21131),
            .I(\line_buffer.n3602_cascade_ ));
    InMux I__4773 (
            .O(N__21128),
            .I(N__21125));
    LocalMux I__4772 (
            .O(N__21125),
            .I(\line_buffer.n3570 ));
    InMux I__4771 (
            .O(N__21122),
            .I(N__21119));
    LocalMux I__4770 (
            .O(N__21119),
            .I(N__21116));
    Span4Mux_h I__4769 (
            .O(N__21116),
            .I(N__21113));
    Span4Mux_h I__4768 (
            .O(N__21113),
            .I(N__21110));
    Odrv4 I__4767 (
            .O(N__21110),
            .I(\line_buffer.n472 ));
    CascadeMux I__4766 (
            .O(N__21107),
            .I(N__21104));
    InMux I__4765 (
            .O(N__21104),
            .I(N__21101));
    LocalMux I__4764 (
            .O(N__21101),
            .I(N__21098));
    Span4Mux_v I__4763 (
            .O(N__21098),
            .I(N__21095));
    Sp12to4 I__4762 (
            .O(N__21095),
            .I(N__21092));
    Span12Mux_h I__4761 (
            .O(N__21092),
            .I(N__21089));
    Odrv12 I__4760 (
            .O(N__21089),
            .I(\line_buffer.n464 ));
    CascadeMux I__4759 (
            .O(N__21086),
            .I(\line_buffer.n3593_cascade_ ));
    InMux I__4758 (
            .O(N__21083),
            .I(N__21080));
    LocalMux I__4757 (
            .O(N__21080),
            .I(N__21077));
    Odrv4 I__4756 (
            .O(N__21077),
            .I(\line_buffer.n3629 ));
    InMux I__4755 (
            .O(N__21074),
            .I(N__21071));
    LocalMux I__4754 (
            .O(N__21071),
            .I(TX_DATA_3));
    InMux I__4753 (
            .O(N__21068),
            .I(N__21065));
    LocalMux I__4752 (
            .O(N__21065),
            .I(N__21062));
    Span4Mux_v I__4751 (
            .O(N__21062),
            .I(N__21059));
    Sp12to4 I__4750 (
            .O(N__21059),
            .I(N__21056));
    Odrv12 I__4749 (
            .O(N__21056),
            .I(\line_buffer.n471 ));
    InMux I__4748 (
            .O(N__21053),
            .I(N__21050));
    LocalMux I__4747 (
            .O(N__21050),
            .I(N__21047));
    Span4Mux_h I__4746 (
            .O(N__21047),
            .I(N__21044));
    Span4Mux_v I__4745 (
            .O(N__21044),
            .I(N__21041));
    Span4Mux_h I__4744 (
            .O(N__21041),
            .I(N__21038));
    Odrv4 I__4743 (
            .O(N__21038),
            .I(\line_buffer.n463 ));
    InMux I__4742 (
            .O(N__21035),
            .I(N__21032));
    LocalMux I__4741 (
            .O(N__21032),
            .I(N__21029));
    Span4Mux_v I__4740 (
            .O(N__21029),
            .I(N__21026));
    Span4Mux_v I__4739 (
            .O(N__21026),
            .I(N__21023));
    Odrv4 I__4738 (
            .O(N__21023),
            .I(\line_buffer.n3552 ));
    CascadeMux I__4737 (
            .O(N__21020),
            .I(\line_buffer.n3551_cascade_ ));
    InMux I__4736 (
            .O(N__21017),
            .I(N__21014));
    LocalMux I__4735 (
            .O(N__21014),
            .I(N__21011));
    Span4Mux_v I__4734 (
            .O(N__21011),
            .I(N__21008));
    Span4Mux_h I__4733 (
            .O(N__21008),
            .I(N__21005));
    Span4Mux_h I__4732 (
            .O(N__21005),
            .I(N__21002));
    Span4Mux_v I__4731 (
            .O(N__21002),
            .I(N__20999));
    Odrv4 I__4730 (
            .O(N__20999),
            .I(\line_buffer.n600 ));
    InMux I__4729 (
            .O(N__20996),
            .I(N__20993));
    LocalMux I__4728 (
            .O(N__20993),
            .I(N__20990));
    Span4Mux_v I__4727 (
            .O(N__20990),
            .I(N__20987));
    Span4Mux_h I__4726 (
            .O(N__20987),
            .I(N__20984));
    Span4Mux_h I__4725 (
            .O(N__20984),
            .I(N__20981));
    Odrv4 I__4724 (
            .O(N__20981),
            .I(\line_buffer.n592 ));
    InMux I__4723 (
            .O(N__20978),
            .I(N__20975));
    LocalMux I__4722 (
            .O(N__20975),
            .I(N__20972));
    Odrv4 I__4721 (
            .O(N__20972),
            .I(TX_DATA_4));
    IoInMux I__4720 (
            .O(N__20969),
            .I(N__20966));
    LocalMux I__4719 (
            .O(N__20966),
            .I(N__20961));
    IoInMux I__4718 (
            .O(N__20965),
            .I(N__20958));
    IoInMux I__4717 (
            .O(N__20964),
            .I(N__20955));
    IoSpan4Mux I__4716 (
            .O(N__20961),
            .I(N__20952));
    LocalMux I__4715 (
            .O(N__20958),
            .I(N__20949));
    LocalMux I__4714 (
            .O(N__20955),
            .I(N__20946));
    Span4Mux_s0_v I__4713 (
            .O(N__20952),
            .I(N__20943));
    IoSpan4Mux I__4712 (
            .O(N__20949),
            .I(N__20940));
    IoSpan4Mux I__4711 (
            .O(N__20946),
            .I(N__20937));
    Span4Mux_v I__4710 (
            .O(N__20943),
            .I(N__20934));
    Span4Mux_s3_h I__4709 (
            .O(N__20940),
            .I(N__20931));
    Span4Mux_s2_v I__4708 (
            .O(N__20937),
            .I(N__20928));
    Span4Mux_v I__4707 (
            .O(N__20934),
            .I(N__20923));
    Span4Mux_h I__4706 (
            .O(N__20931),
            .I(N__20923));
    Sp12to4 I__4705 (
            .O(N__20928),
            .I(N__20920));
    Span4Mux_h I__4704 (
            .O(N__20923),
            .I(N__20917));
    Span12Mux_s8_v I__4703 (
            .O(N__20920),
            .I(N__20914));
    Span4Mux_h I__4702 (
            .O(N__20917),
            .I(N__20911));
    Odrv12 I__4701 (
            .O(N__20914),
            .I(n1817));
    Odrv4 I__4700 (
            .O(N__20911),
            .I(n1817));
    InMux I__4699 (
            .O(N__20906),
            .I(N__20903));
    LocalMux I__4698 (
            .O(N__20903),
            .I(N__20900));
    Span12Mux_s10_v I__4697 (
            .O(N__20900),
            .I(N__20897));
    Odrv12 I__4696 (
            .O(N__20897),
            .I(TX_DATA_1));
    IoInMux I__4695 (
            .O(N__20894),
            .I(N__20891));
    LocalMux I__4694 (
            .O(N__20891),
            .I(N__20887));
    IoInMux I__4693 (
            .O(N__20890),
            .I(N__20884));
    IoSpan4Mux I__4692 (
            .O(N__20887),
            .I(N__20879));
    LocalMux I__4691 (
            .O(N__20884),
            .I(N__20879));
    IoSpan4Mux I__4690 (
            .O(N__20879),
            .I(N__20876));
    Span4Mux_s2_h I__4689 (
            .O(N__20876),
            .I(N__20872));
    IoInMux I__4688 (
            .O(N__20875),
            .I(N__20869));
    Span4Mux_h I__4687 (
            .O(N__20872),
            .I(N__20866));
    LocalMux I__4686 (
            .O(N__20869),
            .I(N__20863));
    Span4Mux_h I__4685 (
            .O(N__20866),
            .I(N__20860));
    Span4Mux_s3_v I__4684 (
            .O(N__20863),
            .I(N__20857));
    Span4Mux_h I__4683 (
            .O(N__20860),
            .I(N__20852));
    Span4Mux_v I__4682 (
            .O(N__20857),
            .I(N__20852));
    Odrv4 I__4681 (
            .O(N__20852),
            .I(n1820));
    InMux I__4680 (
            .O(N__20849),
            .I(N__20846));
    LocalMux I__4679 (
            .O(N__20846),
            .I(N__20843));
    Odrv4 I__4678 (
            .O(N__20843),
            .I(\tvp_hs_buffer.BUFFER_1_0 ));
    InMux I__4677 (
            .O(N__20840),
            .I(N__20837));
    LocalMux I__4676 (
            .O(N__20837),
            .I(N__20834));
    Span4Mux_v I__4675 (
            .O(N__20834),
            .I(N__20831));
    Span4Mux_h I__4674 (
            .O(N__20831),
            .I(N__20828));
    Span4Mux_h I__4673 (
            .O(N__20828),
            .I(N__20825));
    Odrv4 I__4672 (
            .O(N__20825),
            .I(\line_buffer.n536 ));
    InMux I__4671 (
            .O(N__20822),
            .I(N__20819));
    LocalMux I__4670 (
            .O(N__20819),
            .I(N__20816));
    Span12Mux_v I__4669 (
            .O(N__20816),
            .I(N__20813));
    Odrv12 I__4668 (
            .O(N__20813),
            .I(\line_buffer.n528 ));
    InMux I__4667 (
            .O(N__20810),
            .I(N__20807));
    LocalMux I__4666 (
            .O(N__20807),
            .I(N__20801));
    InMux I__4665 (
            .O(N__20806),
            .I(N__20798));
    InMux I__4664 (
            .O(N__20805),
            .I(N__20795));
    InMux I__4663 (
            .O(N__20804),
            .I(N__20792));
    Odrv12 I__4662 (
            .O(N__20801),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__4661 (
            .O(N__20798),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__4660 (
            .O(N__20795),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__4659 (
            .O(N__20792),
            .I(\transmit_module.TX_ADDR_4 ));
    InMux I__4658 (
            .O(N__20783),
            .I(N__20780));
    LocalMux I__4657 (
            .O(N__20780),
            .I(N__20777));
    Odrv4 I__4656 (
            .O(N__20777),
            .I(\transmit_module.ADDR_Y_COMPONENT_4 ));
    CEMux I__4655 (
            .O(N__20774),
            .I(N__20768));
    CEMux I__4654 (
            .O(N__20773),
            .I(N__20765));
    CEMux I__4653 (
            .O(N__20772),
            .I(N__20761));
    CEMux I__4652 (
            .O(N__20771),
            .I(N__20758));
    LocalMux I__4651 (
            .O(N__20768),
            .I(N__20752));
    LocalMux I__4650 (
            .O(N__20765),
            .I(N__20752));
    CEMux I__4649 (
            .O(N__20764),
            .I(N__20749));
    LocalMux I__4648 (
            .O(N__20761),
            .I(N__20745));
    LocalMux I__4647 (
            .O(N__20758),
            .I(N__20742));
    CEMux I__4646 (
            .O(N__20757),
            .I(N__20739));
    Span4Mux_h I__4645 (
            .O(N__20752),
            .I(N__20735));
    LocalMux I__4644 (
            .O(N__20749),
            .I(N__20732));
    CEMux I__4643 (
            .O(N__20748),
            .I(N__20729));
    Span4Mux_v I__4642 (
            .O(N__20745),
            .I(N__20724));
    Span4Mux_h I__4641 (
            .O(N__20742),
            .I(N__20724));
    LocalMux I__4640 (
            .O(N__20739),
            .I(N__20721));
    CEMux I__4639 (
            .O(N__20738),
            .I(N__20718));
    Span4Mux_v I__4638 (
            .O(N__20735),
            .I(N__20713));
    Span4Mux_h I__4637 (
            .O(N__20732),
            .I(N__20713));
    LocalMux I__4636 (
            .O(N__20729),
            .I(N__20710));
    Span4Mux_h I__4635 (
            .O(N__20724),
            .I(N__20707));
    Span4Mux_h I__4634 (
            .O(N__20721),
            .I(N__20704));
    LocalMux I__4633 (
            .O(N__20718),
            .I(N__20701));
    Odrv4 I__4632 (
            .O(N__20713),
            .I(\transmit_module.n2313 ));
    Odrv12 I__4631 (
            .O(N__20710),
            .I(\transmit_module.n2313 ));
    Odrv4 I__4630 (
            .O(N__20707),
            .I(\transmit_module.n2313 ));
    Odrv4 I__4629 (
            .O(N__20704),
            .I(\transmit_module.n2313 ));
    Odrv4 I__4628 (
            .O(N__20701),
            .I(\transmit_module.n2313 ));
    InMux I__4627 (
            .O(N__20690),
            .I(N__20687));
    LocalMux I__4626 (
            .O(N__20687),
            .I(\transmit_module.ADDR_Y_COMPONENT_2 ));
    InMux I__4625 (
            .O(N__20684),
            .I(N__20679));
    InMux I__4624 (
            .O(N__20683),
            .I(N__20673));
    InMux I__4623 (
            .O(N__20682),
            .I(N__20668));
    LocalMux I__4622 (
            .O(N__20679),
            .I(N__20665));
    InMux I__4621 (
            .O(N__20678),
            .I(N__20662));
    InMux I__4620 (
            .O(N__20677),
            .I(N__20656));
    InMux I__4619 (
            .O(N__20676),
            .I(N__20656));
    LocalMux I__4618 (
            .O(N__20673),
            .I(N__20652));
    InMux I__4617 (
            .O(N__20672),
            .I(N__20649));
    InMux I__4616 (
            .O(N__20671),
            .I(N__20644));
    LocalMux I__4615 (
            .O(N__20668),
            .I(N__20641));
    Span4Mux_h I__4614 (
            .O(N__20665),
            .I(N__20636));
    LocalMux I__4613 (
            .O(N__20662),
            .I(N__20636));
    InMux I__4612 (
            .O(N__20661),
            .I(N__20633));
    LocalMux I__4611 (
            .O(N__20656),
            .I(N__20630));
    InMux I__4610 (
            .O(N__20655),
            .I(N__20627));
    Span4Mux_h I__4609 (
            .O(N__20652),
            .I(N__20620));
    LocalMux I__4608 (
            .O(N__20649),
            .I(N__20620));
    InMux I__4607 (
            .O(N__20648),
            .I(N__20615));
    InMux I__4606 (
            .O(N__20647),
            .I(N__20615));
    LocalMux I__4605 (
            .O(N__20644),
            .I(N__20612));
    Span4Mux_v I__4604 (
            .O(N__20641),
            .I(N__20605));
    Span4Mux_v I__4603 (
            .O(N__20636),
            .I(N__20605));
    LocalMux I__4602 (
            .O(N__20633),
            .I(N__20605));
    Span4Mux_v I__4601 (
            .O(N__20630),
            .I(N__20600));
    LocalMux I__4600 (
            .O(N__20627),
            .I(N__20600));
    InMux I__4599 (
            .O(N__20626),
            .I(N__20597));
    InMux I__4598 (
            .O(N__20625),
            .I(N__20594));
    Odrv4 I__4597 (
            .O(N__20620),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4596 (
            .O(N__20615),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4595 (
            .O(N__20612),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4594 (
            .O(N__20605),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4593 (
            .O(N__20600),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4592 (
            .O(N__20597),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4591 (
            .O(N__20594),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    InMux I__4590 (
            .O(N__20579),
            .I(N__20574));
    InMux I__4589 (
            .O(N__20578),
            .I(N__20570));
    InMux I__4588 (
            .O(N__20577),
            .I(N__20567));
    LocalMux I__4587 (
            .O(N__20574),
            .I(N__20564));
    InMux I__4586 (
            .O(N__20573),
            .I(N__20561));
    LocalMux I__4585 (
            .O(N__20570),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__4584 (
            .O(N__20567),
            .I(\transmit_module.TX_ADDR_2 ));
    Odrv4 I__4583 (
            .O(N__20564),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__4582 (
            .O(N__20561),
            .I(\transmit_module.TX_ADDR_2 ));
    InMux I__4581 (
            .O(N__20552),
            .I(N__20549));
    LocalMux I__4580 (
            .O(N__20549),
            .I(N__20545));
    InMux I__4579 (
            .O(N__20548),
            .I(N__20542));
    Odrv4 I__4578 (
            .O(N__20545),
            .I(\transmit_module.n114 ));
    LocalMux I__4577 (
            .O(N__20542),
            .I(\transmit_module.n114 ));
    InMux I__4576 (
            .O(N__20537),
            .I(N__20534));
    LocalMux I__4575 (
            .O(N__20534),
            .I(N__20531));
    Odrv4 I__4574 (
            .O(N__20531),
            .I(\transmit_module.n145 ));
    CascadeMux I__4573 (
            .O(N__20528),
            .I(N__20524));
    CascadeMux I__4572 (
            .O(N__20527),
            .I(N__20521));
    CascadeBuf I__4571 (
            .O(N__20524),
            .I(N__20518));
    CascadeBuf I__4570 (
            .O(N__20521),
            .I(N__20515));
    CascadeMux I__4569 (
            .O(N__20518),
            .I(N__20512));
    CascadeMux I__4568 (
            .O(N__20515),
            .I(N__20509));
    CascadeBuf I__4567 (
            .O(N__20512),
            .I(N__20506));
    CascadeBuf I__4566 (
            .O(N__20509),
            .I(N__20503));
    CascadeMux I__4565 (
            .O(N__20506),
            .I(N__20500));
    CascadeMux I__4564 (
            .O(N__20503),
            .I(N__20497));
    CascadeBuf I__4563 (
            .O(N__20500),
            .I(N__20494));
    CascadeBuf I__4562 (
            .O(N__20497),
            .I(N__20491));
    CascadeMux I__4561 (
            .O(N__20494),
            .I(N__20488));
    CascadeMux I__4560 (
            .O(N__20491),
            .I(N__20485));
    CascadeBuf I__4559 (
            .O(N__20488),
            .I(N__20482));
    CascadeBuf I__4558 (
            .O(N__20485),
            .I(N__20479));
    CascadeMux I__4557 (
            .O(N__20482),
            .I(N__20476));
    CascadeMux I__4556 (
            .O(N__20479),
            .I(N__20473));
    CascadeBuf I__4555 (
            .O(N__20476),
            .I(N__20470));
    CascadeBuf I__4554 (
            .O(N__20473),
            .I(N__20467));
    CascadeMux I__4553 (
            .O(N__20470),
            .I(N__20464));
    CascadeMux I__4552 (
            .O(N__20467),
            .I(N__20461));
    CascadeBuf I__4551 (
            .O(N__20464),
            .I(N__20458));
    CascadeBuf I__4550 (
            .O(N__20461),
            .I(N__20455));
    CascadeMux I__4549 (
            .O(N__20458),
            .I(N__20452));
    CascadeMux I__4548 (
            .O(N__20455),
            .I(N__20449));
    CascadeBuf I__4547 (
            .O(N__20452),
            .I(N__20446));
    CascadeBuf I__4546 (
            .O(N__20449),
            .I(N__20443));
    CascadeMux I__4545 (
            .O(N__20446),
            .I(N__20440));
    CascadeMux I__4544 (
            .O(N__20443),
            .I(N__20437));
    CascadeBuf I__4543 (
            .O(N__20440),
            .I(N__20434));
    CascadeBuf I__4542 (
            .O(N__20437),
            .I(N__20431));
    CascadeMux I__4541 (
            .O(N__20434),
            .I(N__20428));
    CascadeMux I__4540 (
            .O(N__20431),
            .I(N__20425));
    CascadeBuf I__4539 (
            .O(N__20428),
            .I(N__20422));
    CascadeBuf I__4538 (
            .O(N__20425),
            .I(N__20419));
    CascadeMux I__4537 (
            .O(N__20422),
            .I(N__20416));
    CascadeMux I__4536 (
            .O(N__20419),
            .I(N__20413));
    CascadeBuf I__4535 (
            .O(N__20416),
            .I(N__20410));
    CascadeBuf I__4534 (
            .O(N__20413),
            .I(N__20407));
    CascadeMux I__4533 (
            .O(N__20410),
            .I(N__20404));
    CascadeMux I__4532 (
            .O(N__20407),
            .I(N__20401));
    CascadeBuf I__4531 (
            .O(N__20404),
            .I(N__20398));
    CascadeBuf I__4530 (
            .O(N__20401),
            .I(N__20395));
    CascadeMux I__4529 (
            .O(N__20398),
            .I(N__20392));
    CascadeMux I__4528 (
            .O(N__20395),
            .I(N__20389));
    CascadeBuf I__4527 (
            .O(N__20392),
            .I(N__20386));
    CascadeBuf I__4526 (
            .O(N__20389),
            .I(N__20383));
    CascadeMux I__4525 (
            .O(N__20386),
            .I(N__20380));
    CascadeMux I__4524 (
            .O(N__20383),
            .I(N__20377));
    CascadeBuf I__4523 (
            .O(N__20380),
            .I(N__20374));
    CascadeBuf I__4522 (
            .O(N__20377),
            .I(N__20371));
    CascadeMux I__4521 (
            .O(N__20374),
            .I(N__20368));
    CascadeMux I__4520 (
            .O(N__20371),
            .I(N__20365));
    CascadeBuf I__4519 (
            .O(N__20368),
            .I(N__20362));
    CascadeBuf I__4518 (
            .O(N__20365),
            .I(N__20359));
    CascadeMux I__4517 (
            .O(N__20362),
            .I(N__20356));
    CascadeMux I__4516 (
            .O(N__20359),
            .I(N__20353));
    CascadeBuf I__4515 (
            .O(N__20356),
            .I(N__20350));
    CascadeBuf I__4514 (
            .O(N__20353),
            .I(N__20347));
    CascadeMux I__4513 (
            .O(N__20350),
            .I(N__20344));
    CascadeMux I__4512 (
            .O(N__20347),
            .I(N__20341));
    InMux I__4511 (
            .O(N__20344),
            .I(N__20338));
    InMux I__4510 (
            .O(N__20341),
            .I(N__20335));
    LocalMux I__4509 (
            .O(N__20338),
            .I(N__20332));
    LocalMux I__4508 (
            .O(N__20335),
            .I(N__20329));
    Span4Mux_h I__4507 (
            .O(N__20332),
            .I(N__20326));
    Span4Mux_v I__4506 (
            .O(N__20329),
            .I(N__20323));
    Span4Mux_h I__4505 (
            .O(N__20326),
            .I(N__20320));
    Sp12to4 I__4504 (
            .O(N__20323),
            .I(N__20317));
    Sp12to4 I__4503 (
            .O(N__20320),
            .I(N__20314));
    Span12Mux_h I__4502 (
            .O(N__20317),
            .I(N__20309));
    Span12Mux_s5_v I__4501 (
            .O(N__20314),
            .I(N__20309));
    Odrv12 I__4500 (
            .O(N__20309),
            .I(n26));
    InMux I__4499 (
            .O(N__20306),
            .I(N__20303));
    LocalMux I__4498 (
            .O(N__20303),
            .I(N__20300));
    Span4Mux_v I__4497 (
            .O(N__20300),
            .I(N__20297));
    Span4Mux_h I__4496 (
            .O(N__20297),
            .I(N__20294));
    Sp12to4 I__4495 (
            .O(N__20294),
            .I(N__20291));
    Span12Mux_v I__4494 (
            .O(N__20291),
            .I(N__20288));
    Odrv12 I__4493 (
            .O(N__20288),
            .I(\line_buffer.n535 ));
    CascadeMux I__4492 (
            .O(N__20285),
            .I(N__20282));
    InMux I__4491 (
            .O(N__20282),
            .I(N__20279));
    LocalMux I__4490 (
            .O(N__20279),
            .I(N__20276));
    Span4Mux_h I__4489 (
            .O(N__20276),
            .I(N__20273));
    Sp12to4 I__4488 (
            .O(N__20273),
            .I(N__20270));
    Span12Mux_v I__4487 (
            .O(N__20270),
            .I(N__20267));
    Odrv12 I__4486 (
            .O(N__20267),
            .I(\line_buffer.n527 ));
    InMux I__4485 (
            .O(N__20264),
            .I(N__20248));
    InMux I__4484 (
            .O(N__20263),
            .I(N__20243));
    InMux I__4483 (
            .O(N__20262),
            .I(N__20243));
    InMux I__4482 (
            .O(N__20261),
            .I(N__20240));
    CascadeMux I__4481 (
            .O(N__20260),
            .I(N__20237));
    InMux I__4480 (
            .O(N__20259),
            .I(N__20233));
    InMux I__4479 (
            .O(N__20258),
            .I(N__20230));
    InMux I__4478 (
            .O(N__20257),
            .I(N__20227));
    InMux I__4477 (
            .O(N__20256),
            .I(N__20223));
    InMux I__4476 (
            .O(N__20255),
            .I(N__20220));
    InMux I__4475 (
            .O(N__20254),
            .I(N__20217));
    InMux I__4474 (
            .O(N__20253),
            .I(N__20214));
    InMux I__4473 (
            .O(N__20252),
            .I(N__20209));
    InMux I__4472 (
            .O(N__20251),
            .I(N__20209));
    LocalMux I__4471 (
            .O(N__20248),
            .I(N__20206));
    LocalMux I__4470 (
            .O(N__20243),
            .I(N__20201));
    LocalMux I__4469 (
            .O(N__20240),
            .I(N__20201));
    InMux I__4468 (
            .O(N__20237),
            .I(N__20196));
    InMux I__4467 (
            .O(N__20236),
            .I(N__20196));
    LocalMux I__4466 (
            .O(N__20233),
            .I(N__20190));
    LocalMux I__4465 (
            .O(N__20230),
            .I(N__20185));
    LocalMux I__4464 (
            .O(N__20227),
            .I(N__20185));
    InMux I__4463 (
            .O(N__20226),
            .I(N__20182));
    LocalMux I__4462 (
            .O(N__20223),
            .I(N__20172));
    LocalMux I__4461 (
            .O(N__20220),
            .I(N__20172));
    LocalMux I__4460 (
            .O(N__20217),
            .I(N__20172));
    LocalMux I__4459 (
            .O(N__20214),
            .I(N__20167));
    LocalMux I__4458 (
            .O(N__20209),
            .I(N__20167));
    Span4Mux_h I__4457 (
            .O(N__20206),
            .I(N__20164));
    Span4Mux_v I__4456 (
            .O(N__20201),
            .I(N__20156));
    LocalMux I__4455 (
            .O(N__20196),
            .I(N__20156));
    InMux I__4454 (
            .O(N__20195),
            .I(N__20153));
    InMux I__4453 (
            .O(N__20194),
            .I(N__20150));
    InMux I__4452 (
            .O(N__20193),
            .I(N__20147));
    Span4Mux_v I__4451 (
            .O(N__20190),
            .I(N__20144));
    Span4Mux_v I__4450 (
            .O(N__20185),
            .I(N__20141));
    LocalMux I__4449 (
            .O(N__20182),
            .I(N__20138));
    InMux I__4448 (
            .O(N__20181),
            .I(N__20135));
    InMux I__4447 (
            .O(N__20180),
            .I(N__20130));
    InMux I__4446 (
            .O(N__20179),
            .I(N__20130));
    Span4Mux_v I__4445 (
            .O(N__20172),
            .I(N__20122));
    Span4Mux_v I__4444 (
            .O(N__20167),
            .I(N__20122));
    Span4Mux_v I__4443 (
            .O(N__20164),
            .I(N__20119));
    InMux I__4442 (
            .O(N__20163),
            .I(N__20112));
    InMux I__4441 (
            .O(N__20162),
            .I(N__20112));
    InMux I__4440 (
            .O(N__20161),
            .I(N__20112));
    Span4Mux_v I__4439 (
            .O(N__20156),
            .I(N__20109));
    LocalMux I__4438 (
            .O(N__20153),
            .I(N__20104));
    LocalMux I__4437 (
            .O(N__20150),
            .I(N__20104));
    LocalMux I__4436 (
            .O(N__20147),
            .I(N__20091));
    Span4Mux_h I__4435 (
            .O(N__20144),
            .I(N__20091));
    Span4Mux_h I__4434 (
            .O(N__20141),
            .I(N__20091));
    Span4Mux_v I__4433 (
            .O(N__20138),
            .I(N__20091));
    LocalMux I__4432 (
            .O(N__20135),
            .I(N__20091));
    LocalMux I__4431 (
            .O(N__20130),
            .I(N__20091));
    InMux I__4430 (
            .O(N__20129),
            .I(N__20084));
    InMux I__4429 (
            .O(N__20128),
            .I(N__20084));
    InMux I__4428 (
            .O(N__20127),
            .I(N__20084));
    Odrv4 I__4427 (
            .O(N__20122),
            .I(\transmit_module.n3678 ));
    Odrv4 I__4426 (
            .O(N__20119),
            .I(\transmit_module.n3678 ));
    LocalMux I__4425 (
            .O(N__20112),
            .I(\transmit_module.n3678 ));
    Odrv4 I__4424 (
            .O(N__20109),
            .I(\transmit_module.n3678 ));
    Odrv12 I__4423 (
            .O(N__20104),
            .I(\transmit_module.n3678 ));
    Odrv4 I__4422 (
            .O(N__20091),
            .I(\transmit_module.n3678 ));
    LocalMux I__4421 (
            .O(N__20084),
            .I(\transmit_module.n3678 ));
    SRMux I__4420 (
            .O(N__20069),
            .I(N__20062));
    SRMux I__4419 (
            .O(N__20068),
            .I(N__20051));
    SRMux I__4418 (
            .O(N__20067),
            .I(N__20046));
    CascadeMux I__4417 (
            .O(N__20066),
            .I(N__20038));
    SRMux I__4416 (
            .O(N__20065),
            .I(N__20029));
    LocalMux I__4415 (
            .O(N__20062),
            .I(N__20026));
    SRMux I__4414 (
            .O(N__20061),
            .I(N__20023));
    SRMux I__4413 (
            .O(N__20060),
            .I(N__20020));
    CascadeMux I__4412 (
            .O(N__20059),
            .I(N__20014));
    SRMux I__4411 (
            .O(N__20058),
            .I(N__20008));
    SRMux I__4410 (
            .O(N__20057),
            .I(N__20003));
    SRMux I__4409 (
            .O(N__20056),
            .I(N__19998));
    SRMux I__4408 (
            .O(N__20055),
            .I(N__19991));
    SRMux I__4407 (
            .O(N__20054),
            .I(N__19988));
    LocalMux I__4406 (
            .O(N__20051),
            .I(N__19985));
    SRMux I__4405 (
            .O(N__20050),
            .I(N__19982));
    SRMux I__4404 (
            .O(N__20049),
            .I(N__19978));
    LocalMux I__4403 (
            .O(N__20046),
            .I(N__19975));
    SRMux I__4402 (
            .O(N__20045),
            .I(N__19972));
    SRMux I__4401 (
            .O(N__20044),
            .I(N__19968));
    SRMux I__4400 (
            .O(N__20043),
            .I(N__19965));
    SRMux I__4399 (
            .O(N__20042),
            .I(N__19960));
    SRMux I__4398 (
            .O(N__20041),
            .I(N__19957));
    InMux I__4397 (
            .O(N__20038),
            .I(N__19952));
    InMux I__4396 (
            .O(N__20037),
            .I(N__19952));
    SRMux I__4395 (
            .O(N__20036),
            .I(N__19948));
    CascadeMux I__4394 (
            .O(N__20035),
            .I(N__19945));
    CascadeMux I__4393 (
            .O(N__20034),
            .I(N__19942));
    CascadeMux I__4392 (
            .O(N__20033),
            .I(N__19939));
    SRMux I__4391 (
            .O(N__20032),
            .I(N__19936));
    LocalMux I__4390 (
            .O(N__20029),
            .I(N__19932));
    Span4Mux_v I__4389 (
            .O(N__20026),
            .I(N__19925));
    LocalMux I__4388 (
            .O(N__20023),
            .I(N__19925));
    LocalMux I__4387 (
            .O(N__20020),
            .I(N__19925));
    SRMux I__4386 (
            .O(N__20019),
            .I(N__19922));
    SRMux I__4385 (
            .O(N__20018),
            .I(N__19919));
    SRMux I__4384 (
            .O(N__20017),
            .I(N__19916));
    InMux I__4383 (
            .O(N__20014),
            .I(N__19913));
    CascadeMux I__4382 (
            .O(N__20013),
            .I(N__19907));
    SRMux I__4381 (
            .O(N__20012),
            .I(N__19904));
    SRMux I__4380 (
            .O(N__20011),
            .I(N__19901));
    LocalMux I__4379 (
            .O(N__20008),
            .I(N__19898));
    SRMux I__4378 (
            .O(N__20007),
            .I(N__19895));
    SRMux I__4377 (
            .O(N__20006),
            .I(N__19892));
    LocalMux I__4376 (
            .O(N__20003),
            .I(N__19889));
    SRMux I__4375 (
            .O(N__20002),
            .I(N__19886));
    SRMux I__4374 (
            .O(N__20001),
            .I(N__19883));
    LocalMux I__4373 (
            .O(N__19998),
            .I(N__19880));
    SRMux I__4372 (
            .O(N__19997),
            .I(N__19877));
    IoInMux I__4371 (
            .O(N__19996),
            .I(N__19870));
    CascadeMux I__4370 (
            .O(N__19995),
            .I(N__19867));
    SRMux I__4369 (
            .O(N__19994),
            .I(N__19863));
    LocalMux I__4368 (
            .O(N__19991),
            .I(N__19860));
    LocalMux I__4367 (
            .O(N__19988),
            .I(N__19857));
    Span4Mux_v I__4366 (
            .O(N__19985),
            .I(N__19852));
    LocalMux I__4365 (
            .O(N__19982),
            .I(N__19852));
    SRMux I__4364 (
            .O(N__19981),
            .I(N__19849));
    LocalMux I__4363 (
            .O(N__19978),
            .I(N__19842));
    Span4Mux_v I__4362 (
            .O(N__19975),
            .I(N__19842));
    LocalMux I__4361 (
            .O(N__19972),
            .I(N__19842));
    SRMux I__4360 (
            .O(N__19971),
            .I(N__19839));
    LocalMux I__4359 (
            .O(N__19968),
            .I(N__19831));
    LocalMux I__4358 (
            .O(N__19965),
            .I(N__19831));
    SRMux I__4357 (
            .O(N__19964),
            .I(N__19828));
    SRMux I__4356 (
            .O(N__19963),
            .I(N__19825));
    LocalMux I__4355 (
            .O(N__19960),
            .I(N__19818));
    LocalMux I__4354 (
            .O(N__19957),
            .I(N__19818));
    LocalMux I__4353 (
            .O(N__19952),
            .I(N__19818));
    CascadeMux I__4352 (
            .O(N__19951),
            .I(N__19815));
    LocalMux I__4351 (
            .O(N__19948),
            .I(N__19812));
    InMux I__4350 (
            .O(N__19945),
            .I(N__19807));
    InMux I__4349 (
            .O(N__19942),
            .I(N__19807));
    InMux I__4348 (
            .O(N__19939),
            .I(N__19804));
    LocalMux I__4347 (
            .O(N__19936),
            .I(N__19801));
    SRMux I__4346 (
            .O(N__19935),
            .I(N__19798));
    Span4Mux_h I__4345 (
            .O(N__19932),
            .I(N__19791));
    Span4Mux_h I__4344 (
            .O(N__19925),
            .I(N__19791));
    LocalMux I__4343 (
            .O(N__19922),
            .I(N__19791));
    LocalMux I__4342 (
            .O(N__19919),
            .I(N__19786));
    LocalMux I__4341 (
            .O(N__19916),
            .I(N__19786));
    LocalMux I__4340 (
            .O(N__19913),
            .I(N__19783));
    SRMux I__4339 (
            .O(N__19912),
            .I(N__19780));
    SRMux I__4338 (
            .O(N__19911),
            .I(N__19777));
    InMux I__4337 (
            .O(N__19910),
            .I(N__19772));
    InMux I__4336 (
            .O(N__19907),
            .I(N__19772));
    LocalMux I__4335 (
            .O(N__19904),
            .I(N__19769));
    LocalMux I__4334 (
            .O(N__19901),
            .I(N__19766));
    Span4Mux_v I__4333 (
            .O(N__19898),
            .I(N__19763));
    LocalMux I__4332 (
            .O(N__19895),
            .I(N__19758));
    LocalMux I__4331 (
            .O(N__19892),
            .I(N__19758));
    Span4Mux_h I__4330 (
            .O(N__19889),
            .I(N__19751));
    LocalMux I__4329 (
            .O(N__19886),
            .I(N__19751));
    LocalMux I__4328 (
            .O(N__19883),
            .I(N__19751));
    Span4Mux_h I__4327 (
            .O(N__19880),
            .I(N__19746));
    LocalMux I__4326 (
            .O(N__19877),
            .I(N__19746));
    SRMux I__4325 (
            .O(N__19876),
            .I(N__19743));
    CascadeMux I__4324 (
            .O(N__19875),
            .I(N__19740));
    InMux I__4323 (
            .O(N__19874),
            .I(N__19734));
    InMux I__4322 (
            .O(N__19873),
            .I(N__19734));
    LocalMux I__4321 (
            .O(N__19870),
            .I(N__19731));
    InMux I__4320 (
            .O(N__19867),
            .I(N__19728));
    CascadeMux I__4319 (
            .O(N__19866),
            .I(N__19724));
    LocalMux I__4318 (
            .O(N__19863),
            .I(N__19718));
    Span4Mux_v I__4317 (
            .O(N__19860),
            .I(N__19709));
    Span4Mux_h I__4316 (
            .O(N__19857),
            .I(N__19709));
    Span4Mux_v I__4315 (
            .O(N__19852),
            .I(N__19709));
    LocalMux I__4314 (
            .O(N__19849),
            .I(N__19709));
    Span4Mux_v I__4313 (
            .O(N__19842),
            .I(N__19704));
    LocalMux I__4312 (
            .O(N__19839),
            .I(N__19704));
    CascadeMux I__4311 (
            .O(N__19838),
            .I(N__19701));
    CascadeMux I__4310 (
            .O(N__19837),
            .I(N__19698));
    CascadeMux I__4309 (
            .O(N__19836),
            .I(N__19695));
    Span4Mux_h I__4308 (
            .O(N__19831),
            .I(N__19685));
    LocalMux I__4307 (
            .O(N__19828),
            .I(N__19685));
    LocalMux I__4306 (
            .O(N__19825),
            .I(N__19685));
    Span4Mux_v I__4305 (
            .O(N__19818),
            .I(N__19682));
    InMux I__4304 (
            .O(N__19815),
            .I(N__19679));
    Span4Mux_v I__4303 (
            .O(N__19812),
            .I(N__19674));
    LocalMux I__4302 (
            .O(N__19807),
            .I(N__19674));
    LocalMux I__4301 (
            .O(N__19804),
            .I(N__19671));
    Span4Mux_v I__4300 (
            .O(N__19801),
            .I(N__19660));
    LocalMux I__4299 (
            .O(N__19798),
            .I(N__19660));
    Span4Mux_h I__4298 (
            .O(N__19791),
            .I(N__19660));
    Span4Mux_v I__4297 (
            .O(N__19786),
            .I(N__19660));
    Span4Mux_h I__4296 (
            .O(N__19783),
            .I(N__19660));
    LocalMux I__4295 (
            .O(N__19780),
            .I(N__19653));
    LocalMux I__4294 (
            .O(N__19777),
            .I(N__19653));
    LocalMux I__4293 (
            .O(N__19772),
            .I(N__19653));
    Span4Mux_h I__4292 (
            .O(N__19769),
            .I(N__19638));
    Span4Mux_v I__4291 (
            .O(N__19766),
            .I(N__19638));
    Span4Mux_v I__4290 (
            .O(N__19763),
            .I(N__19638));
    Span4Mux_h I__4289 (
            .O(N__19758),
            .I(N__19638));
    Span4Mux_v I__4288 (
            .O(N__19751),
            .I(N__19638));
    Span4Mux_v I__4287 (
            .O(N__19746),
            .I(N__19638));
    LocalMux I__4286 (
            .O(N__19743),
            .I(N__19638));
    InMux I__4285 (
            .O(N__19740),
            .I(N__19633));
    InMux I__4284 (
            .O(N__19739),
            .I(N__19633));
    LocalMux I__4283 (
            .O(N__19734),
            .I(N__19630));
    Span12Mux_s0_h I__4282 (
            .O(N__19731),
            .I(N__19627));
    LocalMux I__4281 (
            .O(N__19728),
            .I(N__19624));
    InMux I__4280 (
            .O(N__19727),
            .I(N__19621));
    InMux I__4279 (
            .O(N__19724),
            .I(N__19616));
    InMux I__4278 (
            .O(N__19723),
            .I(N__19616));
    CascadeMux I__4277 (
            .O(N__19722),
            .I(N__19613));
    CascadeMux I__4276 (
            .O(N__19721),
            .I(N__19609));
    Span4Mux_v I__4275 (
            .O(N__19718),
            .I(N__19604));
    Span4Mux_v I__4274 (
            .O(N__19709),
            .I(N__19599));
    Span4Mux_h I__4273 (
            .O(N__19704),
            .I(N__19599));
    InMux I__4272 (
            .O(N__19701),
            .I(N__19596));
    InMux I__4271 (
            .O(N__19698),
            .I(N__19593));
    InMux I__4270 (
            .O(N__19695),
            .I(N__19586));
    InMux I__4269 (
            .O(N__19694),
            .I(N__19586));
    InMux I__4268 (
            .O(N__19693),
            .I(N__19586));
    InMux I__4267 (
            .O(N__19692),
            .I(N__19583));
    Span4Mux_v I__4266 (
            .O(N__19685),
            .I(N__19568));
    Span4Mux_h I__4265 (
            .O(N__19682),
            .I(N__19568));
    LocalMux I__4264 (
            .O(N__19679),
            .I(N__19568));
    Span4Mux_h I__4263 (
            .O(N__19674),
            .I(N__19568));
    Span4Mux_v I__4262 (
            .O(N__19671),
            .I(N__19568));
    Span4Mux_v I__4261 (
            .O(N__19660),
            .I(N__19568));
    Span4Mux_v I__4260 (
            .O(N__19653),
            .I(N__19568));
    Span4Mux_h I__4259 (
            .O(N__19638),
            .I(N__19561));
    LocalMux I__4258 (
            .O(N__19633),
            .I(N__19561));
    Span4Mux_v I__4257 (
            .O(N__19630),
            .I(N__19561));
    Span12Mux_h I__4256 (
            .O(N__19627),
            .I(N__19552));
    Sp12to4 I__4255 (
            .O(N__19624),
            .I(N__19552));
    LocalMux I__4254 (
            .O(N__19621),
            .I(N__19552));
    LocalMux I__4253 (
            .O(N__19616),
            .I(N__19552));
    InMux I__4252 (
            .O(N__19613),
            .I(N__19547));
    InMux I__4251 (
            .O(N__19612),
            .I(N__19547));
    InMux I__4250 (
            .O(N__19609),
            .I(N__19540));
    InMux I__4249 (
            .O(N__19608),
            .I(N__19540));
    InMux I__4248 (
            .O(N__19607),
            .I(N__19540));
    Odrv4 I__4247 (
            .O(N__19604),
            .I(ADV_VSYNC_c));
    Odrv4 I__4246 (
            .O(N__19599),
            .I(ADV_VSYNC_c));
    LocalMux I__4245 (
            .O(N__19596),
            .I(ADV_VSYNC_c));
    LocalMux I__4244 (
            .O(N__19593),
            .I(ADV_VSYNC_c));
    LocalMux I__4243 (
            .O(N__19586),
            .I(ADV_VSYNC_c));
    LocalMux I__4242 (
            .O(N__19583),
            .I(ADV_VSYNC_c));
    Odrv4 I__4241 (
            .O(N__19568),
            .I(ADV_VSYNC_c));
    Odrv4 I__4240 (
            .O(N__19561),
            .I(ADV_VSYNC_c));
    Odrv12 I__4239 (
            .O(N__19552),
            .I(ADV_VSYNC_c));
    LocalMux I__4238 (
            .O(N__19547),
            .I(ADV_VSYNC_c));
    LocalMux I__4237 (
            .O(N__19540),
            .I(ADV_VSYNC_c));
    InMux I__4236 (
            .O(N__19517),
            .I(N__19513));
    CascadeMux I__4235 (
            .O(N__19516),
            .I(N__19510));
    LocalMux I__4234 (
            .O(N__19513),
            .I(N__19507));
    InMux I__4233 (
            .O(N__19510),
            .I(N__19504));
    Odrv12 I__4232 (
            .O(N__19507),
            .I(\transmit_module.n113 ));
    LocalMux I__4231 (
            .O(N__19504),
            .I(\transmit_module.n113 ));
    InMux I__4230 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__4229 (
            .O(N__19496),
            .I(N__19492));
    InMux I__4228 (
            .O(N__19495),
            .I(N__19489));
    Span4Mux_v I__4227 (
            .O(N__19492),
            .I(N__19486));
    LocalMux I__4226 (
            .O(N__19489),
            .I(\transmit_module.n144 ));
    Odrv4 I__4225 (
            .O(N__19486),
            .I(\transmit_module.n144 ));
    CascadeMux I__4224 (
            .O(N__19481),
            .I(N__19477));
    CascadeMux I__4223 (
            .O(N__19480),
            .I(N__19474));
    CascadeBuf I__4222 (
            .O(N__19477),
            .I(N__19471));
    CascadeBuf I__4221 (
            .O(N__19474),
            .I(N__19468));
    CascadeMux I__4220 (
            .O(N__19471),
            .I(N__19465));
    CascadeMux I__4219 (
            .O(N__19468),
            .I(N__19462));
    CascadeBuf I__4218 (
            .O(N__19465),
            .I(N__19459));
    CascadeBuf I__4217 (
            .O(N__19462),
            .I(N__19456));
    CascadeMux I__4216 (
            .O(N__19459),
            .I(N__19453));
    CascadeMux I__4215 (
            .O(N__19456),
            .I(N__19450));
    CascadeBuf I__4214 (
            .O(N__19453),
            .I(N__19447));
    CascadeBuf I__4213 (
            .O(N__19450),
            .I(N__19444));
    CascadeMux I__4212 (
            .O(N__19447),
            .I(N__19441));
    CascadeMux I__4211 (
            .O(N__19444),
            .I(N__19438));
    CascadeBuf I__4210 (
            .O(N__19441),
            .I(N__19435));
    CascadeBuf I__4209 (
            .O(N__19438),
            .I(N__19432));
    CascadeMux I__4208 (
            .O(N__19435),
            .I(N__19429));
    CascadeMux I__4207 (
            .O(N__19432),
            .I(N__19426));
    CascadeBuf I__4206 (
            .O(N__19429),
            .I(N__19423));
    CascadeBuf I__4205 (
            .O(N__19426),
            .I(N__19420));
    CascadeMux I__4204 (
            .O(N__19423),
            .I(N__19417));
    CascadeMux I__4203 (
            .O(N__19420),
            .I(N__19414));
    CascadeBuf I__4202 (
            .O(N__19417),
            .I(N__19411));
    CascadeBuf I__4201 (
            .O(N__19414),
            .I(N__19408));
    CascadeMux I__4200 (
            .O(N__19411),
            .I(N__19405));
    CascadeMux I__4199 (
            .O(N__19408),
            .I(N__19402));
    CascadeBuf I__4198 (
            .O(N__19405),
            .I(N__19399));
    CascadeBuf I__4197 (
            .O(N__19402),
            .I(N__19396));
    CascadeMux I__4196 (
            .O(N__19399),
            .I(N__19393));
    CascadeMux I__4195 (
            .O(N__19396),
            .I(N__19390));
    CascadeBuf I__4194 (
            .O(N__19393),
            .I(N__19387));
    CascadeBuf I__4193 (
            .O(N__19390),
            .I(N__19384));
    CascadeMux I__4192 (
            .O(N__19387),
            .I(N__19381));
    CascadeMux I__4191 (
            .O(N__19384),
            .I(N__19378));
    CascadeBuf I__4190 (
            .O(N__19381),
            .I(N__19375));
    CascadeBuf I__4189 (
            .O(N__19378),
            .I(N__19372));
    CascadeMux I__4188 (
            .O(N__19375),
            .I(N__19369));
    CascadeMux I__4187 (
            .O(N__19372),
            .I(N__19366));
    CascadeBuf I__4186 (
            .O(N__19369),
            .I(N__19363));
    CascadeBuf I__4185 (
            .O(N__19366),
            .I(N__19360));
    CascadeMux I__4184 (
            .O(N__19363),
            .I(N__19357));
    CascadeMux I__4183 (
            .O(N__19360),
            .I(N__19354));
    CascadeBuf I__4182 (
            .O(N__19357),
            .I(N__19351));
    CascadeBuf I__4181 (
            .O(N__19354),
            .I(N__19348));
    CascadeMux I__4180 (
            .O(N__19351),
            .I(N__19345));
    CascadeMux I__4179 (
            .O(N__19348),
            .I(N__19342));
    CascadeBuf I__4178 (
            .O(N__19345),
            .I(N__19339));
    CascadeBuf I__4177 (
            .O(N__19342),
            .I(N__19336));
    CascadeMux I__4176 (
            .O(N__19339),
            .I(N__19333));
    CascadeMux I__4175 (
            .O(N__19336),
            .I(N__19330));
    CascadeBuf I__4174 (
            .O(N__19333),
            .I(N__19327));
    CascadeBuf I__4173 (
            .O(N__19330),
            .I(N__19324));
    CascadeMux I__4172 (
            .O(N__19327),
            .I(N__19321));
    CascadeMux I__4171 (
            .O(N__19324),
            .I(N__19318));
    CascadeBuf I__4170 (
            .O(N__19321),
            .I(N__19315));
    CascadeBuf I__4169 (
            .O(N__19318),
            .I(N__19312));
    CascadeMux I__4168 (
            .O(N__19315),
            .I(N__19309));
    CascadeMux I__4167 (
            .O(N__19312),
            .I(N__19306));
    CascadeBuf I__4166 (
            .O(N__19309),
            .I(N__19303));
    CascadeBuf I__4165 (
            .O(N__19306),
            .I(N__19300));
    CascadeMux I__4164 (
            .O(N__19303),
            .I(N__19297));
    CascadeMux I__4163 (
            .O(N__19300),
            .I(N__19294));
    InMux I__4162 (
            .O(N__19297),
            .I(N__19291));
    InMux I__4161 (
            .O(N__19294),
            .I(N__19288));
    LocalMux I__4160 (
            .O(N__19291),
            .I(N__19285));
    LocalMux I__4159 (
            .O(N__19288),
            .I(N__19282));
    Span12Mux_s11_h I__4158 (
            .O(N__19285),
            .I(N__19279));
    Sp12to4 I__4157 (
            .O(N__19282),
            .I(N__19276));
    Span12Mux_v I__4156 (
            .O(N__19279),
            .I(N__19271));
    Span12Mux_v I__4155 (
            .O(N__19276),
            .I(N__19271));
    Odrv12 I__4154 (
            .O(N__19271),
            .I(n25));
    IoInMux I__4153 (
            .O(N__19268),
            .I(N__19265));
    LocalMux I__4152 (
            .O(N__19265),
            .I(N__19260));
    IoInMux I__4151 (
            .O(N__19264),
            .I(N__19257));
    IoInMux I__4150 (
            .O(N__19263),
            .I(N__19254));
    IoSpan4Mux I__4149 (
            .O(N__19260),
            .I(N__19251));
    LocalMux I__4148 (
            .O(N__19257),
            .I(N__19248));
    LocalMux I__4147 (
            .O(N__19254),
            .I(N__19245));
    Span4Mux_s2_v I__4146 (
            .O(N__19251),
            .I(N__19242));
    IoSpan4Mux I__4145 (
            .O(N__19248),
            .I(N__19239));
    Span4Mux_s3_h I__4144 (
            .O(N__19245),
            .I(N__19236));
    Sp12to4 I__4143 (
            .O(N__19242),
            .I(N__19233));
    Span4Mux_s1_v I__4142 (
            .O(N__19239),
            .I(N__19230));
    Span4Mux_h I__4141 (
            .O(N__19236),
            .I(N__19227));
    Span12Mux_v I__4140 (
            .O(N__19233),
            .I(N__19224));
    Sp12to4 I__4139 (
            .O(N__19230),
            .I(N__19221));
    Span4Mux_h I__4138 (
            .O(N__19227),
            .I(N__19218));
    Span12Mux_h I__4137 (
            .O(N__19224),
            .I(N__19213));
    Span12Mux_h I__4136 (
            .O(N__19221),
            .I(N__19213));
    Span4Mux_h I__4135 (
            .O(N__19218),
            .I(N__19210));
    Odrv12 I__4134 (
            .O(N__19213),
            .I(n1818));
    Odrv4 I__4133 (
            .O(N__19210),
            .I(n1818));
    InMux I__4132 (
            .O(N__19205),
            .I(N__19202));
    LocalMux I__4131 (
            .O(N__19202),
            .I(N__19199));
    Sp12to4 I__4130 (
            .O(N__19199),
            .I(N__19196));
    Odrv12 I__4129 (
            .O(N__19196),
            .I(\line_buffer.n470 ));
    CascadeMux I__4128 (
            .O(N__19193),
            .I(N__19190));
    InMux I__4127 (
            .O(N__19190),
            .I(N__19187));
    LocalMux I__4126 (
            .O(N__19187),
            .I(N__19184));
    Span4Mux_v I__4125 (
            .O(N__19184),
            .I(N__19181));
    Sp12to4 I__4124 (
            .O(N__19181),
            .I(N__19178));
    Span12Mux_h I__4123 (
            .O(N__19178),
            .I(N__19175));
    Odrv12 I__4122 (
            .O(N__19175),
            .I(\line_buffer.n462 ));
    InMux I__4121 (
            .O(N__19172),
            .I(N__19169));
    LocalMux I__4120 (
            .O(N__19169),
            .I(N__19166));
    Odrv12 I__4119 (
            .O(N__19166),
            .I(\line_buffer.n3590 ));
    SRMux I__4118 (
            .O(N__19163),
            .I(N__19160));
    LocalMux I__4117 (
            .O(N__19160),
            .I(\receive_module.rx_counter.n2550 ));
    InMux I__4116 (
            .O(N__19157),
            .I(N__19154));
    LocalMux I__4115 (
            .O(N__19154),
            .I(N__19151));
    Odrv4 I__4114 (
            .O(N__19151),
            .I(\tvp_video_buffer.BUFFER_1_6 ));
    InMux I__4113 (
            .O(N__19148),
            .I(N__19143));
    InMux I__4112 (
            .O(N__19147),
            .I(N__19140));
    InMux I__4111 (
            .O(N__19146),
            .I(N__19137));
    LocalMux I__4110 (
            .O(N__19143),
            .I(N__19130));
    LocalMux I__4109 (
            .O(N__19140),
            .I(N__19130));
    LocalMux I__4108 (
            .O(N__19137),
            .I(N__19127));
    InMux I__4107 (
            .O(N__19136),
            .I(N__19124));
    InMux I__4106 (
            .O(N__19135),
            .I(N__19121));
    Span4Mux_v I__4105 (
            .O(N__19130),
            .I(N__19112));
    Span4Mux_h I__4104 (
            .O(N__19127),
            .I(N__19112));
    LocalMux I__4103 (
            .O(N__19124),
            .I(N__19112));
    LocalMux I__4102 (
            .O(N__19121),
            .I(N__19108));
    InMux I__4101 (
            .O(N__19120),
            .I(N__19105));
    InMux I__4100 (
            .O(N__19119),
            .I(N__19102));
    Span4Mux_v I__4099 (
            .O(N__19112),
            .I(N__19099));
    InMux I__4098 (
            .O(N__19111),
            .I(N__19096));
    Span4Mux_v I__4097 (
            .O(N__19108),
            .I(N__19093));
    LocalMux I__4096 (
            .O(N__19105),
            .I(N__19090));
    LocalMux I__4095 (
            .O(N__19102),
            .I(N__19087));
    Span4Mux_v I__4094 (
            .O(N__19099),
            .I(N__19082));
    LocalMux I__4093 (
            .O(N__19096),
            .I(N__19082));
    Sp12to4 I__4092 (
            .O(N__19093),
            .I(N__19078));
    Span4Mux_s2_v I__4091 (
            .O(N__19090),
            .I(N__19073));
    Span4Mux_v I__4090 (
            .O(N__19087),
            .I(N__19073));
    Span4Mux_v I__4089 (
            .O(N__19082),
            .I(N__19070));
    InMux I__4088 (
            .O(N__19081),
            .I(N__19067));
    Span12Mux_h I__4087 (
            .O(N__19078),
            .I(N__19064));
    Sp12to4 I__4086 (
            .O(N__19073),
            .I(N__19061));
    Span4Mux_h I__4085 (
            .O(N__19070),
            .I(N__19056));
    LocalMux I__4084 (
            .O(N__19067),
            .I(N__19056));
    Span12Mux_v I__4083 (
            .O(N__19064),
            .I(N__19051));
    Span12Mux_h I__4082 (
            .O(N__19061),
            .I(N__19051));
    Span4Mux_h I__4081 (
            .O(N__19056),
            .I(N__19048));
    Odrv12 I__4080 (
            .O(N__19051),
            .I(RX_DATA_6));
    Odrv4 I__4079 (
            .O(N__19048),
            .I(RX_DATA_6));
    InMux I__4078 (
            .O(N__19043),
            .I(N__19040));
    LocalMux I__4077 (
            .O(N__19040),
            .I(N__19037));
    Span4Mux_v I__4076 (
            .O(N__19037),
            .I(N__19031));
    InMux I__4075 (
            .O(N__19036),
            .I(N__19028));
    InMux I__4074 (
            .O(N__19035),
            .I(N__19025));
    InMux I__4073 (
            .O(N__19034),
            .I(N__19022));
    Span4Mux_v I__4072 (
            .O(N__19031),
            .I(N__19016));
    LocalMux I__4071 (
            .O(N__19028),
            .I(N__19016));
    LocalMux I__4070 (
            .O(N__19025),
            .I(N__19013));
    LocalMux I__4069 (
            .O(N__19022),
            .I(N__19010));
    InMux I__4068 (
            .O(N__19021),
            .I(N__19007));
    Span4Mux_v I__4067 (
            .O(N__19016),
            .I(N__19003));
    Sp12to4 I__4066 (
            .O(N__19013),
            .I(N__18998));
    Span4Mux_h I__4065 (
            .O(N__19010),
            .I(N__18995));
    LocalMux I__4064 (
            .O(N__19007),
            .I(N__18992));
    InMux I__4063 (
            .O(N__19006),
            .I(N__18989));
    Span4Mux_v I__4062 (
            .O(N__19003),
            .I(N__18986));
    InMux I__4061 (
            .O(N__19002),
            .I(N__18983));
    InMux I__4060 (
            .O(N__19001),
            .I(N__18980));
    Span12Mux_s9_v I__4059 (
            .O(N__18998),
            .I(N__18977));
    Span4Mux_h I__4058 (
            .O(N__18995),
            .I(N__18974));
    Span4Mux_h I__4057 (
            .O(N__18992),
            .I(N__18971));
    LocalMux I__4056 (
            .O(N__18989),
            .I(N__18968));
    Sp12to4 I__4055 (
            .O(N__18986),
            .I(N__18963));
    LocalMux I__4054 (
            .O(N__18983),
            .I(N__18963));
    LocalMux I__4053 (
            .O(N__18980),
            .I(N__18960));
    Span12Mux_v I__4052 (
            .O(N__18977),
            .I(N__18956));
    Span4Mux_h I__4051 (
            .O(N__18974),
            .I(N__18951));
    Span4Mux_h I__4050 (
            .O(N__18971),
            .I(N__18951));
    Span12Mux_h I__4049 (
            .O(N__18968),
            .I(N__18944));
    Span12Mux_h I__4048 (
            .O(N__18963),
            .I(N__18944));
    Span12Mux_h I__4047 (
            .O(N__18960),
            .I(N__18944));
    InMux I__4046 (
            .O(N__18959),
            .I(N__18941));
    Odrv12 I__4045 (
            .O(N__18956),
            .I(RX_DATA_4));
    Odrv4 I__4044 (
            .O(N__18951),
            .I(RX_DATA_4));
    Odrv12 I__4043 (
            .O(N__18944),
            .I(RX_DATA_4));
    LocalMux I__4042 (
            .O(N__18941),
            .I(RX_DATA_4));
    CascadeMux I__4041 (
            .O(N__18932),
            .I(\receive_module.sync_wd.n6_cascade_ ));
    CascadeMux I__4040 (
            .O(N__18929),
            .I(\receive_module.sync_wd.n4_cascade_ ));
    InMux I__4039 (
            .O(N__18926),
            .I(N__18920));
    InMux I__4038 (
            .O(N__18925),
            .I(N__18920));
    LocalMux I__4037 (
            .O(N__18920),
            .I(N__18915));
    InMux I__4036 (
            .O(N__18919),
            .I(N__18912));
    InMux I__4035 (
            .O(N__18918),
            .I(N__18909));
    Span4Mux_s2_v I__4034 (
            .O(N__18915),
            .I(N__18901));
    LocalMux I__4033 (
            .O(N__18912),
            .I(N__18901));
    LocalMux I__4032 (
            .O(N__18909),
            .I(N__18901));
    InMux I__4031 (
            .O(N__18908),
            .I(N__18898));
    Span4Mux_v I__4030 (
            .O(N__18901),
            .I(N__18887));
    LocalMux I__4029 (
            .O(N__18898),
            .I(N__18887));
    InMux I__4028 (
            .O(N__18897),
            .I(N__18880));
    InMux I__4027 (
            .O(N__18896),
            .I(N__18880));
    InMux I__4026 (
            .O(N__18895),
            .I(N__18880));
    InMux I__4025 (
            .O(N__18894),
            .I(N__18873));
    InMux I__4024 (
            .O(N__18893),
            .I(N__18873));
    InMux I__4023 (
            .O(N__18892),
            .I(N__18873));
    Span4Mux_v I__4022 (
            .O(N__18887),
            .I(N__18863));
    LocalMux I__4021 (
            .O(N__18880),
            .I(N__18863));
    LocalMux I__4020 (
            .O(N__18873),
            .I(N__18863));
    InMux I__4019 (
            .O(N__18872),
            .I(N__18855));
    InMux I__4018 (
            .O(N__18871),
            .I(N__18855));
    InMux I__4017 (
            .O(N__18870),
            .I(N__18855));
    Span4Mux_v I__4016 (
            .O(N__18863),
            .I(N__18851));
    InMux I__4015 (
            .O(N__18862),
            .I(N__18848));
    LocalMux I__4014 (
            .O(N__18855),
            .I(N__18845));
    InMux I__4013 (
            .O(N__18854),
            .I(N__18840));
    Span4Mux_v I__4012 (
            .O(N__18851),
            .I(N__18835));
    LocalMux I__4011 (
            .O(N__18848),
            .I(N__18835));
    Span4Mux_h I__4010 (
            .O(N__18845),
            .I(N__18832));
    InMux I__4009 (
            .O(N__18844),
            .I(N__18827));
    InMux I__4008 (
            .O(N__18843),
            .I(N__18827));
    LocalMux I__4007 (
            .O(N__18840),
            .I(TVP_VSYNC_buff));
    Odrv4 I__4006 (
            .O(N__18835),
            .I(TVP_VSYNC_buff));
    Odrv4 I__4005 (
            .O(N__18832),
            .I(TVP_VSYNC_buff));
    LocalMux I__4004 (
            .O(N__18827),
            .I(TVP_VSYNC_buff));
    IoInMux I__4003 (
            .O(N__18818),
            .I(N__18815));
    LocalMux I__4002 (
            .O(N__18815),
            .I(N__18812));
    Span4Mux_s3_h I__4001 (
            .O(N__18812),
            .I(N__18809));
    Sp12to4 I__4000 (
            .O(N__18809),
            .I(N__18806));
    Span12Mux_v I__3999 (
            .O(N__18806),
            .I(N__18802));
    InMux I__3998 (
            .O(N__18805),
            .I(N__18799));
    Span12Mux_h I__3997 (
            .O(N__18802),
            .I(N__18793));
    LocalMux I__3996 (
            .O(N__18799),
            .I(N__18793));
    InMux I__3995 (
            .O(N__18798),
            .I(N__18790));
    Odrv12 I__3994 (
            .O(N__18793),
            .I(DEBUG_c_0));
    LocalMux I__3993 (
            .O(N__18790),
            .I(DEBUG_c_0));
    CascadeMux I__3992 (
            .O(N__18785),
            .I(N__18781));
    CascadeMux I__3991 (
            .O(N__18784),
            .I(N__18778));
    InMux I__3990 (
            .O(N__18781),
            .I(N__18772));
    InMux I__3989 (
            .O(N__18778),
            .I(N__18772));
    CascadeMux I__3988 (
            .O(N__18777),
            .I(N__18769));
    LocalMux I__3987 (
            .O(N__18772),
            .I(N__18763));
    InMux I__3986 (
            .O(N__18769),
            .I(N__18760));
    CascadeMux I__3985 (
            .O(N__18768),
            .I(N__18757));
    IoInMux I__3984 (
            .O(N__18767),
            .I(N__18750));
    CascadeMux I__3983 (
            .O(N__18766),
            .I(N__18747));
    Span4Mux_h I__3982 (
            .O(N__18763),
            .I(N__18744));
    LocalMux I__3981 (
            .O(N__18760),
            .I(N__18741));
    InMux I__3980 (
            .O(N__18757),
            .I(N__18738));
    CascadeMux I__3979 (
            .O(N__18756),
            .I(N__18734));
    CascadeMux I__3978 (
            .O(N__18755),
            .I(N__18730));
    CascadeMux I__3977 (
            .O(N__18754),
            .I(N__18727));
    CascadeMux I__3976 (
            .O(N__18753),
            .I(N__18724));
    LocalMux I__3975 (
            .O(N__18750),
            .I(N__18721));
    InMux I__3974 (
            .O(N__18747),
            .I(N__18718));
    Span4Mux_v I__3973 (
            .O(N__18744),
            .I(N__18713));
    Span4Mux_h I__3972 (
            .O(N__18741),
            .I(N__18713));
    LocalMux I__3971 (
            .O(N__18738),
            .I(N__18710));
    InMux I__3970 (
            .O(N__18737),
            .I(N__18697));
    InMux I__3969 (
            .O(N__18734),
            .I(N__18697));
    InMux I__3968 (
            .O(N__18733),
            .I(N__18697));
    InMux I__3967 (
            .O(N__18730),
            .I(N__18697));
    InMux I__3966 (
            .O(N__18727),
            .I(N__18697));
    InMux I__3965 (
            .O(N__18724),
            .I(N__18697));
    Span12Mux_s1_h I__3964 (
            .O(N__18721),
            .I(N__18694));
    LocalMux I__3963 (
            .O(N__18718),
            .I(N__18691));
    Span4Mux_v I__3962 (
            .O(N__18713),
            .I(N__18686));
    Span4Mux_h I__3961 (
            .O(N__18710),
            .I(N__18686));
    LocalMux I__3960 (
            .O(N__18697),
            .I(N__18683));
    Span12Mux_h I__3959 (
            .O(N__18694),
            .I(N__18675));
    Span12Mux_h I__3958 (
            .O(N__18691),
            .I(N__18675));
    Span4Mux_v I__3957 (
            .O(N__18686),
            .I(N__18670));
    Span4Mux_h I__3956 (
            .O(N__18683),
            .I(N__18670));
    InMux I__3955 (
            .O(N__18682),
            .I(N__18666));
    InMux I__3954 (
            .O(N__18681),
            .I(N__18654));
    InMux I__3953 (
            .O(N__18680),
            .I(N__18654));
    Span12Mux_v I__3952 (
            .O(N__18675),
            .I(N__18651));
    Span4Mux_v I__3951 (
            .O(N__18670),
            .I(N__18648));
    InMux I__3950 (
            .O(N__18669),
            .I(N__18645));
    LocalMux I__3949 (
            .O(N__18666),
            .I(N__18642));
    InMux I__3948 (
            .O(N__18665),
            .I(N__18635));
    InMux I__3947 (
            .O(N__18664),
            .I(N__18635));
    InMux I__3946 (
            .O(N__18663),
            .I(N__18635));
    InMux I__3945 (
            .O(N__18662),
            .I(N__18632));
    InMux I__3944 (
            .O(N__18661),
            .I(N__18627));
    InMux I__3943 (
            .O(N__18660),
            .I(N__18627));
    InMux I__3942 (
            .O(N__18659),
            .I(N__18624));
    LocalMux I__3941 (
            .O(N__18654),
            .I(N__18621));
    Odrv12 I__3940 (
            .O(N__18651),
            .I(DEBUG_c_4));
    Odrv4 I__3939 (
            .O(N__18648),
            .I(DEBUG_c_4));
    LocalMux I__3938 (
            .O(N__18645),
            .I(DEBUG_c_4));
    Odrv4 I__3937 (
            .O(N__18642),
            .I(DEBUG_c_4));
    LocalMux I__3936 (
            .O(N__18635),
            .I(DEBUG_c_4));
    LocalMux I__3935 (
            .O(N__18632),
            .I(DEBUG_c_4));
    LocalMux I__3934 (
            .O(N__18627),
            .I(DEBUG_c_4));
    LocalMux I__3933 (
            .O(N__18624),
            .I(DEBUG_c_4));
    Odrv4 I__3932 (
            .O(N__18621),
            .I(DEBUG_c_4));
    InMux I__3931 (
            .O(N__18602),
            .I(N__18599));
    LocalMux I__3930 (
            .O(N__18599),
            .I(\receive_module.sync_wd.old_visible ));
    InMux I__3929 (
            .O(N__18596),
            .I(N__18593));
    LocalMux I__3928 (
            .O(N__18593),
            .I(N__18588));
    InMux I__3927 (
            .O(N__18592),
            .I(N__18585));
    InMux I__3926 (
            .O(N__18591),
            .I(N__18582));
    Span4Mux_v I__3925 (
            .O(N__18588),
            .I(N__18572));
    LocalMux I__3924 (
            .O(N__18585),
            .I(N__18572));
    LocalMux I__3923 (
            .O(N__18582),
            .I(N__18572));
    InMux I__3922 (
            .O(N__18581),
            .I(N__18569));
    InMux I__3921 (
            .O(N__18580),
            .I(N__18566));
    InMux I__3920 (
            .O(N__18579),
            .I(N__18563));
    Span4Mux_v I__3919 (
            .O(N__18572),
            .I(N__18558));
    LocalMux I__3918 (
            .O(N__18569),
            .I(N__18558));
    LocalMux I__3917 (
            .O(N__18566),
            .I(N__18553));
    LocalMux I__3916 (
            .O(N__18563),
            .I(N__18550));
    Span4Mux_v I__3915 (
            .O(N__18558),
            .I(N__18547));
    InMux I__3914 (
            .O(N__18557),
            .I(N__18544));
    InMux I__3913 (
            .O(N__18556),
            .I(N__18541));
    Span12Mux_s10_h I__3912 (
            .O(N__18553),
            .I(N__18538));
    Span12Mux_s10_h I__3911 (
            .O(N__18550),
            .I(N__18535));
    Span4Mux_h I__3910 (
            .O(N__18547),
            .I(N__18532));
    LocalMux I__3909 (
            .O(N__18544),
            .I(N__18529));
    LocalMux I__3908 (
            .O(N__18541),
            .I(N__18526));
    Span12Mux_v I__3907 (
            .O(N__18538),
            .I(N__18520));
    Span12Mux_v I__3906 (
            .O(N__18535),
            .I(N__18520));
    Span4Mux_v I__3905 (
            .O(N__18532),
            .I(N__18517));
    Span12Mux_h I__3904 (
            .O(N__18529),
            .I(N__18512));
    Span12Mux_h I__3903 (
            .O(N__18526),
            .I(N__18512));
    InMux I__3902 (
            .O(N__18525),
            .I(N__18509));
    Odrv12 I__3901 (
            .O(N__18520),
            .I(RX_DATA_7));
    Odrv4 I__3900 (
            .O(N__18517),
            .I(RX_DATA_7));
    Odrv12 I__3899 (
            .O(N__18512),
            .I(RX_DATA_7));
    LocalMux I__3898 (
            .O(N__18509),
            .I(RX_DATA_7));
    InMux I__3897 (
            .O(N__18500),
            .I(N__18497));
    LocalMux I__3896 (
            .O(N__18497),
            .I(N__18494));
    Span4Mux_v I__3895 (
            .O(N__18494),
            .I(N__18491));
    Span4Mux_h I__3894 (
            .O(N__18491),
            .I(N__18488));
    Span4Mux_h I__3893 (
            .O(N__18488),
            .I(N__18485));
    Odrv4 I__3892 (
            .O(N__18485),
            .I(\line_buffer.n569 ));
    InMux I__3891 (
            .O(N__18482),
            .I(N__18479));
    LocalMux I__3890 (
            .O(N__18479),
            .I(N__18476));
    Span4Mux_v I__3889 (
            .O(N__18476),
            .I(N__18473));
    Sp12to4 I__3888 (
            .O(N__18473),
            .I(N__18470));
    Odrv12 I__3887 (
            .O(N__18470),
            .I(\line_buffer.n561 ));
    InMux I__3886 (
            .O(N__18467),
            .I(N__18464));
    LocalMux I__3885 (
            .O(N__18464),
            .I(N__18461));
    Span4Mux_v I__3884 (
            .O(N__18461),
            .I(N__18458));
    Span4Mux_h I__3883 (
            .O(N__18458),
            .I(N__18455));
    Span4Mux_h I__3882 (
            .O(N__18455),
            .I(N__18452));
    Odrv4 I__3881 (
            .O(N__18452),
            .I(\line_buffer.n567 ));
    InMux I__3880 (
            .O(N__18449),
            .I(N__18446));
    LocalMux I__3879 (
            .O(N__18446),
            .I(N__18443));
    Span12Mux_h I__3878 (
            .O(N__18443),
            .I(N__18440));
    Odrv12 I__3877 (
            .O(N__18440),
            .I(\line_buffer.n559 ));
    CascadeMux I__3876 (
            .O(N__18437),
            .I(\receive_module.rx_counter.n3522_cascade_ ));
    InMux I__3875 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__3874 (
            .O(N__18431),
            .I(\receive_module.rx_counter.n7_adj_619 ));
    InMux I__3873 (
            .O(N__18428),
            .I(N__18424));
    InMux I__3872 (
            .O(N__18427),
            .I(N__18421));
    LocalMux I__3871 (
            .O(N__18424),
            .I(\receive_module.rx_counter.n11 ));
    LocalMux I__3870 (
            .O(N__18421),
            .I(\receive_module.rx_counter.n11 ));
    InMux I__3869 (
            .O(N__18416),
            .I(N__18412));
    InMux I__3868 (
            .O(N__18415),
            .I(N__18409));
    LocalMux I__3867 (
            .O(N__18412),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    LocalMux I__3866 (
            .O(N__18409),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    InMux I__3865 (
            .O(N__18404),
            .I(bfn_16_10_0_));
    InMux I__3864 (
            .O(N__18401),
            .I(N__18397));
    InMux I__3863 (
            .O(N__18400),
            .I(N__18394));
    LocalMux I__3862 (
            .O(N__18397),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    LocalMux I__3861 (
            .O(N__18394),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    InMux I__3860 (
            .O(N__18389),
            .I(\receive_module.rx_counter.n3205 ));
    InMux I__3859 (
            .O(N__18386),
            .I(N__18382));
    InMux I__3858 (
            .O(N__18385),
            .I(N__18379));
    LocalMux I__3857 (
            .O(N__18382),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    LocalMux I__3856 (
            .O(N__18379),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    InMux I__3855 (
            .O(N__18374),
            .I(\receive_module.rx_counter.n3206 ));
    InMux I__3854 (
            .O(N__18371),
            .I(N__18367));
    InMux I__3853 (
            .O(N__18370),
            .I(N__18364));
    LocalMux I__3852 (
            .O(N__18367),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    LocalMux I__3851 (
            .O(N__18364),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    InMux I__3850 (
            .O(N__18359),
            .I(\receive_module.rx_counter.n3207 ));
    InMux I__3849 (
            .O(N__18356),
            .I(N__18352));
    InMux I__3848 (
            .O(N__18355),
            .I(N__18349));
    LocalMux I__3847 (
            .O(N__18352),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    LocalMux I__3846 (
            .O(N__18349),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    InMux I__3845 (
            .O(N__18344),
            .I(\receive_module.rx_counter.n3208 ));
    InMux I__3844 (
            .O(N__18341),
            .I(\receive_module.rx_counter.n3209 ));
    InMux I__3843 (
            .O(N__18338),
            .I(N__18334));
    InMux I__3842 (
            .O(N__18337),
            .I(N__18331));
    LocalMux I__3841 (
            .O(N__18334),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    LocalMux I__3840 (
            .O(N__18331),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    CEMux I__3839 (
            .O(N__18326),
            .I(N__18322));
    CEMux I__3838 (
            .O(N__18325),
            .I(N__18319));
    LocalMux I__3837 (
            .O(N__18322),
            .I(N__18316));
    LocalMux I__3836 (
            .O(N__18319),
            .I(N__18313));
    Span4Mux_v I__3835 (
            .O(N__18316),
            .I(N__18310));
    Span4Mux_h I__3834 (
            .O(N__18313),
            .I(N__18307));
    Odrv4 I__3833 (
            .O(N__18310),
            .I(\receive_module.rx_counter.n3675 ));
    Odrv4 I__3832 (
            .O(N__18307),
            .I(\receive_module.rx_counter.n3675 ));
    InMux I__3831 (
            .O(N__18302),
            .I(N__18299));
    LocalMux I__3830 (
            .O(N__18299),
            .I(N__18296));
    Span12Mux_s9_v I__3829 (
            .O(N__18296),
            .I(N__18293));
    Span12Mux_v I__3828 (
            .O(N__18293),
            .I(N__18290));
    Odrv12 I__3827 (
            .O(N__18290),
            .I(\receive_module.n137 ));
    CascadeMux I__3826 (
            .O(N__18287),
            .I(N__18284));
    CascadeBuf I__3825 (
            .O(N__18284),
            .I(N__18281));
    CascadeMux I__3824 (
            .O(N__18281),
            .I(N__18277));
    CascadeMux I__3823 (
            .O(N__18280),
            .I(N__18274));
    CascadeBuf I__3822 (
            .O(N__18277),
            .I(N__18271));
    CascadeBuf I__3821 (
            .O(N__18274),
            .I(N__18268));
    CascadeMux I__3820 (
            .O(N__18271),
            .I(N__18265));
    CascadeMux I__3819 (
            .O(N__18268),
            .I(N__18262));
    CascadeBuf I__3818 (
            .O(N__18265),
            .I(N__18259));
    CascadeBuf I__3817 (
            .O(N__18262),
            .I(N__18256));
    CascadeMux I__3816 (
            .O(N__18259),
            .I(N__18253));
    CascadeMux I__3815 (
            .O(N__18256),
            .I(N__18250));
    CascadeBuf I__3814 (
            .O(N__18253),
            .I(N__18247));
    CascadeBuf I__3813 (
            .O(N__18250),
            .I(N__18244));
    CascadeMux I__3812 (
            .O(N__18247),
            .I(N__18241));
    CascadeMux I__3811 (
            .O(N__18244),
            .I(N__18238));
    CascadeBuf I__3810 (
            .O(N__18241),
            .I(N__18235));
    CascadeBuf I__3809 (
            .O(N__18238),
            .I(N__18232));
    CascadeMux I__3808 (
            .O(N__18235),
            .I(N__18229));
    CascadeMux I__3807 (
            .O(N__18232),
            .I(N__18226));
    CascadeBuf I__3806 (
            .O(N__18229),
            .I(N__18223));
    CascadeBuf I__3805 (
            .O(N__18226),
            .I(N__18220));
    CascadeMux I__3804 (
            .O(N__18223),
            .I(N__18217));
    CascadeMux I__3803 (
            .O(N__18220),
            .I(N__18214));
    CascadeBuf I__3802 (
            .O(N__18217),
            .I(N__18211));
    CascadeBuf I__3801 (
            .O(N__18214),
            .I(N__18208));
    CascadeMux I__3800 (
            .O(N__18211),
            .I(N__18205));
    CascadeMux I__3799 (
            .O(N__18208),
            .I(N__18202));
    CascadeBuf I__3798 (
            .O(N__18205),
            .I(N__18199));
    CascadeBuf I__3797 (
            .O(N__18202),
            .I(N__18196));
    CascadeMux I__3796 (
            .O(N__18199),
            .I(N__18193));
    CascadeMux I__3795 (
            .O(N__18196),
            .I(N__18190));
    CascadeBuf I__3794 (
            .O(N__18193),
            .I(N__18187));
    CascadeBuf I__3793 (
            .O(N__18190),
            .I(N__18184));
    CascadeMux I__3792 (
            .O(N__18187),
            .I(N__18181));
    CascadeMux I__3791 (
            .O(N__18184),
            .I(N__18178));
    CascadeBuf I__3790 (
            .O(N__18181),
            .I(N__18175));
    CascadeBuf I__3789 (
            .O(N__18178),
            .I(N__18172));
    CascadeMux I__3788 (
            .O(N__18175),
            .I(N__18169));
    CascadeMux I__3787 (
            .O(N__18172),
            .I(N__18166));
    CascadeBuf I__3786 (
            .O(N__18169),
            .I(N__18163));
    CascadeBuf I__3785 (
            .O(N__18166),
            .I(N__18160));
    CascadeMux I__3784 (
            .O(N__18163),
            .I(N__18157));
    CascadeMux I__3783 (
            .O(N__18160),
            .I(N__18154));
    CascadeBuf I__3782 (
            .O(N__18157),
            .I(N__18151));
    CascadeBuf I__3781 (
            .O(N__18154),
            .I(N__18148));
    CascadeMux I__3780 (
            .O(N__18151),
            .I(N__18145));
    CascadeMux I__3779 (
            .O(N__18148),
            .I(N__18142));
    CascadeBuf I__3778 (
            .O(N__18145),
            .I(N__18139));
    CascadeBuf I__3777 (
            .O(N__18142),
            .I(N__18136));
    CascadeMux I__3776 (
            .O(N__18139),
            .I(N__18133));
    CascadeMux I__3775 (
            .O(N__18136),
            .I(N__18130));
    CascadeBuf I__3774 (
            .O(N__18133),
            .I(N__18127));
    CascadeBuf I__3773 (
            .O(N__18130),
            .I(N__18124));
    CascadeMux I__3772 (
            .O(N__18127),
            .I(N__18121));
    CascadeMux I__3771 (
            .O(N__18124),
            .I(N__18118));
    CascadeBuf I__3770 (
            .O(N__18121),
            .I(N__18115));
    CascadeBuf I__3769 (
            .O(N__18118),
            .I(N__18112));
    CascadeMux I__3768 (
            .O(N__18115),
            .I(N__18109));
    CascadeMux I__3767 (
            .O(N__18112),
            .I(N__18106));
    InMux I__3766 (
            .O(N__18109),
            .I(N__18103));
    CascadeBuf I__3765 (
            .O(N__18106),
            .I(N__18100));
    LocalMux I__3764 (
            .O(N__18103),
            .I(N__18096));
    CascadeMux I__3763 (
            .O(N__18100),
            .I(N__18093));
    InMux I__3762 (
            .O(N__18099),
            .I(N__18090));
    Span4Mux_h I__3761 (
            .O(N__18096),
            .I(N__18087));
    InMux I__3760 (
            .O(N__18093),
            .I(N__18084));
    LocalMux I__3759 (
            .O(N__18090),
            .I(N__18081));
    Span4Mux_v I__3758 (
            .O(N__18087),
            .I(N__18077));
    LocalMux I__3757 (
            .O(N__18084),
            .I(N__18074));
    Span12Mux_v I__3756 (
            .O(N__18081),
            .I(N__18071));
    InMux I__3755 (
            .O(N__18080),
            .I(N__18068));
    Sp12to4 I__3754 (
            .O(N__18077),
            .I(N__18063));
    Span12Mux_s4_v I__3753 (
            .O(N__18074),
            .I(N__18063));
    Odrv12 I__3752 (
            .O(N__18071),
            .I(RX_ADDR_0));
    LocalMux I__3751 (
            .O(N__18068),
            .I(RX_ADDR_0));
    Odrv12 I__3750 (
            .O(N__18063),
            .I(RX_ADDR_0));
    InMux I__3749 (
            .O(N__18056),
            .I(N__18053));
    LocalMux I__3748 (
            .O(N__18053),
            .I(N__18050));
    Span12Mux_s10_v I__3747 (
            .O(N__18050),
            .I(N__18047));
    Odrv12 I__3746 (
            .O(N__18047),
            .I(\receive_module.n134 ));
    CascadeMux I__3745 (
            .O(N__18044),
            .I(N__18040));
    CascadeMux I__3744 (
            .O(N__18043),
            .I(N__18037));
    CascadeBuf I__3743 (
            .O(N__18040),
            .I(N__18034));
    CascadeBuf I__3742 (
            .O(N__18037),
            .I(N__18031));
    CascadeMux I__3741 (
            .O(N__18034),
            .I(N__18028));
    CascadeMux I__3740 (
            .O(N__18031),
            .I(N__18025));
    CascadeBuf I__3739 (
            .O(N__18028),
            .I(N__18022));
    CascadeBuf I__3738 (
            .O(N__18025),
            .I(N__18019));
    CascadeMux I__3737 (
            .O(N__18022),
            .I(N__18016));
    CascadeMux I__3736 (
            .O(N__18019),
            .I(N__18013));
    CascadeBuf I__3735 (
            .O(N__18016),
            .I(N__18010));
    CascadeBuf I__3734 (
            .O(N__18013),
            .I(N__18007));
    CascadeMux I__3733 (
            .O(N__18010),
            .I(N__18004));
    CascadeMux I__3732 (
            .O(N__18007),
            .I(N__18001));
    CascadeBuf I__3731 (
            .O(N__18004),
            .I(N__17998));
    CascadeBuf I__3730 (
            .O(N__18001),
            .I(N__17995));
    CascadeMux I__3729 (
            .O(N__17998),
            .I(N__17992));
    CascadeMux I__3728 (
            .O(N__17995),
            .I(N__17989));
    CascadeBuf I__3727 (
            .O(N__17992),
            .I(N__17986));
    CascadeBuf I__3726 (
            .O(N__17989),
            .I(N__17983));
    CascadeMux I__3725 (
            .O(N__17986),
            .I(N__17980));
    CascadeMux I__3724 (
            .O(N__17983),
            .I(N__17977));
    CascadeBuf I__3723 (
            .O(N__17980),
            .I(N__17974));
    CascadeBuf I__3722 (
            .O(N__17977),
            .I(N__17971));
    CascadeMux I__3721 (
            .O(N__17974),
            .I(N__17968));
    CascadeMux I__3720 (
            .O(N__17971),
            .I(N__17965));
    CascadeBuf I__3719 (
            .O(N__17968),
            .I(N__17962));
    CascadeBuf I__3718 (
            .O(N__17965),
            .I(N__17959));
    CascadeMux I__3717 (
            .O(N__17962),
            .I(N__17956));
    CascadeMux I__3716 (
            .O(N__17959),
            .I(N__17953));
    CascadeBuf I__3715 (
            .O(N__17956),
            .I(N__17950));
    CascadeBuf I__3714 (
            .O(N__17953),
            .I(N__17947));
    CascadeMux I__3713 (
            .O(N__17950),
            .I(N__17944));
    CascadeMux I__3712 (
            .O(N__17947),
            .I(N__17941));
    CascadeBuf I__3711 (
            .O(N__17944),
            .I(N__17938));
    CascadeBuf I__3710 (
            .O(N__17941),
            .I(N__17935));
    CascadeMux I__3709 (
            .O(N__17938),
            .I(N__17932));
    CascadeMux I__3708 (
            .O(N__17935),
            .I(N__17929));
    CascadeBuf I__3707 (
            .O(N__17932),
            .I(N__17926));
    CascadeBuf I__3706 (
            .O(N__17929),
            .I(N__17923));
    CascadeMux I__3705 (
            .O(N__17926),
            .I(N__17920));
    CascadeMux I__3704 (
            .O(N__17923),
            .I(N__17917));
    CascadeBuf I__3703 (
            .O(N__17920),
            .I(N__17914));
    CascadeBuf I__3702 (
            .O(N__17917),
            .I(N__17911));
    CascadeMux I__3701 (
            .O(N__17914),
            .I(N__17908));
    CascadeMux I__3700 (
            .O(N__17911),
            .I(N__17905));
    CascadeBuf I__3699 (
            .O(N__17908),
            .I(N__17902));
    CascadeBuf I__3698 (
            .O(N__17905),
            .I(N__17899));
    CascadeMux I__3697 (
            .O(N__17902),
            .I(N__17896));
    CascadeMux I__3696 (
            .O(N__17899),
            .I(N__17893));
    CascadeBuf I__3695 (
            .O(N__17896),
            .I(N__17890));
    CascadeBuf I__3694 (
            .O(N__17893),
            .I(N__17887));
    CascadeMux I__3693 (
            .O(N__17890),
            .I(N__17884));
    CascadeMux I__3692 (
            .O(N__17887),
            .I(N__17881));
    CascadeBuf I__3691 (
            .O(N__17884),
            .I(N__17878));
    CascadeBuf I__3690 (
            .O(N__17881),
            .I(N__17875));
    CascadeMux I__3689 (
            .O(N__17878),
            .I(N__17872));
    CascadeMux I__3688 (
            .O(N__17875),
            .I(N__17869));
    CascadeBuf I__3687 (
            .O(N__17872),
            .I(N__17866));
    CascadeBuf I__3686 (
            .O(N__17869),
            .I(N__17863));
    CascadeMux I__3685 (
            .O(N__17866),
            .I(N__17859));
    CascadeMux I__3684 (
            .O(N__17863),
            .I(N__17856));
    InMux I__3683 (
            .O(N__17862),
            .I(N__17853));
    InMux I__3682 (
            .O(N__17859),
            .I(N__17850));
    InMux I__3681 (
            .O(N__17856),
            .I(N__17847));
    LocalMux I__3680 (
            .O(N__17853),
            .I(N__17843));
    LocalMux I__3679 (
            .O(N__17850),
            .I(N__17840));
    LocalMux I__3678 (
            .O(N__17847),
            .I(N__17837));
    InMux I__3677 (
            .O(N__17846),
            .I(N__17834));
    Span12Mux_v I__3676 (
            .O(N__17843),
            .I(N__17827));
    Span12Mux_h I__3675 (
            .O(N__17840),
            .I(N__17827));
    Span12Mux_h I__3674 (
            .O(N__17837),
            .I(N__17827));
    LocalMux I__3673 (
            .O(N__17834),
            .I(RX_ADDR_3));
    Odrv12 I__3672 (
            .O(N__17827),
            .I(RX_ADDR_3));
    InMux I__3671 (
            .O(N__17822),
            .I(N__17819));
    LocalMux I__3670 (
            .O(N__17819),
            .I(N__17816));
    Span12Mux_s10_v I__3669 (
            .O(N__17816),
            .I(N__17813));
    Odrv12 I__3668 (
            .O(N__17813),
            .I(\receive_module.n127 ));
    CascadeMux I__3667 (
            .O(N__17810),
            .I(N__17807));
    CascadeBuf I__3666 (
            .O(N__17807),
            .I(N__17803));
    CascadeMux I__3665 (
            .O(N__17806),
            .I(N__17800));
    CascadeMux I__3664 (
            .O(N__17803),
            .I(N__17797));
    CascadeBuf I__3663 (
            .O(N__17800),
            .I(N__17794));
    CascadeBuf I__3662 (
            .O(N__17797),
            .I(N__17791));
    CascadeMux I__3661 (
            .O(N__17794),
            .I(N__17788));
    CascadeMux I__3660 (
            .O(N__17791),
            .I(N__17785));
    CascadeBuf I__3659 (
            .O(N__17788),
            .I(N__17782));
    CascadeBuf I__3658 (
            .O(N__17785),
            .I(N__17779));
    CascadeMux I__3657 (
            .O(N__17782),
            .I(N__17776));
    CascadeMux I__3656 (
            .O(N__17779),
            .I(N__17773));
    CascadeBuf I__3655 (
            .O(N__17776),
            .I(N__17770));
    CascadeBuf I__3654 (
            .O(N__17773),
            .I(N__17767));
    CascadeMux I__3653 (
            .O(N__17770),
            .I(N__17764));
    CascadeMux I__3652 (
            .O(N__17767),
            .I(N__17761));
    CascadeBuf I__3651 (
            .O(N__17764),
            .I(N__17758));
    CascadeBuf I__3650 (
            .O(N__17761),
            .I(N__17755));
    CascadeMux I__3649 (
            .O(N__17758),
            .I(N__17752));
    CascadeMux I__3648 (
            .O(N__17755),
            .I(N__17749));
    CascadeBuf I__3647 (
            .O(N__17752),
            .I(N__17746));
    CascadeBuf I__3646 (
            .O(N__17749),
            .I(N__17743));
    CascadeMux I__3645 (
            .O(N__17746),
            .I(N__17740));
    CascadeMux I__3644 (
            .O(N__17743),
            .I(N__17737));
    CascadeBuf I__3643 (
            .O(N__17740),
            .I(N__17734));
    CascadeBuf I__3642 (
            .O(N__17737),
            .I(N__17731));
    CascadeMux I__3641 (
            .O(N__17734),
            .I(N__17728));
    CascadeMux I__3640 (
            .O(N__17731),
            .I(N__17725));
    CascadeBuf I__3639 (
            .O(N__17728),
            .I(N__17722));
    CascadeBuf I__3638 (
            .O(N__17725),
            .I(N__17719));
    CascadeMux I__3637 (
            .O(N__17722),
            .I(N__17716));
    CascadeMux I__3636 (
            .O(N__17719),
            .I(N__17713));
    CascadeBuf I__3635 (
            .O(N__17716),
            .I(N__17710));
    CascadeBuf I__3634 (
            .O(N__17713),
            .I(N__17707));
    CascadeMux I__3633 (
            .O(N__17710),
            .I(N__17704));
    CascadeMux I__3632 (
            .O(N__17707),
            .I(N__17701));
    CascadeBuf I__3631 (
            .O(N__17704),
            .I(N__17698));
    CascadeBuf I__3630 (
            .O(N__17701),
            .I(N__17695));
    CascadeMux I__3629 (
            .O(N__17698),
            .I(N__17692));
    CascadeMux I__3628 (
            .O(N__17695),
            .I(N__17689));
    CascadeBuf I__3627 (
            .O(N__17692),
            .I(N__17686));
    CascadeBuf I__3626 (
            .O(N__17689),
            .I(N__17683));
    CascadeMux I__3625 (
            .O(N__17686),
            .I(N__17680));
    CascadeMux I__3624 (
            .O(N__17683),
            .I(N__17677));
    CascadeBuf I__3623 (
            .O(N__17680),
            .I(N__17674));
    CascadeBuf I__3622 (
            .O(N__17677),
            .I(N__17671));
    CascadeMux I__3621 (
            .O(N__17674),
            .I(N__17668));
    CascadeMux I__3620 (
            .O(N__17671),
            .I(N__17665));
    CascadeBuf I__3619 (
            .O(N__17668),
            .I(N__17662));
    CascadeBuf I__3618 (
            .O(N__17665),
            .I(N__17659));
    CascadeMux I__3617 (
            .O(N__17662),
            .I(N__17656));
    CascadeMux I__3616 (
            .O(N__17659),
            .I(N__17653));
    CascadeBuf I__3615 (
            .O(N__17656),
            .I(N__17650));
    CascadeBuf I__3614 (
            .O(N__17653),
            .I(N__17647));
    CascadeMux I__3613 (
            .O(N__17650),
            .I(N__17644));
    CascadeMux I__3612 (
            .O(N__17647),
            .I(N__17641));
    CascadeBuf I__3611 (
            .O(N__17644),
            .I(N__17638));
    CascadeBuf I__3610 (
            .O(N__17641),
            .I(N__17635));
    CascadeMux I__3609 (
            .O(N__17638),
            .I(N__17632));
    CascadeMux I__3608 (
            .O(N__17635),
            .I(N__17629));
    CascadeBuf I__3607 (
            .O(N__17632),
            .I(N__17626));
    InMux I__3606 (
            .O(N__17629),
            .I(N__17622));
    CascadeMux I__3605 (
            .O(N__17626),
            .I(N__17619));
    InMux I__3604 (
            .O(N__17625),
            .I(N__17616));
    LocalMux I__3603 (
            .O(N__17622),
            .I(N__17613));
    InMux I__3602 (
            .O(N__17619),
            .I(N__17610));
    LocalMux I__3601 (
            .O(N__17616),
            .I(N__17607));
    Span4Mux_s1_v I__3600 (
            .O(N__17613),
            .I(N__17604));
    LocalMux I__3599 (
            .O(N__17610),
            .I(N__17601));
    Span12Mux_v I__3598 (
            .O(N__17607),
            .I(N__17598));
    Span4Mux_h I__3597 (
            .O(N__17604),
            .I(N__17594));
    Span4Mux_s1_v I__3596 (
            .O(N__17601),
            .I(N__17591));
    Span12Mux_v I__3595 (
            .O(N__17598),
            .I(N__17588));
    InMux I__3594 (
            .O(N__17597),
            .I(N__17585));
    Span4Mux_h I__3593 (
            .O(N__17594),
            .I(N__17582));
    Span4Mux_h I__3592 (
            .O(N__17591),
            .I(N__17579));
    Odrv12 I__3591 (
            .O(N__17588),
            .I(RX_ADDR_10));
    LocalMux I__3590 (
            .O(N__17585),
            .I(RX_ADDR_10));
    Odrv4 I__3589 (
            .O(N__17582),
            .I(RX_ADDR_10));
    Odrv4 I__3588 (
            .O(N__17579),
            .I(RX_ADDR_10));
    SRMux I__3587 (
            .O(N__17570),
            .I(N__17567));
    LocalMux I__3586 (
            .O(N__17567),
            .I(N__17562));
    SRMux I__3585 (
            .O(N__17566),
            .I(N__17559));
    SRMux I__3584 (
            .O(N__17565),
            .I(N__17556));
    Span4Mux_v I__3583 (
            .O(N__17562),
            .I(N__17549));
    LocalMux I__3582 (
            .O(N__17559),
            .I(N__17549));
    LocalMux I__3581 (
            .O(N__17556),
            .I(N__17546));
    SRMux I__3580 (
            .O(N__17555),
            .I(N__17543));
    SRMux I__3579 (
            .O(N__17554),
            .I(N__17538));
    Span4Mux_v I__3578 (
            .O(N__17549),
            .I(N__17531));
    Span4Mux_v I__3577 (
            .O(N__17546),
            .I(N__17531));
    LocalMux I__3576 (
            .O(N__17543),
            .I(N__17531));
    SRMux I__3575 (
            .O(N__17542),
            .I(N__17528));
    SRMux I__3574 (
            .O(N__17541),
            .I(N__17525));
    LocalMux I__3573 (
            .O(N__17538),
            .I(N__17522));
    Span4Mux_v I__3572 (
            .O(N__17531),
            .I(N__17517));
    LocalMux I__3571 (
            .O(N__17528),
            .I(N__17517));
    LocalMux I__3570 (
            .O(N__17525),
            .I(N__17514));
    Span4Mux_h I__3569 (
            .O(N__17522),
            .I(N__17510));
    Span4Mux_v I__3568 (
            .O(N__17517),
            .I(N__17505));
    Span4Mux_h I__3567 (
            .O(N__17514),
            .I(N__17505));
    SRMux I__3566 (
            .O(N__17513),
            .I(N__17502));
    Odrv4 I__3565 (
            .O(N__17510),
            .I(\receive_module.n3677 ));
    Odrv4 I__3564 (
            .O(N__17505),
            .I(\receive_module.n3677 ));
    LocalMux I__3563 (
            .O(N__17502),
            .I(\receive_module.n3677 ));
    IoInMux I__3562 (
            .O(N__17495),
            .I(N__17492));
    LocalMux I__3561 (
            .O(N__17492),
            .I(N__17489));
    Span4Mux_s1_v I__3560 (
            .O(N__17489),
            .I(N__17486));
    Span4Mux_v I__3559 (
            .O(N__17486),
            .I(N__17483));
    Span4Mux_h I__3558 (
            .O(N__17483),
            .I(N__17480));
    Odrv4 I__3557 (
            .O(N__17480),
            .I(LED_c));
    InMux I__3556 (
            .O(N__17477),
            .I(N__17474));
    LocalMux I__3555 (
            .O(N__17474),
            .I(N__17470));
    InMux I__3554 (
            .O(N__17473),
            .I(N__17467));
    Odrv4 I__3553 (
            .O(N__17470),
            .I(PULSE_1HZ));
    LocalMux I__3552 (
            .O(N__17467),
            .I(PULSE_1HZ));
    InMux I__3551 (
            .O(N__17462),
            .I(N__17456));
    InMux I__3550 (
            .O(N__17461),
            .I(N__17456));
    LocalMux I__3549 (
            .O(N__17456),
            .I(\receive_module.rx_counter.old_VS ));
    InMux I__3548 (
            .O(N__17453),
            .I(N__17450));
    LocalMux I__3547 (
            .O(N__17450),
            .I(N__17447));
    Span4Mux_v I__3546 (
            .O(N__17447),
            .I(N__17444));
    Span4Mux_v I__3545 (
            .O(N__17444),
            .I(N__17441));
    Odrv4 I__3544 (
            .O(N__17441),
            .I(\receive_module.n133 ));
    CascadeMux I__3543 (
            .O(N__17438),
            .I(N__17434));
    CascadeMux I__3542 (
            .O(N__17437),
            .I(N__17431));
    CascadeBuf I__3541 (
            .O(N__17434),
            .I(N__17428));
    CascadeBuf I__3540 (
            .O(N__17431),
            .I(N__17425));
    CascadeMux I__3539 (
            .O(N__17428),
            .I(N__17422));
    CascadeMux I__3538 (
            .O(N__17425),
            .I(N__17419));
    CascadeBuf I__3537 (
            .O(N__17422),
            .I(N__17416));
    CascadeBuf I__3536 (
            .O(N__17419),
            .I(N__17413));
    CascadeMux I__3535 (
            .O(N__17416),
            .I(N__17410));
    CascadeMux I__3534 (
            .O(N__17413),
            .I(N__17407));
    CascadeBuf I__3533 (
            .O(N__17410),
            .I(N__17404));
    CascadeBuf I__3532 (
            .O(N__17407),
            .I(N__17401));
    CascadeMux I__3531 (
            .O(N__17404),
            .I(N__17398));
    CascadeMux I__3530 (
            .O(N__17401),
            .I(N__17395));
    CascadeBuf I__3529 (
            .O(N__17398),
            .I(N__17392));
    CascadeBuf I__3528 (
            .O(N__17395),
            .I(N__17389));
    CascadeMux I__3527 (
            .O(N__17392),
            .I(N__17386));
    CascadeMux I__3526 (
            .O(N__17389),
            .I(N__17383));
    CascadeBuf I__3525 (
            .O(N__17386),
            .I(N__17380));
    CascadeBuf I__3524 (
            .O(N__17383),
            .I(N__17377));
    CascadeMux I__3523 (
            .O(N__17380),
            .I(N__17374));
    CascadeMux I__3522 (
            .O(N__17377),
            .I(N__17371));
    CascadeBuf I__3521 (
            .O(N__17374),
            .I(N__17368));
    CascadeBuf I__3520 (
            .O(N__17371),
            .I(N__17365));
    CascadeMux I__3519 (
            .O(N__17368),
            .I(N__17362));
    CascadeMux I__3518 (
            .O(N__17365),
            .I(N__17359));
    CascadeBuf I__3517 (
            .O(N__17362),
            .I(N__17356));
    CascadeBuf I__3516 (
            .O(N__17359),
            .I(N__17353));
    CascadeMux I__3515 (
            .O(N__17356),
            .I(N__17350));
    CascadeMux I__3514 (
            .O(N__17353),
            .I(N__17347));
    CascadeBuf I__3513 (
            .O(N__17350),
            .I(N__17344));
    CascadeBuf I__3512 (
            .O(N__17347),
            .I(N__17341));
    CascadeMux I__3511 (
            .O(N__17344),
            .I(N__17338));
    CascadeMux I__3510 (
            .O(N__17341),
            .I(N__17335));
    CascadeBuf I__3509 (
            .O(N__17338),
            .I(N__17332));
    CascadeBuf I__3508 (
            .O(N__17335),
            .I(N__17329));
    CascadeMux I__3507 (
            .O(N__17332),
            .I(N__17326));
    CascadeMux I__3506 (
            .O(N__17329),
            .I(N__17323));
    CascadeBuf I__3505 (
            .O(N__17326),
            .I(N__17320));
    CascadeBuf I__3504 (
            .O(N__17323),
            .I(N__17317));
    CascadeMux I__3503 (
            .O(N__17320),
            .I(N__17314));
    CascadeMux I__3502 (
            .O(N__17317),
            .I(N__17311));
    CascadeBuf I__3501 (
            .O(N__17314),
            .I(N__17308));
    CascadeBuf I__3500 (
            .O(N__17311),
            .I(N__17305));
    CascadeMux I__3499 (
            .O(N__17308),
            .I(N__17302));
    CascadeMux I__3498 (
            .O(N__17305),
            .I(N__17299));
    CascadeBuf I__3497 (
            .O(N__17302),
            .I(N__17296));
    CascadeBuf I__3496 (
            .O(N__17299),
            .I(N__17293));
    CascadeMux I__3495 (
            .O(N__17296),
            .I(N__17290));
    CascadeMux I__3494 (
            .O(N__17293),
            .I(N__17287));
    CascadeBuf I__3493 (
            .O(N__17290),
            .I(N__17284));
    CascadeBuf I__3492 (
            .O(N__17287),
            .I(N__17281));
    CascadeMux I__3491 (
            .O(N__17284),
            .I(N__17278));
    CascadeMux I__3490 (
            .O(N__17281),
            .I(N__17275));
    CascadeBuf I__3489 (
            .O(N__17278),
            .I(N__17272));
    CascadeBuf I__3488 (
            .O(N__17275),
            .I(N__17269));
    CascadeMux I__3487 (
            .O(N__17272),
            .I(N__17266));
    CascadeMux I__3486 (
            .O(N__17269),
            .I(N__17263));
    CascadeBuf I__3485 (
            .O(N__17266),
            .I(N__17260));
    CascadeBuf I__3484 (
            .O(N__17263),
            .I(N__17257));
    CascadeMux I__3483 (
            .O(N__17260),
            .I(N__17254));
    CascadeMux I__3482 (
            .O(N__17257),
            .I(N__17251));
    InMux I__3481 (
            .O(N__17254),
            .I(N__17248));
    InMux I__3480 (
            .O(N__17251),
            .I(N__17245));
    LocalMux I__3479 (
            .O(N__17248),
            .I(N__17241));
    LocalMux I__3478 (
            .O(N__17245),
            .I(N__17238));
    InMux I__3477 (
            .O(N__17244),
            .I(N__17235));
    Span4Mux_s1_v I__3476 (
            .O(N__17241),
            .I(N__17232));
    Span4Mux_s1_v I__3475 (
            .O(N__17238),
            .I(N__17229));
    LocalMux I__3474 (
            .O(N__17235),
            .I(N__17226));
    Sp12to4 I__3473 (
            .O(N__17232),
            .I(N__17223));
    Sp12to4 I__3472 (
            .O(N__17229),
            .I(N__17220));
    Span4Mux_h I__3471 (
            .O(N__17226),
            .I(N__17216));
    Span12Mux_s6_h I__3470 (
            .O(N__17223),
            .I(N__17213));
    Span12Mux_s5_h I__3469 (
            .O(N__17220),
            .I(N__17210));
    InMux I__3468 (
            .O(N__17219),
            .I(N__17207));
    Span4Mux_v I__3467 (
            .O(N__17216),
            .I(N__17204));
    Span12Mux_v I__3466 (
            .O(N__17213),
            .I(N__17201));
    Span12Mux_v I__3465 (
            .O(N__17210),
            .I(N__17198));
    LocalMux I__3464 (
            .O(N__17207),
            .I(RX_ADDR_4));
    Odrv4 I__3463 (
            .O(N__17204),
            .I(RX_ADDR_4));
    Odrv12 I__3462 (
            .O(N__17201),
            .I(RX_ADDR_4));
    Odrv12 I__3461 (
            .O(N__17198),
            .I(RX_ADDR_4));
    InMux I__3460 (
            .O(N__17189),
            .I(N__17186));
    LocalMux I__3459 (
            .O(N__17186),
            .I(N__17183));
    Span12Mux_v I__3458 (
            .O(N__17183),
            .I(N__17180));
    Odrv12 I__3457 (
            .O(N__17180),
            .I(\receive_module.n132 ));
    CascadeMux I__3456 (
            .O(N__17177),
            .I(N__17173));
    CascadeMux I__3455 (
            .O(N__17176),
            .I(N__17170));
    CascadeBuf I__3454 (
            .O(N__17173),
            .I(N__17167));
    CascadeBuf I__3453 (
            .O(N__17170),
            .I(N__17164));
    CascadeMux I__3452 (
            .O(N__17167),
            .I(N__17161));
    CascadeMux I__3451 (
            .O(N__17164),
            .I(N__17158));
    CascadeBuf I__3450 (
            .O(N__17161),
            .I(N__17155));
    CascadeBuf I__3449 (
            .O(N__17158),
            .I(N__17152));
    CascadeMux I__3448 (
            .O(N__17155),
            .I(N__17149));
    CascadeMux I__3447 (
            .O(N__17152),
            .I(N__17146));
    CascadeBuf I__3446 (
            .O(N__17149),
            .I(N__17143));
    CascadeBuf I__3445 (
            .O(N__17146),
            .I(N__17140));
    CascadeMux I__3444 (
            .O(N__17143),
            .I(N__17137));
    CascadeMux I__3443 (
            .O(N__17140),
            .I(N__17134));
    CascadeBuf I__3442 (
            .O(N__17137),
            .I(N__17131));
    CascadeBuf I__3441 (
            .O(N__17134),
            .I(N__17128));
    CascadeMux I__3440 (
            .O(N__17131),
            .I(N__17125));
    CascadeMux I__3439 (
            .O(N__17128),
            .I(N__17122));
    CascadeBuf I__3438 (
            .O(N__17125),
            .I(N__17119));
    CascadeBuf I__3437 (
            .O(N__17122),
            .I(N__17116));
    CascadeMux I__3436 (
            .O(N__17119),
            .I(N__17113));
    CascadeMux I__3435 (
            .O(N__17116),
            .I(N__17110));
    CascadeBuf I__3434 (
            .O(N__17113),
            .I(N__17107));
    CascadeBuf I__3433 (
            .O(N__17110),
            .I(N__17104));
    CascadeMux I__3432 (
            .O(N__17107),
            .I(N__17101));
    CascadeMux I__3431 (
            .O(N__17104),
            .I(N__17098));
    CascadeBuf I__3430 (
            .O(N__17101),
            .I(N__17095));
    CascadeBuf I__3429 (
            .O(N__17098),
            .I(N__17092));
    CascadeMux I__3428 (
            .O(N__17095),
            .I(N__17089));
    CascadeMux I__3427 (
            .O(N__17092),
            .I(N__17086));
    CascadeBuf I__3426 (
            .O(N__17089),
            .I(N__17083));
    CascadeBuf I__3425 (
            .O(N__17086),
            .I(N__17080));
    CascadeMux I__3424 (
            .O(N__17083),
            .I(N__17077));
    CascadeMux I__3423 (
            .O(N__17080),
            .I(N__17074));
    CascadeBuf I__3422 (
            .O(N__17077),
            .I(N__17071));
    CascadeBuf I__3421 (
            .O(N__17074),
            .I(N__17068));
    CascadeMux I__3420 (
            .O(N__17071),
            .I(N__17065));
    CascadeMux I__3419 (
            .O(N__17068),
            .I(N__17062));
    CascadeBuf I__3418 (
            .O(N__17065),
            .I(N__17059));
    CascadeBuf I__3417 (
            .O(N__17062),
            .I(N__17056));
    CascadeMux I__3416 (
            .O(N__17059),
            .I(N__17053));
    CascadeMux I__3415 (
            .O(N__17056),
            .I(N__17050));
    CascadeBuf I__3414 (
            .O(N__17053),
            .I(N__17047));
    CascadeBuf I__3413 (
            .O(N__17050),
            .I(N__17044));
    CascadeMux I__3412 (
            .O(N__17047),
            .I(N__17041));
    CascadeMux I__3411 (
            .O(N__17044),
            .I(N__17038));
    CascadeBuf I__3410 (
            .O(N__17041),
            .I(N__17035));
    CascadeBuf I__3409 (
            .O(N__17038),
            .I(N__17032));
    CascadeMux I__3408 (
            .O(N__17035),
            .I(N__17029));
    CascadeMux I__3407 (
            .O(N__17032),
            .I(N__17026));
    CascadeBuf I__3406 (
            .O(N__17029),
            .I(N__17023));
    CascadeBuf I__3405 (
            .O(N__17026),
            .I(N__17020));
    CascadeMux I__3404 (
            .O(N__17023),
            .I(N__17017));
    CascadeMux I__3403 (
            .O(N__17020),
            .I(N__17014));
    CascadeBuf I__3402 (
            .O(N__17017),
            .I(N__17011));
    CascadeBuf I__3401 (
            .O(N__17014),
            .I(N__17008));
    CascadeMux I__3400 (
            .O(N__17011),
            .I(N__17005));
    CascadeMux I__3399 (
            .O(N__17008),
            .I(N__17002));
    CascadeBuf I__3398 (
            .O(N__17005),
            .I(N__16999));
    CascadeBuf I__3397 (
            .O(N__17002),
            .I(N__16996));
    CascadeMux I__3396 (
            .O(N__16999),
            .I(N__16993));
    CascadeMux I__3395 (
            .O(N__16996),
            .I(N__16989));
    InMux I__3394 (
            .O(N__16993),
            .I(N__16986));
    InMux I__3393 (
            .O(N__16992),
            .I(N__16983));
    InMux I__3392 (
            .O(N__16989),
            .I(N__16980));
    LocalMux I__3391 (
            .O(N__16986),
            .I(N__16977));
    LocalMux I__3390 (
            .O(N__16983),
            .I(N__16973));
    LocalMux I__3389 (
            .O(N__16980),
            .I(N__16970));
    Span4Mux_h I__3388 (
            .O(N__16977),
            .I(N__16967));
    CascadeMux I__3387 (
            .O(N__16976),
            .I(N__16964));
    Span4Mux_h I__3386 (
            .O(N__16973),
            .I(N__16961));
    Sp12to4 I__3385 (
            .O(N__16970),
            .I(N__16958));
    Sp12to4 I__3384 (
            .O(N__16967),
            .I(N__16955));
    InMux I__3383 (
            .O(N__16964),
            .I(N__16952));
    Span4Mux_v I__3382 (
            .O(N__16961),
            .I(N__16949));
    Span12Mux_v I__3381 (
            .O(N__16958),
            .I(N__16946));
    Span12Mux_v I__3380 (
            .O(N__16955),
            .I(N__16943));
    LocalMux I__3379 (
            .O(N__16952),
            .I(RX_ADDR_5));
    Odrv4 I__3378 (
            .O(N__16949),
            .I(RX_ADDR_5));
    Odrv12 I__3377 (
            .O(N__16946),
            .I(RX_ADDR_5));
    Odrv12 I__3376 (
            .O(N__16943),
            .I(RX_ADDR_5));
    InMux I__3375 (
            .O(N__16934),
            .I(N__16931));
    LocalMux I__3374 (
            .O(N__16931),
            .I(N__16928));
    Span4Mux_v I__3373 (
            .O(N__16928),
            .I(N__16925));
    Span4Mux_v I__3372 (
            .O(N__16925),
            .I(N__16922));
    Odrv4 I__3371 (
            .O(N__16922),
            .I(\receive_module.n131 ));
    CascadeMux I__3370 (
            .O(N__16919),
            .I(N__16915));
    CascadeMux I__3369 (
            .O(N__16918),
            .I(N__16912));
    CascadeBuf I__3368 (
            .O(N__16915),
            .I(N__16909));
    CascadeBuf I__3367 (
            .O(N__16912),
            .I(N__16906));
    CascadeMux I__3366 (
            .O(N__16909),
            .I(N__16903));
    CascadeMux I__3365 (
            .O(N__16906),
            .I(N__16900));
    CascadeBuf I__3364 (
            .O(N__16903),
            .I(N__16897));
    CascadeBuf I__3363 (
            .O(N__16900),
            .I(N__16894));
    CascadeMux I__3362 (
            .O(N__16897),
            .I(N__16891));
    CascadeMux I__3361 (
            .O(N__16894),
            .I(N__16888));
    CascadeBuf I__3360 (
            .O(N__16891),
            .I(N__16885));
    CascadeBuf I__3359 (
            .O(N__16888),
            .I(N__16882));
    CascadeMux I__3358 (
            .O(N__16885),
            .I(N__16879));
    CascadeMux I__3357 (
            .O(N__16882),
            .I(N__16876));
    CascadeBuf I__3356 (
            .O(N__16879),
            .I(N__16873));
    CascadeBuf I__3355 (
            .O(N__16876),
            .I(N__16870));
    CascadeMux I__3354 (
            .O(N__16873),
            .I(N__16867));
    CascadeMux I__3353 (
            .O(N__16870),
            .I(N__16864));
    CascadeBuf I__3352 (
            .O(N__16867),
            .I(N__16861));
    CascadeBuf I__3351 (
            .O(N__16864),
            .I(N__16858));
    CascadeMux I__3350 (
            .O(N__16861),
            .I(N__16855));
    CascadeMux I__3349 (
            .O(N__16858),
            .I(N__16852));
    CascadeBuf I__3348 (
            .O(N__16855),
            .I(N__16849));
    CascadeBuf I__3347 (
            .O(N__16852),
            .I(N__16846));
    CascadeMux I__3346 (
            .O(N__16849),
            .I(N__16843));
    CascadeMux I__3345 (
            .O(N__16846),
            .I(N__16840));
    CascadeBuf I__3344 (
            .O(N__16843),
            .I(N__16837));
    CascadeBuf I__3343 (
            .O(N__16840),
            .I(N__16834));
    CascadeMux I__3342 (
            .O(N__16837),
            .I(N__16831));
    CascadeMux I__3341 (
            .O(N__16834),
            .I(N__16828));
    CascadeBuf I__3340 (
            .O(N__16831),
            .I(N__16825));
    CascadeBuf I__3339 (
            .O(N__16828),
            .I(N__16822));
    CascadeMux I__3338 (
            .O(N__16825),
            .I(N__16819));
    CascadeMux I__3337 (
            .O(N__16822),
            .I(N__16816));
    CascadeBuf I__3336 (
            .O(N__16819),
            .I(N__16813));
    CascadeBuf I__3335 (
            .O(N__16816),
            .I(N__16810));
    CascadeMux I__3334 (
            .O(N__16813),
            .I(N__16807));
    CascadeMux I__3333 (
            .O(N__16810),
            .I(N__16804));
    CascadeBuf I__3332 (
            .O(N__16807),
            .I(N__16801));
    CascadeBuf I__3331 (
            .O(N__16804),
            .I(N__16798));
    CascadeMux I__3330 (
            .O(N__16801),
            .I(N__16795));
    CascadeMux I__3329 (
            .O(N__16798),
            .I(N__16792));
    CascadeBuf I__3328 (
            .O(N__16795),
            .I(N__16789));
    CascadeBuf I__3327 (
            .O(N__16792),
            .I(N__16786));
    CascadeMux I__3326 (
            .O(N__16789),
            .I(N__16783));
    CascadeMux I__3325 (
            .O(N__16786),
            .I(N__16780));
    CascadeBuf I__3324 (
            .O(N__16783),
            .I(N__16777));
    CascadeBuf I__3323 (
            .O(N__16780),
            .I(N__16774));
    CascadeMux I__3322 (
            .O(N__16777),
            .I(N__16771));
    CascadeMux I__3321 (
            .O(N__16774),
            .I(N__16768));
    CascadeBuf I__3320 (
            .O(N__16771),
            .I(N__16765));
    CascadeBuf I__3319 (
            .O(N__16768),
            .I(N__16762));
    CascadeMux I__3318 (
            .O(N__16765),
            .I(N__16759));
    CascadeMux I__3317 (
            .O(N__16762),
            .I(N__16756));
    CascadeBuf I__3316 (
            .O(N__16759),
            .I(N__16753));
    CascadeBuf I__3315 (
            .O(N__16756),
            .I(N__16750));
    CascadeMux I__3314 (
            .O(N__16753),
            .I(N__16747));
    CascadeMux I__3313 (
            .O(N__16750),
            .I(N__16744));
    CascadeBuf I__3312 (
            .O(N__16747),
            .I(N__16741));
    CascadeBuf I__3311 (
            .O(N__16744),
            .I(N__16738));
    CascadeMux I__3310 (
            .O(N__16741),
            .I(N__16735));
    CascadeMux I__3309 (
            .O(N__16738),
            .I(N__16732));
    InMux I__3308 (
            .O(N__16735),
            .I(N__16729));
    InMux I__3307 (
            .O(N__16732),
            .I(N__16726));
    LocalMux I__3306 (
            .O(N__16729),
            .I(N__16722));
    LocalMux I__3305 (
            .O(N__16726),
            .I(N__16719));
    InMux I__3304 (
            .O(N__16725),
            .I(N__16716));
    Span4Mux_s3_v I__3303 (
            .O(N__16722),
            .I(N__16713));
    Span4Mux_s1_v I__3302 (
            .O(N__16719),
            .I(N__16710));
    LocalMux I__3301 (
            .O(N__16716),
            .I(N__16707));
    Span4Mux_v I__3300 (
            .O(N__16713),
            .I(N__16704));
    Span4Mux_h I__3299 (
            .O(N__16710),
            .I(N__16701));
    Span4Mux_v I__3298 (
            .O(N__16707),
            .I(N__16697));
    Sp12to4 I__3297 (
            .O(N__16704),
            .I(N__16694));
    Sp12to4 I__3296 (
            .O(N__16701),
            .I(N__16691));
    InMux I__3295 (
            .O(N__16700),
            .I(N__16688));
    Sp12to4 I__3294 (
            .O(N__16697),
            .I(N__16683));
    Span12Mux_h I__3293 (
            .O(N__16694),
            .I(N__16683));
    Span12Mux_v I__3292 (
            .O(N__16691),
            .I(N__16680));
    LocalMux I__3291 (
            .O(N__16688),
            .I(RX_ADDR_6));
    Odrv12 I__3290 (
            .O(N__16683),
            .I(RX_ADDR_6));
    Odrv12 I__3289 (
            .O(N__16680),
            .I(RX_ADDR_6));
    InMux I__3288 (
            .O(N__16673),
            .I(N__16670));
    LocalMux I__3287 (
            .O(N__16670),
            .I(N__16667));
    Span4Mux_v I__3286 (
            .O(N__16667),
            .I(N__16664));
    Span4Mux_v I__3285 (
            .O(N__16664),
            .I(N__16661));
    Odrv4 I__3284 (
            .O(N__16661),
            .I(\receive_module.n130 ));
    CascadeMux I__3283 (
            .O(N__16658),
            .I(N__16654));
    CascadeMux I__3282 (
            .O(N__16657),
            .I(N__16651));
    CascadeBuf I__3281 (
            .O(N__16654),
            .I(N__16648));
    CascadeBuf I__3280 (
            .O(N__16651),
            .I(N__16645));
    CascadeMux I__3279 (
            .O(N__16648),
            .I(N__16642));
    CascadeMux I__3278 (
            .O(N__16645),
            .I(N__16639));
    CascadeBuf I__3277 (
            .O(N__16642),
            .I(N__16636));
    CascadeBuf I__3276 (
            .O(N__16639),
            .I(N__16633));
    CascadeMux I__3275 (
            .O(N__16636),
            .I(N__16630));
    CascadeMux I__3274 (
            .O(N__16633),
            .I(N__16627));
    CascadeBuf I__3273 (
            .O(N__16630),
            .I(N__16624));
    CascadeBuf I__3272 (
            .O(N__16627),
            .I(N__16621));
    CascadeMux I__3271 (
            .O(N__16624),
            .I(N__16618));
    CascadeMux I__3270 (
            .O(N__16621),
            .I(N__16615));
    CascadeBuf I__3269 (
            .O(N__16618),
            .I(N__16612));
    CascadeBuf I__3268 (
            .O(N__16615),
            .I(N__16609));
    CascadeMux I__3267 (
            .O(N__16612),
            .I(N__16606));
    CascadeMux I__3266 (
            .O(N__16609),
            .I(N__16603));
    CascadeBuf I__3265 (
            .O(N__16606),
            .I(N__16600));
    CascadeBuf I__3264 (
            .O(N__16603),
            .I(N__16597));
    CascadeMux I__3263 (
            .O(N__16600),
            .I(N__16594));
    CascadeMux I__3262 (
            .O(N__16597),
            .I(N__16591));
    CascadeBuf I__3261 (
            .O(N__16594),
            .I(N__16588));
    CascadeBuf I__3260 (
            .O(N__16591),
            .I(N__16585));
    CascadeMux I__3259 (
            .O(N__16588),
            .I(N__16582));
    CascadeMux I__3258 (
            .O(N__16585),
            .I(N__16579));
    CascadeBuf I__3257 (
            .O(N__16582),
            .I(N__16576));
    CascadeBuf I__3256 (
            .O(N__16579),
            .I(N__16573));
    CascadeMux I__3255 (
            .O(N__16576),
            .I(N__16570));
    CascadeMux I__3254 (
            .O(N__16573),
            .I(N__16567));
    CascadeBuf I__3253 (
            .O(N__16570),
            .I(N__16564));
    CascadeBuf I__3252 (
            .O(N__16567),
            .I(N__16561));
    CascadeMux I__3251 (
            .O(N__16564),
            .I(N__16558));
    CascadeMux I__3250 (
            .O(N__16561),
            .I(N__16555));
    CascadeBuf I__3249 (
            .O(N__16558),
            .I(N__16552));
    CascadeBuf I__3248 (
            .O(N__16555),
            .I(N__16549));
    CascadeMux I__3247 (
            .O(N__16552),
            .I(N__16546));
    CascadeMux I__3246 (
            .O(N__16549),
            .I(N__16543));
    CascadeBuf I__3245 (
            .O(N__16546),
            .I(N__16540));
    CascadeBuf I__3244 (
            .O(N__16543),
            .I(N__16537));
    CascadeMux I__3243 (
            .O(N__16540),
            .I(N__16534));
    CascadeMux I__3242 (
            .O(N__16537),
            .I(N__16531));
    CascadeBuf I__3241 (
            .O(N__16534),
            .I(N__16528));
    CascadeBuf I__3240 (
            .O(N__16531),
            .I(N__16525));
    CascadeMux I__3239 (
            .O(N__16528),
            .I(N__16522));
    CascadeMux I__3238 (
            .O(N__16525),
            .I(N__16519));
    CascadeBuf I__3237 (
            .O(N__16522),
            .I(N__16516));
    CascadeBuf I__3236 (
            .O(N__16519),
            .I(N__16513));
    CascadeMux I__3235 (
            .O(N__16516),
            .I(N__16510));
    CascadeMux I__3234 (
            .O(N__16513),
            .I(N__16507));
    CascadeBuf I__3233 (
            .O(N__16510),
            .I(N__16504));
    CascadeBuf I__3232 (
            .O(N__16507),
            .I(N__16501));
    CascadeMux I__3231 (
            .O(N__16504),
            .I(N__16498));
    CascadeMux I__3230 (
            .O(N__16501),
            .I(N__16495));
    CascadeBuf I__3229 (
            .O(N__16498),
            .I(N__16492));
    CascadeBuf I__3228 (
            .O(N__16495),
            .I(N__16489));
    CascadeMux I__3227 (
            .O(N__16492),
            .I(N__16486));
    CascadeMux I__3226 (
            .O(N__16489),
            .I(N__16483));
    CascadeBuf I__3225 (
            .O(N__16486),
            .I(N__16480));
    CascadeBuf I__3224 (
            .O(N__16483),
            .I(N__16477));
    CascadeMux I__3223 (
            .O(N__16480),
            .I(N__16474));
    CascadeMux I__3222 (
            .O(N__16477),
            .I(N__16471));
    InMux I__3221 (
            .O(N__16474),
            .I(N__16468));
    InMux I__3220 (
            .O(N__16471),
            .I(N__16465));
    LocalMux I__3219 (
            .O(N__16468),
            .I(N__16461));
    LocalMux I__3218 (
            .O(N__16465),
            .I(N__16458));
    InMux I__3217 (
            .O(N__16464),
            .I(N__16454));
    Span4Mux_h I__3216 (
            .O(N__16461),
            .I(N__16451));
    Span4Mux_h I__3215 (
            .O(N__16458),
            .I(N__16448));
    CascadeMux I__3214 (
            .O(N__16457),
            .I(N__16445));
    LocalMux I__3213 (
            .O(N__16454),
            .I(N__16442));
    Sp12to4 I__3212 (
            .O(N__16451),
            .I(N__16439));
    Sp12to4 I__3211 (
            .O(N__16448),
            .I(N__16436));
    InMux I__3210 (
            .O(N__16445),
            .I(N__16433));
    Span12Mux_v I__3209 (
            .O(N__16442),
            .I(N__16430));
    Span12Mux_v I__3208 (
            .O(N__16439),
            .I(N__16425));
    Span12Mux_v I__3207 (
            .O(N__16436),
            .I(N__16425));
    LocalMux I__3206 (
            .O(N__16433),
            .I(RX_ADDR_7));
    Odrv12 I__3205 (
            .O(N__16430),
            .I(RX_ADDR_7));
    Odrv12 I__3204 (
            .O(N__16425),
            .I(RX_ADDR_7));
    InMux I__3203 (
            .O(N__16418),
            .I(N__16415));
    LocalMux I__3202 (
            .O(N__16415),
            .I(N__16412));
    Odrv12 I__3201 (
            .O(N__16412),
            .I(\transmit_module.ADDR_Y_COMPONENT_3 ));
    InMux I__3200 (
            .O(N__16409),
            .I(N__16406));
    LocalMux I__3199 (
            .O(N__16406),
            .I(N__16401));
    InMux I__3198 (
            .O(N__16405),
            .I(N__16398));
    CascadeMux I__3197 (
            .O(N__16404),
            .I(N__16394));
    Span4Mux_v I__3196 (
            .O(N__16401),
            .I(N__16391));
    LocalMux I__3195 (
            .O(N__16398),
            .I(N__16388));
    InMux I__3194 (
            .O(N__16397),
            .I(N__16385));
    InMux I__3193 (
            .O(N__16394),
            .I(N__16382));
    Odrv4 I__3192 (
            .O(N__16391),
            .I(\transmit_module.TX_ADDR_3 ));
    Odrv12 I__3191 (
            .O(N__16388),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__3190 (
            .O(N__16385),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__3189 (
            .O(N__16382),
            .I(\transmit_module.TX_ADDR_3 ));
    InMux I__3188 (
            .O(N__16373),
            .I(N__16370));
    LocalMux I__3187 (
            .O(N__16370),
            .I(N__16367));
    Span12Mux_v I__3186 (
            .O(N__16367),
            .I(N__16364));
    Odrv12 I__3185 (
            .O(N__16364),
            .I(\receive_module.n128 ));
    CascadeMux I__3184 (
            .O(N__16361),
            .I(N__16358));
    CascadeBuf I__3183 (
            .O(N__16358),
            .I(N__16355));
    CascadeMux I__3182 (
            .O(N__16355),
            .I(N__16351));
    CascadeMux I__3181 (
            .O(N__16354),
            .I(N__16348));
    CascadeBuf I__3180 (
            .O(N__16351),
            .I(N__16345));
    CascadeBuf I__3179 (
            .O(N__16348),
            .I(N__16342));
    CascadeMux I__3178 (
            .O(N__16345),
            .I(N__16339));
    CascadeMux I__3177 (
            .O(N__16342),
            .I(N__16336));
    CascadeBuf I__3176 (
            .O(N__16339),
            .I(N__16333));
    CascadeBuf I__3175 (
            .O(N__16336),
            .I(N__16330));
    CascadeMux I__3174 (
            .O(N__16333),
            .I(N__16327));
    CascadeMux I__3173 (
            .O(N__16330),
            .I(N__16324));
    CascadeBuf I__3172 (
            .O(N__16327),
            .I(N__16321));
    CascadeBuf I__3171 (
            .O(N__16324),
            .I(N__16318));
    CascadeMux I__3170 (
            .O(N__16321),
            .I(N__16315));
    CascadeMux I__3169 (
            .O(N__16318),
            .I(N__16312));
    CascadeBuf I__3168 (
            .O(N__16315),
            .I(N__16309));
    CascadeBuf I__3167 (
            .O(N__16312),
            .I(N__16306));
    CascadeMux I__3166 (
            .O(N__16309),
            .I(N__16303));
    CascadeMux I__3165 (
            .O(N__16306),
            .I(N__16300));
    CascadeBuf I__3164 (
            .O(N__16303),
            .I(N__16297));
    CascadeBuf I__3163 (
            .O(N__16300),
            .I(N__16294));
    CascadeMux I__3162 (
            .O(N__16297),
            .I(N__16291));
    CascadeMux I__3161 (
            .O(N__16294),
            .I(N__16288));
    CascadeBuf I__3160 (
            .O(N__16291),
            .I(N__16285));
    CascadeBuf I__3159 (
            .O(N__16288),
            .I(N__16282));
    CascadeMux I__3158 (
            .O(N__16285),
            .I(N__16279));
    CascadeMux I__3157 (
            .O(N__16282),
            .I(N__16276));
    CascadeBuf I__3156 (
            .O(N__16279),
            .I(N__16273));
    CascadeBuf I__3155 (
            .O(N__16276),
            .I(N__16270));
    CascadeMux I__3154 (
            .O(N__16273),
            .I(N__16267));
    CascadeMux I__3153 (
            .O(N__16270),
            .I(N__16264));
    CascadeBuf I__3152 (
            .O(N__16267),
            .I(N__16261));
    CascadeBuf I__3151 (
            .O(N__16264),
            .I(N__16258));
    CascadeMux I__3150 (
            .O(N__16261),
            .I(N__16255));
    CascadeMux I__3149 (
            .O(N__16258),
            .I(N__16252));
    CascadeBuf I__3148 (
            .O(N__16255),
            .I(N__16249));
    CascadeBuf I__3147 (
            .O(N__16252),
            .I(N__16246));
    CascadeMux I__3146 (
            .O(N__16249),
            .I(N__16243));
    CascadeMux I__3145 (
            .O(N__16246),
            .I(N__16240));
    CascadeBuf I__3144 (
            .O(N__16243),
            .I(N__16237));
    CascadeBuf I__3143 (
            .O(N__16240),
            .I(N__16234));
    CascadeMux I__3142 (
            .O(N__16237),
            .I(N__16231));
    CascadeMux I__3141 (
            .O(N__16234),
            .I(N__16228));
    CascadeBuf I__3140 (
            .O(N__16231),
            .I(N__16225));
    CascadeBuf I__3139 (
            .O(N__16228),
            .I(N__16222));
    CascadeMux I__3138 (
            .O(N__16225),
            .I(N__16219));
    CascadeMux I__3137 (
            .O(N__16222),
            .I(N__16216));
    CascadeBuf I__3136 (
            .O(N__16219),
            .I(N__16213));
    CascadeBuf I__3135 (
            .O(N__16216),
            .I(N__16210));
    CascadeMux I__3134 (
            .O(N__16213),
            .I(N__16207));
    CascadeMux I__3133 (
            .O(N__16210),
            .I(N__16204));
    CascadeBuf I__3132 (
            .O(N__16207),
            .I(N__16201));
    CascadeBuf I__3131 (
            .O(N__16204),
            .I(N__16198));
    CascadeMux I__3130 (
            .O(N__16201),
            .I(N__16195));
    CascadeMux I__3129 (
            .O(N__16198),
            .I(N__16192));
    CascadeBuf I__3128 (
            .O(N__16195),
            .I(N__16189));
    CascadeBuf I__3127 (
            .O(N__16192),
            .I(N__16186));
    CascadeMux I__3126 (
            .O(N__16189),
            .I(N__16183));
    CascadeMux I__3125 (
            .O(N__16186),
            .I(N__16180));
    InMux I__3124 (
            .O(N__16183),
            .I(N__16177));
    CascadeBuf I__3123 (
            .O(N__16180),
            .I(N__16174));
    LocalMux I__3122 (
            .O(N__16177),
            .I(N__16170));
    CascadeMux I__3121 (
            .O(N__16174),
            .I(N__16167));
    InMux I__3120 (
            .O(N__16173),
            .I(N__16164));
    Span4Mux_h I__3119 (
            .O(N__16170),
            .I(N__16161));
    InMux I__3118 (
            .O(N__16167),
            .I(N__16158));
    LocalMux I__3117 (
            .O(N__16164),
            .I(N__16155));
    Span4Mux_h I__3116 (
            .O(N__16161),
            .I(N__16152));
    LocalMux I__3115 (
            .O(N__16158),
            .I(N__16149));
    Span4Mux_v I__3114 (
            .O(N__16155),
            .I(N__16146));
    Sp12to4 I__3113 (
            .O(N__16152),
            .I(N__16142));
    Sp12to4 I__3112 (
            .O(N__16149),
            .I(N__16139));
    Span4Mux_v I__3111 (
            .O(N__16146),
            .I(N__16136));
    InMux I__3110 (
            .O(N__16145),
            .I(N__16133));
    Span12Mux_s9_v I__3109 (
            .O(N__16142),
            .I(N__16128));
    Span12Mux_s9_v I__3108 (
            .O(N__16139),
            .I(N__16128));
    Odrv4 I__3107 (
            .O(N__16136),
            .I(RX_ADDR_9));
    LocalMux I__3106 (
            .O(N__16133),
            .I(RX_ADDR_9));
    Odrv12 I__3105 (
            .O(N__16128),
            .I(RX_ADDR_9));
    IoInMux I__3104 (
            .O(N__16121),
            .I(N__16117));
    IoInMux I__3103 (
            .O(N__16120),
            .I(N__16114));
    LocalMux I__3102 (
            .O(N__16117),
            .I(N__16111));
    LocalMux I__3101 (
            .O(N__16114),
            .I(N__16108));
    Span12Mux_s2_h I__3100 (
            .O(N__16111),
            .I(N__16105));
    IoSpan4Mux I__3099 (
            .O(N__16108),
            .I(N__16102));
    Span12Mux_v I__3098 (
            .O(N__16105),
            .I(N__16099));
    Span4Mux_s1_v I__3097 (
            .O(N__16102),
            .I(N__16096));
    Span12Mux_h I__3096 (
            .O(N__16099),
            .I(N__16093));
    Span4Mux_v I__3095 (
            .O(N__16096),
            .I(N__16090));
    Odrv12 I__3094 (
            .O(N__16093),
            .I(GB_BUFFER_DEBUG_c_3_c_THRU_CO));
    Odrv4 I__3093 (
            .O(N__16090),
            .I(GB_BUFFER_DEBUG_c_3_c_THRU_CO));
    IoInMux I__3092 (
            .O(N__16085),
            .I(N__16081));
    IoInMux I__3091 (
            .O(N__16084),
            .I(N__16078));
    LocalMux I__3090 (
            .O(N__16081),
            .I(N__16075));
    LocalMux I__3089 (
            .O(N__16078),
            .I(N__16071));
    IoSpan4Mux I__3088 (
            .O(N__16075),
            .I(N__16068));
    IoInMux I__3087 (
            .O(N__16074),
            .I(N__16065));
    IoSpan4Mux I__3086 (
            .O(N__16071),
            .I(N__16062));
    IoSpan4Mux I__3085 (
            .O(N__16068),
            .I(N__16057));
    LocalMux I__3084 (
            .O(N__16065),
            .I(N__16057));
    Span4Mux_s2_h I__3083 (
            .O(N__16062),
            .I(N__16054));
    IoSpan4Mux I__3082 (
            .O(N__16057),
            .I(N__16051));
    Sp12to4 I__3081 (
            .O(N__16054),
            .I(N__16048));
    Span4Mux_s3_v I__3080 (
            .O(N__16051),
            .I(N__16045));
    Span12Mux_h I__3079 (
            .O(N__16048),
            .I(N__16042));
    Span4Mux_v I__3078 (
            .O(N__16045),
            .I(N__16039));
    Odrv12 I__3077 (
            .O(N__16042),
            .I(n1821));
    Odrv4 I__3076 (
            .O(N__16039),
            .I(n1821));
    InMux I__3075 (
            .O(N__16034),
            .I(N__16031));
    LocalMux I__3074 (
            .O(N__16031),
            .I(N__16028));
    Span12Mux_v I__3073 (
            .O(N__16028),
            .I(N__16025));
    Odrv12 I__3072 (
            .O(N__16025),
            .I(\receive_module.n129 ));
    CascadeMux I__3071 (
            .O(N__16022),
            .I(N__16018));
    CascadeMux I__3070 (
            .O(N__16021),
            .I(N__16015));
    CascadeBuf I__3069 (
            .O(N__16018),
            .I(N__16012));
    CascadeBuf I__3068 (
            .O(N__16015),
            .I(N__16009));
    CascadeMux I__3067 (
            .O(N__16012),
            .I(N__16006));
    CascadeMux I__3066 (
            .O(N__16009),
            .I(N__16003));
    CascadeBuf I__3065 (
            .O(N__16006),
            .I(N__16000));
    CascadeBuf I__3064 (
            .O(N__16003),
            .I(N__15997));
    CascadeMux I__3063 (
            .O(N__16000),
            .I(N__15994));
    CascadeMux I__3062 (
            .O(N__15997),
            .I(N__15991));
    CascadeBuf I__3061 (
            .O(N__15994),
            .I(N__15988));
    CascadeBuf I__3060 (
            .O(N__15991),
            .I(N__15985));
    CascadeMux I__3059 (
            .O(N__15988),
            .I(N__15982));
    CascadeMux I__3058 (
            .O(N__15985),
            .I(N__15979));
    CascadeBuf I__3057 (
            .O(N__15982),
            .I(N__15976));
    CascadeBuf I__3056 (
            .O(N__15979),
            .I(N__15973));
    CascadeMux I__3055 (
            .O(N__15976),
            .I(N__15970));
    CascadeMux I__3054 (
            .O(N__15973),
            .I(N__15967));
    CascadeBuf I__3053 (
            .O(N__15970),
            .I(N__15964));
    CascadeBuf I__3052 (
            .O(N__15967),
            .I(N__15961));
    CascadeMux I__3051 (
            .O(N__15964),
            .I(N__15958));
    CascadeMux I__3050 (
            .O(N__15961),
            .I(N__15955));
    CascadeBuf I__3049 (
            .O(N__15958),
            .I(N__15952));
    CascadeBuf I__3048 (
            .O(N__15955),
            .I(N__15949));
    CascadeMux I__3047 (
            .O(N__15952),
            .I(N__15946));
    CascadeMux I__3046 (
            .O(N__15949),
            .I(N__15943));
    CascadeBuf I__3045 (
            .O(N__15946),
            .I(N__15940));
    CascadeBuf I__3044 (
            .O(N__15943),
            .I(N__15937));
    CascadeMux I__3043 (
            .O(N__15940),
            .I(N__15934));
    CascadeMux I__3042 (
            .O(N__15937),
            .I(N__15931));
    CascadeBuf I__3041 (
            .O(N__15934),
            .I(N__15928));
    CascadeBuf I__3040 (
            .O(N__15931),
            .I(N__15925));
    CascadeMux I__3039 (
            .O(N__15928),
            .I(N__15922));
    CascadeMux I__3038 (
            .O(N__15925),
            .I(N__15919));
    CascadeBuf I__3037 (
            .O(N__15922),
            .I(N__15916));
    CascadeBuf I__3036 (
            .O(N__15919),
            .I(N__15913));
    CascadeMux I__3035 (
            .O(N__15916),
            .I(N__15910));
    CascadeMux I__3034 (
            .O(N__15913),
            .I(N__15907));
    CascadeBuf I__3033 (
            .O(N__15910),
            .I(N__15904));
    CascadeBuf I__3032 (
            .O(N__15907),
            .I(N__15901));
    CascadeMux I__3031 (
            .O(N__15904),
            .I(N__15898));
    CascadeMux I__3030 (
            .O(N__15901),
            .I(N__15895));
    CascadeBuf I__3029 (
            .O(N__15898),
            .I(N__15892));
    CascadeBuf I__3028 (
            .O(N__15895),
            .I(N__15889));
    CascadeMux I__3027 (
            .O(N__15892),
            .I(N__15886));
    CascadeMux I__3026 (
            .O(N__15889),
            .I(N__15883));
    CascadeBuf I__3025 (
            .O(N__15886),
            .I(N__15880));
    CascadeBuf I__3024 (
            .O(N__15883),
            .I(N__15877));
    CascadeMux I__3023 (
            .O(N__15880),
            .I(N__15874));
    CascadeMux I__3022 (
            .O(N__15877),
            .I(N__15871));
    CascadeBuf I__3021 (
            .O(N__15874),
            .I(N__15868));
    CascadeBuf I__3020 (
            .O(N__15871),
            .I(N__15865));
    CascadeMux I__3019 (
            .O(N__15868),
            .I(N__15862));
    CascadeMux I__3018 (
            .O(N__15865),
            .I(N__15859));
    CascadeBuf I__3017 (
            .O(N__15862),
            .I(N__15856));
    CascadeBuf I__3016 (
            .O(N__15859),
            .I(N__15853));
    CascadeMux I__3015 (
            .O(N__15856),
            .I(N__15850));
    CascadeMux I__3014 (
            .O(N__15853),
            .I(N__15847));
    CascadeBuf I__3013 (
            .O(N__15850),
            .I(N__15844));
    CascadeBuf I__3012 (
            .O(N__15847),
            .I(N__15841));
    CascadeMux I__3011 (
            .O(N__15844),
            .I(N__15838));
    CascadeMux I__3010 (
            .O(N__15841),
            .I(N__15835));
    InMux I__3009 (
            .O(N__15838),
            .I(N__15832));
    InMux I__3008 (
            .O(N__15835),
            .I(N__15829));
    LocalMux I__3007 (
            .O(N__15832),
            .I(N__15825));
    LocalMux I__3006 (
            .O(N__15829),
            .I(N__15822));
    InMux I__3005 (
            .O(N__15828),
            .I(N__15819));
    Span4Mux_s1_v I__3004 (
            .O(N__15825),
            .I(N__15816));
    Span4Mux_s1_v I__3003 (
            .O(N__15822),
            .I(N__15813));
    LocalMux I__3002 (
            .O(N__15819),
            .I(N__15809));
    Sp12to4 I__3001 (
            .O(N__15816),
            .I(N__15806));
    Span4Mux_h I__3000 (
            .O(N__15813),
            .I(N__15803));
    InMux I__2999 (
            .O(N__15812),
            .I(N__15800));
    Span12Mux_v I__2998 (
            .O(N__15809),
            .I(N__15795));
    Span12Mux_h I__2997 (
            .O(N__15806),
            .I(N__15795));
    Span4Mux_v I__2996 (
            .O(N__15803),
            .I(N__15792));
    LocalMux I__2995 (
            .O(N__15800),
            .I(RX_ADDR_8));
    Odrv12 I__2994 (
            .O(N__15795),
            .I(RX_ADDR_8));
    Odrv4 I__2993 (
            .O(N__15792),
            .I(RX_ADDR_8));
    CascadeMux I__2992 (
            .O(N__15785),
            .I(\transmit_module.n145_cascade_ ));
    InMux I__2991 (
            .O(N__15782),
            .I(N__15779));
    LocalMux I__2990 (
            .O(N__15779),
            .I(\transmit_module.Y_DELTA_PATTERN_2 ));
    InMux I__2989 (
            .O(N__15776),
            .I(N__15773));
    LocalMux I__2988 (
            .O(N__15773),
            .I(N__15770));
    Odrv12 I__2987 (
            .O(N__15770),
            .I(\transmit_module.Y_DELTA_PATTERN_5 ));
    InMux I__2986 (
            .O(N__15767),
            .I(N__15764));
    LocalMux I__2985 (
            .O(N__15764),
            .I(\transmit_module.Y_DELTA_PATTERN_4 ));
    InMux I__2984 (
            .O(N__15761),
            .I(N__15758));
    LocalMux I__2983 (
            .O(N__15758),
            .I(\transmit_module.Y_DELTA_PATTERN_3 ));
    InMux I__2982 (
            .O(N__15755),
            .I(N__15752));
    LocalMux I__2981 (
            .O(N__15752),
            .I(\transmit_module.Y_DELTA_PATTERN_1 ));
    InMux I__2980 (
            .O(N__15749),
            .I(N__15746));
    LocalMux I__2979 (
            .O(N__15746),
            .I(N__15743));
    Span4Mux_v I__2978 (
            .O(N__15743),
            .I(N__15740));
    Span4Mux_v I__2977 (
            .O(N__15740),
            .I(N__15737));
    Odrv4 I__2976 (
            .O(N__15737),
            .I(\receive_module.n136 ));
    CascadeMux I__2975 (
            .O(N__15734),
            .I(N__15730));
    CascadeMux I__2974 (
            .O(N__15733),
            .I(N__15727));
    CascadeBuf I__2973 (
            .O(N__15730),
            .I(N__15724));
    CascadeBuf I__2972 (
            .O(N__15727),
            .I(N__15721));
    CascadeMux I__2971 (
            .O(N__15724),
            .I(N__15718));
    CascadeMux I__2970 (
            .O(N__15721),
            .I(N__15715));
    CascadeBuf I__2969 (
            .O(N__15718),
            .I(N__15712));
    CascadeBuf I__2968 (
            .O(N__15715),
            .I(N__15709));
    CascadeMux I__2967 (
            .O(N__15712),
            .I(N__15706));
    CascadeMux I__2966 (
            .O(N__15709),
            .I(N__15703));
    CascadeBuf I__2965 (
            .O(N__15706),
            .I(N__15700));
    CascadeBuf I__2964 (
            .O(N__15703),
            .I(N__15697));
    CascadeMux I__2963 (
            .O(N__15700),
            .I(N__15694));
    CascadeMux I__2962 (
            .O(N__15697),
            .I(N__15691));
    CascadeBuf I__2961 (
            .O(N__15694),
            .I(N__15688));
    CascadeBuf I__2960 (
            .O(N__15691),
            .I(N__15685));
    CascadeMux I__2959 (
            .O(N__15688),
            .I(N__15682));
    CascadeMux I__2958 (
            .O(N__15685),
            .I(N__15679));
    CascadeBuf I__2957 (
            .O(N__15682),
            .I(N__15676));
    CascadeBuf I__2956 (
            .O(N__15679),
            .I(N__15673));
    CascadeMux I__2955 (
            .O(N__15676),
            .I(N__15670));
    CascadeMux I__2954 (
            .O(N__15673),
            .I(N__15667));
    CascadeBuf I__2953 (
            .O(N__15670),
            .I(N__15664));
    CascadeBuf I__2952 (
            .O(N__15667),
            .I(N__15661));
    CascadeMux I__2951 (
            .O(N__15664),
            .I(N__15658));
    CascadeMux I__2950 (
            .O(N__15661),
            .I(N__15655));
    CascadeBuf I__2949 (
            .O(N__15658),
            .I(N__15652));
    CascadeBuf I__2948 (
            .O(N__15655),
            .I(N__15649));
    CascadeMux I__2947 (
            .O(N__15652),
            .I(N__15646));
    CascadeMux I__2946 (
            .O(N__15649),
            .I(N__15643));
    CascadeBuf I__2945 (
            .O(N__15646),
            .I(N__15640));
    CascadeBuf I__2944 (
            .O(N__15643),
            .I(N__15637));
    CascadeMux I__2943 (
            .O(N__15640),
            .I(N__15634));
    CascadeMux I__2942 (
            .O(N__15637),
            .I(N__15631));
    CascadeBuf I__2941 (
            .O(N__15634),
            .I(N__15628));
    CascadeBuf I__2940 (
            .O(N__15631),
            .I(N__15625));
    CascadeMux I__2939 (
            .O(N__15628),
            .I(N__15622));
    CascadeMux I__2938 (
            .O(N__15625),
            .I(N__15619));
    CascadeBuf I__2937 (
            .O(N__15622),
            .I(N__15616));
    CascadeBuf I__2936 (
            .O(N__15619),
            .I(N__15613));
    CascadeMux I__2935 (
            .O(N__15616),
            .I(N__15610));
    CascadeMux I__2934 (
            .O(N__15613),
            .I(N__15607));
    CascadeBuf I__2933 (
            .O(N__15610),
            .I(N__15604));
    CascadeBuf I__2932 (
            .O(N__15607),
            .I(N__15601));
    CascadeMux I__2931 (
            .O(N__15604),
            .I(N__15598));
    CascadeMux I__2930 (
            .O(N__15601),
            .I(N__15595));
    CascadeBuf I__2929 (
            .O(N__15598),
            .I(N__15592));
    CascadeBuf I__2928 (
            .O(N__15595),
            .I(N__15589));
    CascadeMux I__2927 (
            .O(N__15592),
            .I(N__15586));
    CascadeMux I__2926 (
            .O(N__15589),
            .I(N__15583));
    CascadeBuf I__2925 (
            .O(N__15586),
            .I(N__15580));
    CascadeBuf I__2924 (
            .O(N__15583),
            .I(N__15577));
    CascadeMux I__2923 (
            .O(N__15580),
            .I(N__15574));
    CascadeMux I__2922 (
            .O(N__15577),
            .I(N__15571));
    CascadeBuf I__2921 (
            .O(N__15574),
            .I(N__15568));
    CascadeBuf I__2920 (
            .O(N__15571),
            .I(N__15565));
    CascadeMux I__2919 (
            .O(N__15568),
            .I(N__15562));
    CascadeMux I__2918 (
            .O(N__15565),
            .I(N__15559));
    CascadeBuf I__2917 (
            .O(N__15562),
            .I(N__15556));
    CascadeBuf I__2916 (
            .O(N__15559),
            .I(N__15553));
    CascadeMux I__2915 (
            .O(N__15556),
            .I(N__15550));
    CascadeMux I__2914 (
            .O(N__15553),
            .I(N__15547));
    InMux I__2913 (
            .O(N__15550),
            .I(N__15544));
    InMux I__2912 (
            .O(N__15547),
            .I(N__15541));
    LocalMux I__2911 (
            .O(N__15544),
            .I(N__15537));
    LocalMux I__2910 (
            .O(N__15541),
            .I(N__15534));
    InMux I__2909 (
            .O(N__15540),
            .I(N__15531));
    Span4Mux_s1_v I__2908 (
            .O(N__15537),
            .I(N__15528));
    Span4Mux_s1_v I__2907 (
            .O(N__15534),
            .I(N__15525));
    LocalMux I__2906 (
            .O(N__15531),
            .I(N__15522));
    Span4Mux_v I__2905 (
            .O(N__15528),
            .I(N__15519));
    Span4Mux_v I__2904 (
            .O(N__15525),
            .I(N__15516));
    Span4Mux_v I__2903 (
            .O(N__15522),
            .I(N__15512));
    Sp12to4 I__2902 (
            .O(N__15519),
            .I(N__15509));
    Sp12to4 I__2901 (
            .O(N__15516),
            .I(N__15506));
    InMux I__2900 (
            .O(N__15515),
            .I(N__15503));
    Sp12to4 I__2899 (
            .O(N__15512),
            .I(N__15496));
    Span12Mux_h I__2898 (
            .O(N__15509),
            .I(N__15496));
    Span12Mux_h I__2897 (
            .O(N__15506),
            .I(N__15496));
    LocalMux I__2896 (
            .O(N__15503),
            .I(RX_ADDR_1));
    Odrv12 I__2895 (
            .O(N__15496),
            .I(RX_ADDR_1));
    InMux I__2894 (
            .O(N__15491),
            .I(N__15488));
    LocalMux I__2893 (
            .O(N__15488),
            .I(N__15485));
    Odrv12 I__2892 (
            .O(N__15485),
            .I(\receive_module.n135 ));
    CascadeMux I__2891 (
            .O(N__15482),
            .I(N__15478));
    CascadeMux I__2890 (
            .O(N__15481),
            .I(N__15475));
    CascadeBuf I__2889 (
            .O(N__15478),
            .I(N__15472));
    CascadeBuf I__2888 (
            .O(N__15475),
            .I(N__15469));
    CascadeMux I__2887 (
            .O(N__15472),
            .I(N__15466));
    CascadeMux I__2886 (
            .O(N__15469),
            .I(N__15463));
    CascadeBuf I__2885 (
            .O(N__15466),
            .I(N__15460));
    CascadeBuf I__2884 (
            .O(N__15463),
            .I(N__15457));
    CascadeMux I__2883 (
            .O(N__15460),
            .I(N__15454));
    CascadeMux I__2882 (
            .O(N__15457),
            .I(N__15451));
    CascadeBuf I__2881 (
            .O(N__15454),
            .I(N__15448));
    CascadeBuf I__2880 (
            .O(N__15451),
            .I(N__15445));
    CascadeMux I__2879 (
            .O(N__15448),
            .I(N__15442));
    CascadeMux I__2878 (
            .O(N__15445),
            .I(N__15439));
    CascadeBuf I__2877 (
            .O(N__15442),
            .I(N__15436));
    CascadeBuf I__2876 (
            .O(N__15439),
            .I(N__15433));
    CascadeMux I__2875 (
            .O(N__15436),
            .I(N__15430));
    CascadeMux I__2874 (
            .O(N__15433),
            .I(N__15427));
    CascadeBuf I__2873 (
            .O(N__15430),
            .I(N__15424));
    CascadeBuf I__2872 (
            .O(N__15427),
            .I(N__15421));
    CascadeMux I__2871 (
            .O(N__15424),
            .I(N__15418));
    CascadeMux I__2870 (
            .O(N__15421),
            .I(N__15415));
    CascadeBuf I__2869 (
            .O(N__15418),
            .I(N__15412));
    CascadeBuf I__2868 (
            .O(N__15415),
            .I(N__15409));
    CascadeMux I__2867 (
            .O(N__15412),
            .I(N__15406));
    CascadeMux I__2866 (
            .O(N__15409),
            .I(N__15403));
    CascadeBuf I__2865 (
            .O(N__15406),
            .I(N__15400));
    CascadeBuf I__2864 (
            .O(N__15403),
            .I(N__15397));
    CascadeMux I__2863 (
            .O(N__15400),
            .I(N__15394));
    CascadeMux I__2862 (
            .O(N__15397),
            .I(N__15391));
    CascadeBuf I__2861 (
            .O(N__15394),
            .I(N__15388));
    CascadeBuf I__2860 (
            .O(N__15391),
            .I(N__15385));
    CascadeMux I__2859 (
            .O(N__15388),
            .I(N__15382));
    CascadeMux I__2858 (
            .O(N__15385),
            .I(N__15379));
    CascadeBuf I__2857 (
            .O(N__15382),
            .I(N__15376));
    CascadeBuf I__2856 (
            .O(N__15379),
            .I(N__15373));
    CascadeMux I__2855 (
            .O(N__15376),
            .I(N__15370));
    CascadeMux I__2854 (
            .O(N__15373),
            .I(N__15367));
    CascadeBuf I__2853 (
            .O(N__15370),
            .I(N__15364));
    CascadeBuf I__2852 (
            .O(N__15367),
            .I(N__15361));
    CascadeMux I__2851 (
            .O(N__15364),
            .I(N__15358));
    CascadeMux I__2850 (
            .O(N__15361),
            .I(N__15355));
    CascadeBuf I__2849 (
            .O(N__15358),
            .I(N__15352));
    CascadeBuf I__2848 (
            .O(N__15355),
            .I(N__15349));
    CascadeMux I__2847 (
            .O(N__15352),
            .I(N__15346));
    CascadeMux I__2846 (
            .O(N__15349),
            .I(N__15343));
    CascadeBuf I__2845 (
            .O(N__15346),
            .I(N__15340));
    CascadeBuf I__2844 (
            .O(N__15343),
            .I(N__15337));
    CascadeMux I__2843 (
            .O(N__15340),
            .I(N__15334));
    CascadeMux I__2842 (
            .O(N__15337),
            .I(N__15331));
    CascadeBuf I__2841 (
            .O(N__15334),
            .I(N__15328));
    CascadeBuf I__2840 (
            .O(N__15331),
            .I(N__15325));
    CascadeMux I__2839 (
            .O(N__15328),
            .I(N__15322));
    CascadeMux I__2838 (
            .O(N__15325),
            .I(N__15319));
    CascadeBuf I__2837 (
            .O(N__15322),
            .I(N__15316));
    CascadeBuf I__2836 (
            .O(N__15319),
            .I(N__15313));
    CascadeMux I__2835 (
            .O(N__15316),
            .I(N__15310));
    CascadeMux I__2834 (
            .O(N__15313),
            .I(N__15307));
    CascadeBuf I__2833 (
            .O(N__15310),
            .I(N__15304));
    CascadeBuf I__2832 (
            .O(N__15307),
            .I(N__15301));
    CascadeMux I__2831 (
            .O(N__15304),
            .I(N__15298));
    CascadeMux I__2830 (
            .O(N__15301),
            .I(N__15295));
    InMux I__2829 (
            .O(N__15298),
            .I(N__15292));
    InMux I__2828 (
            .O(N__15295),
            .I(N__15289));
    LocalMux I__2827 (
            .O(N__15292),
            .I(N__15285));
    LocalMux I__2826 (
            .O(N__15289),
            .I(N__15282));
    InMux I__2825 (
            .O(N__15288),
            .I(N__15279));
    Span4Mux_s3_v I__2824 (
            .O(N__15285),
            .I(N__15276));
    Span4Mux_s3_v I__2823 (
            .O(N__15282),
            .I(N__15273));
    LocalMux I__2822 (
            .O(N__15279),
            .I(N__15269));
    Sp12to4 I__2821 (
            .O(N__15276),
            .I(N__15266));
    Sp12to4 I__2820 (
            .O(N__15273),
            .I(N__15263));
    InMux I__2819 (
            .O(N__15272),
            .I(N__15260));
    Span12Mux_v I__2818 (
            .O(N__15269),
            .I(N__15255));
    Span12Mux_h I__2817 (
            .O(N__15266),
            .I(N__15255));
    Span12Mux_v I__2816 (
            .O(N__15263),
            .I(N__15252));
    LocalMux I__2815 (
            .O(N__15260),
            .I(RX_ADDR_2));
    Odrv12 I__2814 (
            .O(N__15255),
            .I(RX_ADDR_2));
    Odrv12 I__2813 (
            .O(N__15252),
            .I(RX_ADDR_2));
    InMux I__2812 (
            .O(N__15245),
            .I(N__15242));
    LocalMux I__2811 (
            .O(N__15242),
            .I(\transmit_module.X_DELTA_PATTERN_1 ));
    InMux I__2810 (
            .O(N__15239),
            .I(N__15236));
    LocalMux I__2809 (
            .O(N__15236),
            .I(N__15233));
    Odrv12 I__2808 (
            .O(N__15233),
            .I(\transmit_module.X_DELTA_PATTERN_8 ));
    InMux I__2807 (
            .O(N__15230),
            .I(N__15227));
    LocalMux I__2806 (
            .O(N__15227),
            .I(\transmit_module.X_DELTA_PATTERN_2 ));
    InMux I__2805 (
            .O(N__15224),
            .I(N__15221));
    LocalMux I__2804 (
            .O(N__15221),
            .I(\transmit_module.X_DELTA_PATTERN_3 ));
    InMux I__2803 (
            .O(N__15218),
            .I(N__15215));
    LocalMux I__2802 (
            .O(N__15215),
            .I(\transmit_module.X_DELTA_PATTERN_7 ));
    InMux I__2801 (
            .O(N__15212),
            .I(N__15209));
    LocalMux I__2800 (
            .O(N__15209),
            .I(\transmit_module.X_DELTA_PATTERN_4 ));
    InMux I__2799 (
            .O(N__15206),
            .I(N__15203));
    LocalMux I__2798 (
            .O(N__15203),
            .I(\transmit_module.n129 ));
    InMux I__2797 (
            .O(N__15200),
            .I(N__15196));
    InMux I__2796 (
            .O(N__15199),
            .I(N__15193));
    LocalMux I__2795 (
            .O(N__15196),
            .I(\transmit_module.n110 ));
    LocalMux I__2794 (
            .O(N__15193),
            .I(\transmit_module.n110 ));
    InMux I__2793 (
            .O(N__15188),
            .I(N__15185));
    LocalMux I__2792 (
            .O(N__15185),
            .I(N__15182));
    Odrv4 I__2791 (
            .O(N__15182),
            .I(\transmit_module.n141 ));
    InMux I__2790 (
            .O(N__15179),
            .I(N__15176));
    LocalMux I__2789 (
            .O(N__15176),
            .I(N__15170));
    InMux I__2788 (
            .O(N__15175),
            .I(N__15167));
    CascadeMux I__2787 (
            .O(N__15174),
            .I(N__15164));
    InMux I__2786 (
            .O(N__15173),
            .I(N__15161));
    Span4Mux_v I__2785 (
            .O(N__15170),
            .I(N__15156));
    LocalMux I__2784 (
            .O(N__15167),
            .I(N__15156));
    InMux I__2783 (
            .O(N__15164),
            .I(N__15153));
    LocalMux I__2782 (
            .O(N__15161),
            .I(\transmit_module.TX_ADDR_6 ));
    Odrv4 I__2781 (
            .O(N__15156),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__2780 (
            .O(N__15153),
            .I(\transmit_module.TX_ADDR_6 ));
    InMux I__2779 (
            .O(N__15146),
            .I(N__15137));
    InMux I__2778 (
            .O(N__15145),
            .I(N__15134));
    InMux I__2777 (
            .O(N__15144),
            .I(N__15131));
    CascadeMux I__2776 (
            .O(N__15143),
            .I(N__15128));
    InMux I__2775 (
            .O(N__15142),
            .I(N__15123));
    InMux I__2774 (
            .O(N__15141),
            .I(N__15120));
    InMux I__2773 (
            .O(N__15140),
            .I(N__15116));
    LocalMux I__2772 (
            .O(N__15137),
            .I(N__15111));
    LocalMux I__2771 (
            .O(N__15134),
            .I(N__15106));
    LocalMux I__2770 (
            .O(N__15131),
            .I(N__15106));
    InMux I__2769 (
            .O(N__15128),
            .I(N__15103));
    InMux I__2768 (
            .O(N__15127),
            .I(N__15098));
    InMux I__2767 (
            .O(N__15126),
            .I(N__15098));
    LocalMux I__2766 (
            .O(N__15123),
            .I(N__15093));
    LocalMux I__2765 (
            .O(N__15120),
            .I(N__15090));
    InMux I__2764 (
            .O(N__15119),
            .I(N__15087));
    LocalMux I__2763 (
            .O(N__15116),
            .I(N__15084));
    InMux I__2762 (
            .O(N__15115),
            .I(N__15081));
    InMux I__2761 (
            .O(N__15114),
            .I(N__15078));
    Span4Mux_h I__2760 (
            .O(N__15111),
            .I(N__15069));
    Span4Mux_v I__2759 (
            .O(N__15106),
            .I(N__15069));
    LocalMux I__2758 (
            .O(N__15103),
            .I(N__15069));
    LocalMux I__2757 (
            .O(N__15098),
            .I(N__15069));
    InMux I__2756 (
            .O(N__15097),
            .I(N__15066));
    InMux I__2755 (
            .O(N__15096),
            .I(N__15063));
    Odrv4 I__2754 (
            .O(N__15093),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__2753 (
            .O(N__15090),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__2752 (
            .O(N__15087),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__2751 (
            .O(N__15084),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__2750 (
            .O(N__15081),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__2749 (
            .O(N__15078),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__2748 (
            .O(N__15069),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__2747 (
            .O(N__15066),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__2746 (
            .O(N__15063),
            .I(\transmit_module.VGA_VISIBLE ));
    InMux I__2745 (
            .O(N__15044),
            .I(N__15041));
    LocalMux I__2744 (
            .O(N__15041),
            .I(\transmit_module.n130 ));
    InMux I__2743 (
            .O(N__15038),
            .I(\receive_module.n3161 ));
    SRMux I__2742 (
            .O(N__15035),
            .I(N__15032));
    LocalMux I__2741 (
            .O(N__15032),
            .I(N__15028));
    SRMux I__2740 (
            .O(N__15031),
            .I(N__15025));
    Span4Mux_v I__2739 (
            .O(N__15028),
            .I(N__15019));
    LocalMux I__2738 (
            .O(N__15025),
            .I(N__15019));
    SRMux I__2737 (
            .O(N__15024),
            .I(N__15016));
    Span4Mux_v I__2736 (
            .O(N__15019),
            .I(N__15010));
    LocalMux I__2735 (
            .O(N__15016),
            .I(N__15010));
    SRMux I__2734 (
            .O(N__15015),
            .I(N__15007));
    Span4Mux_v I__2733 (
            .O(N__15010),
            .I(N__15002));
    LocalMux I__2732 (
            .O(N__15007),
            .I(N__15002));
    Span4Mux_h I__2731 (
            .O(N__15002),
            .I(N__14999));
    Span4Mux_h I__2730 (
            .O(N__14999),
            .I(N__14996));
    Odrv4 I__2729 (
            .O(N__14996),
            .I(\line_buffer.n606 ));
    SRMux I__2728 (
            .O(N__14993),
            .I(N__14989));
    SRMux I__2727 (
            .O(N__14992),
            .I(N__14984));
    LocalMux I__2726 (
            .O(N__14989),
            .I(N__14981));
    SRMux I__2725 (
            .O(N__14988),
            .I(N__14978));
    SRMux I__2724 (
            .O(N__14987),
            .I(N__14975));
    LocalMux I__2723 (
            .O(N__14984),
            .I(N__14972));
    Span4Mux_s2_v I__2722 (
            .O(N__14981),
            .I(N__14965));
    LocalMux I__2721 (
            .O(N__14978),
            .I(N__14965));
    LocalMux I__2720 (
            .O(N__14975),
            .I(N__14965));
    Span4Mux_h I__2719 (
            .O(N__14972),
            .I(N__14962));
    Span4Mux_v I__2718 (
            .O(N__14965),
            .I(N__14959));
    Span4Mux_v I__2717 (
            .O(N__14962),
            .I(N__14956));
    Sp12to4 I__2716 (
            .O(N__14959),
            .I(N__14953));
    Span4Mux_h I__2715 (
            .O(N__14956),
            .I(N__14950));
    Span12Mux_v I__2714 (
            .O(N__14953),
            .I(N__14947));
    Span4Mux_h I__2713 (
            .O(N__14950),
            .I(N__14944));
    Odrv12 I__2712 (
            .O(N__14947),
            .I(\line_buffer.n476 ));
    Odrv4 I__2711 (
            .O(N__14944),
            .I(\line_buffer.n476 ));
    CEMux I__2710 (
            .O(N__14939),
            .I(N__14936));
    LocalMux I__2709 (
            .O(N__14936),
            .I(N__14933));
    Span4Mux_h I__2708 (
            .O(N__14933),
            .I(N__14930));
    Odrv4 I__2707 (
            .O(N__14930),
            .I(\receive_module.n3674 ));
    InMux I__2706 (
            .O(N__14927),
            .I(N__14924));
    LocalMux I__2705 (
            .O(N__14924),
            .I(N__14913));
    InMux I__2704 (
            .O(N__14923),
            .I(N__14910));
    InMux I__2703 (
            .O(N__14922),
            .I(N__14903));
    InMux I__2702 (
            .O(N__14921),
            .I(N__14903));
    InMux I__2701 (
            .O(N__14920),
            .I(N__14903));
    InMux I__2700 (
            .O(N__14919),
            .I(N__14896));
    InMux I__2699 (
            .O(N__14918),
            .I(N__14896));
    InMux I__2698 (
            .O(N__14917),
            .I(N__14896));
    InMux I__2697 (
            .O(N__14916),
            .I(N__14893));
    Odrv4 I__2696 (
            .O(N__14913),
            .I(RX_ADDR_11));
    LocalMux I__2695 (
            .O(N__14910),
            .I(RX_ADDR_11));
    LocalMux I__2694 (
            .O(N__14903),
            .I(RX_ADDR_11));
    LocalMux I__2693 (
            .O(N__14896),
            .I(RX_ADDR_11));
    LocalMux I__2692 (
            .O(N__14893),
            .I(RX_ADDR_11));
    CascadeMux I__2691 (
            .O(N__14882),
            .I(N__14876));
    InMux I__2690 (
            .O(N__14881),
            .I(N__14869));
    InMux I__2689 (
            .O(N__14880),
            .I(N__14869));
    InMux I__2688 (
            .O(N__14879),
            .I(N__14869));
    InMux I__2687 (
            .O(N__14876),
            .I(N__14861));
    LocalMux I__2686 (
            .O(N__14869),
            .I(N__14858));
    InMux I__2685 (
            .O(N__14868),
            .I(N__14855));
    InMux I__2684 (
            .O(N__14867),
            .I(N__14852));
    InMux I__2683 (
            .O(N__14866),
            .I(N__14847));
    InMux I__2682 (
            .O(N__14865),
            .I(N__14847));
    InMux I__2681 (
            .O(N__14864),
            .I(N__14844));
    LocalMux I__2680 (
            .O(N__14861),
            .I(N__14839));
    Span4Mux_v I__2679 (
            .O(N__14858),
            .I(N__14839));
    LocalMux I__2678 (
            .O(N__14855),
            .I(RX_ADDR_12));
    LocalMux I__2677 (
            .O(N__14852),
            .I(RX_ADDR_12));
    LocalMux I__2676 (
            .O(N__14847),
            .I(RX_ADDR_12));
    LocalMux I__2675 (
            .O(N__14844),
            .I(RX_ADDR_12));
    Odrv4 I__2674 (
            .O(N__14839),
            .I(RX_ADDR_12));
    InMux I__2673 (
            .O(N__14828),
            .I(N__14818));
    CascadeMux I__2672 (
            .O(N__14827),
            .I(N__14814));
    CascadeMux I__2671 (
            .O(N__14826),
            .I(N__14811));
    CascadeMux I__2670 (
            .O(N__14825),
            .I(N__14808));
    CascadeMux I__2669 (
            .O(N__14824),
            .I(N__14805));
    CascadeMux I__2668 (
            .O(N__14823),
            .I(N__14802));
    CascadeMux I__2667 (
            .O(N__14822),
            .I(N__14799));
    CascadeMux I__2666 (
            .O(N__14821),
            .I(N__14796));
    LocalMux I__2665 (
            .O(N__14818),
            .I(N__14793));
    InMux I__2664 (
            .O(N__14817),
            .I(N__14790));
    InMux I__2663 (
            .O(N__14814),
            .I(N__14787));
    InMux I__2662 (
            .O(N__14811),
            .I(N__14784));
    InMux I__2661 (
            .O(N__14808),
            .I(N__14781));
    InMux I__2660 (
            .O(N__14805),
            .I(N__14776));
    InMux I__2659 (
            .O(N__14802),
            .I(N__14776));
    InMux I__2658 (
            .O(N__14799),
            .I(N__14771));
    InMux I__2657 (
            .O(N__14796),
            .I(N__14771));
    Span4Mux_v I__2656 (
            .O(N__14793),
            .I(N__14768));
    LocalMux I__2655 (
            .O(N__14790),
            .I(RX_ADDR_13));
    LocalMux I__2654 (
            .O(N__14787),
            .I(RX_ADDR_13));
    LocalMux I__2653 (
            .O(N__14784),
            .I(RX_ADDR_13));
    LocalMux I__2652 (
            .O(N__14781),
            .I(RX_ADDR_13));
    LocalMux I__2651 (
            .O(N__14776),
            .I(RX_ADDR_13));
    LocalMux I__2650 (
            .O(N__14771),
            .I(RX_ADDR_13));
    Odrv4 I__2649 (
            .O(N__14768),
            .I(RX_ADDR_13));
    SRMux I__2648 (
            .O(N__14753),
            .I(N__14750));
    LocalMux I__2647 (
            .O(N__14750),
            .I(N__14745));
    SRMux I__2646 (
            .O(N__14749),
            .I(N__14742));
    SRMux I__2645 (
            .O(N__14748),
            .I(N__14738));
    Span4Mux_h I__2644 (
            .O(N__14745),
            .I(N__14735));
    LocalMux I__2643 (
            .O(N__14742),
            .I(N__14732));
    SRMux I__2642 (
            .O(N__14741),
            .I(N__14729));
    LocalMux I__2641 (
            .O(N__14738),
            .I(N__14726));
    Span4Mux_h I__2640 (
            .O(N__14735),
            .I(N__14723));
    Span4Mux_h I__2639 (
            .O(N__14732),
            .I(N__14720));
    LocalMux I__2638 (
            .O(N__14729),
            .I(N__14717));
    Span4Mux_h I__2637 (
            .O(N__14726),
            .I(N__14714));
    Span4Mux_v I__2636 (
            .O(N__14723),
            .I(N__14711));
    Span4Mux_v I__2635 (
            .O(N__14720),
            .I(N__14706));
    Span4Mux_h I__2634 (
            .O(N__14717),
            .I(N__14706));
    Span4Mux_h I__2633 (
            .O(N__14714),
            .I(N__14703));
    Span4Mux_v I__2632 (
            .O(N__14711),
            .I(N__14698));
    Span4Mux_h I__2631 (
            .O(N__14706),
            .I(N__14698));
    Odrv4 I__2630 (
            .O(N__14703),
            .I(\line_buffer.n574 ));
    Odrv4 I__2629 (
            .O(N__14698),
            .I(\line_buffer.n574 ));
    InMux I__2628 (
            .O(N__14693),
            .I(N__14690));
    LocalMux I__2627 (
            .O(N__14690),
            .I(N__14687));
    Span4Mux_v I__2626 (
            .O(N__14687),
            .I(N__14684));
    Odrv4 I__2625 (
            .O(N__14684),
            .I(\tvp_vs_buffer.BUFFER_1_0 ));
    InMux I__2624 (
            .O(N__14681),
            .I(N__14678));
    LocalMux I__2623 (
            .O(N__14678),
            .I(\tvp_vs_buffer.BUFFER_2_0 ));
    InMux I__2622 (
            .O(N__14675),
            .I(N__14672));
    LocalMux I__2621 (
            .O(N__14672),
            .I(N__14668));
    CascadeMux I__2620 (
            .O(N__14671),
            .I(N__14665));
    Span4Mux_h I__2619 (
            .O(N__14668),
            .I(N__14662));
    InMux I__2618 (
            .O(N__14665),
            .I(N__14659));
    Odrv4 I__2617 (
            .O(N__14662),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    LocalMux I__2616 (
            .O(N__14659),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    InMux I__2615 (
            .O(N__14654),
            .I(\receive_module.n3152 ));
    InMux I__2614 (
            .O(N__14651),
            .I(\receive_module.n3153 ));
    InMux I__2613 (
            .O(N__14648),
            .I(\receive_module.n3154 ));
    InMux I__2612 (
            .O(N__14645),
            .I(\receive_module.n3155 ));
    InMux I__2611 (
            .O(N__14642),
            .I(bfn_15_12_0_));
    InMux I__2610 (
            .O(N__14639),
            .I(\receive_module.n3157 ));
    InMux I__2609 (
            .O(N__14636),
            .I(\receive_module.n3158 ));
    InMux I__2608 (
            .O(N__14633),
            .I(\receive_module.n3159 ));
    InMux I__2607 (
            .O(N__14630),
            .I(\receive_module.n3160 ));
    InMux I__2606 (
            .O(N__14627),
            .I(N__14624));
    LocalMux I__2605 (
            .O(N__14624),
            .I(\transmit_module.X_DELTA_PATTERN_10 ));
    InMux I__2604 (
            .O(N__14621),
            .I(N__14618));
    LocalMux I__2603 (
            .O(N__14618),
            .I(\transmit_module.X_DELTA_PATTERN_9 ));
    InMux I__2602 (
            .O(N__14615),
            .I(N__14612));
    LocalMux I__2601 (
            .O(N__14612),
            .I(\transmit_module.X_DELTA_PATTERN_11 ));
    InMux I__2600 (
            .O(N__14609),
            .I(N__14606));
    LocalMux I__2599 (
            .O(N__14606),
            .I(N__14603));
    Span4Mux_h I__2598 (
            .O(N__14603),
            .I(N__14600));
    Odrv4 I__2597 (
            .O(N__14600),
            .I(\transmit_module.X_DELTA_PATTERN_13 ));
    InMux I__2596 (
            .O(N__14597),
            .I(N__14594));
    LocalMux I__2595 (
            .O(N__14594),
            .I(\transmit_module.X_DELTA_PATTERN_12 ));
    InMux I__2594 (
            .O(N__14591),
            .I(bfn_15_11_0_));
    InMux I__2593 (
            .O(N__14588),
            .I(\receive_module.n3149 ));
    InMux I__2592 (
            .O(N__14585),
            .I(\receive_module.n3150 ));
    InMux I__2591 (
            .O(N__14582),
            .I(\receive_module.n3151 ));
    InMux I__2590 (
            .O(N__14579),
            .I(N__14575));
    CascadeMux I__2589 (
            .O(N__14578),
            .I(N__14570));
    LocalMux I__2588 (
            .O(N__14575),
            .I(N__14567));
    InMux I__2587 (
            .O(N__14574),
            .I(N__14564));
    InMux I__2586 (
            .O(N__14573),
            .I(N__14561));
    InMux I__2585 (
            .O(N__14570),
            .I(N__14558));
    Odrv4 I__2584 (
            .O(N__14567),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__2583 (
            .O(N__14564),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__2582 (
            .O(N__14561),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__2581 (
            .O(N__14558),
            .I(\transmit_module.TX_ADDR_10 ));
    InMux I__2580 (
            .O(N__14549),
            .I(N__14546));
    LocalMux I__2579 (
            .O(N__14546),
            .I(N__14543));
    Odrv4 I__2578 (
            .O(N__14543),
            .I(\transmit_module.ADDR_Y_COMPONENT_10 ));
    InMux I__2577 (
            .O(N__14540),
            .I(N__14536));
    CascadeMux I__2576 (
            .O(N__14539),
            .I(N__14531));
    LocalMux I__2575 (
            .O(N__14536),
            .I(N__14528));
    InMux I__2574 (
            .O(N__14535),
            .I(N__14523));
    InMux I__2573 (
            .O(N__14534),
            .I(N__14523));
    InMux I__2572 (
            .O(N__14531),
            .I(N__14520));
    Odrv4 I__2571 (
            .O(N__14528),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__2570 (
            .O(N__14523),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__2569 (
            .O(N__14520),
            .I(\transmit_module.TX_ADDR_8 ));
    InMux I__2568 (
            .O(N__14513),
            .I(N__14510));
    LocalMux I__2567 (
            .O(N__14510),
            .I(N__14507));
    Odrv4 I__2566 (
            .O(N__14507),
            .I(\transmit_module.ADDR_Y_COMPONENT_8 ));
    InMux I__2565 (
            .O(N__14504),
            .I(N__14499));
    InMux I__2564 (
            .O(N__14503),
            .I(N__14496));
    InMux I__2563 (
            .O(N__14502),
            .I(N__14493));
    LocalMux I__2562 (
            .O(N__14499),
            .I(N__14489));
    LocalMux I__2561 (
            .O(N__14496),
            .I(N__14486));
    LocalMux I__2560 (
            .O(N__14493),
            .I(N__14483));
    InMux I__2559 (
            .O(N__14492),
            .I(N__14480));
    Odrv12 I__2558 (
            .O(N__14489),
            .I(\transmit_module.TX_ADDR_1 ));
    Odrv4 I__2557 (
            .O(N__14486),
            .I(\transmit_module.TX_ADDR_1 ));
    Odrv4 I__2556 (
            .O(N__14483),
            .I(\transmit_module.TX_ADDR_1 ));
    LocalMux I__2555 (
            .O(N__14480),
            .I(\transmit_module.TX_ADDR_1 ));
    InMux I__2554 (
            .O(N__14471),
            .I(N__14468));
    LocalMux I__2553 (
            .O(N__14468),
            .I(\transmit_module.ADDR_Y_COMPONENT_1 ));
    InMux I__2552 (
            .O(N__14465),
            .I(N__14462));
    LocalMux I__2551 (
            .O(N__14462),
            .I(N__14457));
    InMux I__2550 (
            .O(N__14461),
            .I(N__14454));
    InMux I__2549 (
            .O(N__14460),
            .I(N__14451));
    Span12Mux_v I__2548 (
            .O(N__14457),
            .I(N__14443));
    LocalMux I__2547 (
            .O(N__14454),
            .I(N__14443));
    LocalMux I__2546 (
            .O(N__14451),
            .I(N__14443));
    InMux I__2545 (
            .O(N__14450),
            .I(N__14440));
    Odrv12 I__2544 (
            .O(N__14443),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__2543 (
            .O(N__14440),
            .I(\transmit_module.TX_ADDR_0 ));
    InMux I__2542 (
            .O(N__14435),
            .I(N__14432));
    LocalMux I__2541 (
            .O(N__14432),
            .I(N__14429));
    Odrv4 I__2540 (
            .O(N__14429),
            .I(\transmit_module.ADDR_Y_COMPONENT_0 ));
    IoInMux I__2539 (
            .O(N__14426),
            .I(N__14423));
    LocalMux I__2538 (
            .O(N__14423),
            .I(N__14420));
    IoSpan4Mux I__2537 (
            .O(N__14420),
            .I(N__14417));
    Span4Mux_s1_h I__2536 (
            .O(N__14417),
            .I(N__14414));
    Sp12to4 I__2535 (
            .O(N__14414),
            .I(N__14410));
    InMux I__2534 (
            .O(N__14413),
            .I(N__14407));
    Span12Mux_h I__2533 (
            .O(N__14410),
            .I(N__14402));
    LocalMux I__2532 (
            .O(N__14407),
            .I(N__14402));
    Odrv12 I__2531 (
            .O(N__14402),
            .I(DEBUG_c_1_c));
    IoInMux I__2530 (
            .O(N__14399),
            .I(N__14396));
    LocalMux I__2529 (
            .O(N__14396),
            .I(N__14393));
    IoSpan4Mux I__2528 (
            .O(N__14393),
            .I(N__14390));
    Span4Mux_s0_h I__2527 (
            .O(N__14390),
            .I(N__14386));
    InMux I__2526 (
            .O(N__14389),
            .I(N__14383));
    Sp12to4 I__2525 (
            .O(N__14386),
            .I(N__14380));
    LocalMux I__2524 (
            .O(N__14383),
            .I(N__14377));
    Span12Mux_s11_h I__2523 (
            .O(N__14380),
            .I(N__14374));
    Span4Mux_h I__2522 (
            .O(N__14377),
            .I(N__14371));
    Span12Mux_v I__2521 (
            .O(N__14374),
            .I(N__14368));
    Span4Mux_v I__2520 (
            .O(N__14371),
            .I(N__14365));
    Odrv12 I__2519 (
            .O(N__14368),
            .I(DEBUG_c_6_c));
    Odrv4 I__2518 (
            .O(N__14365),
            .I(DEBUG_c_6_c));
    InMux I__2517 (
            .O(N__14360),
            .I(N__14357));
    LocalMux I__2516 (
            .O(N__14357),
            .I(N__14354));
    Odrv4 I__2515 (
            .O(N__14354),
            .I(\tvp_vs_buffer.BUFFER_0_0 ));
    InMux I__2514 (
            .O(N__14351),
            .I(N__14348));
    LocalMux I__2513 (
            .O(N__14348),
            .I(\tvp_video_buffer.BUFFER_0_6 ));
    CascadeMux I__2512 (
            .O(N__14345),
            .I(N__14341));
    InMux I__2511 (
            .O(N__14344),
            .I(N__14336));
    InMux I__2510 (
            .O(N__14341),
            .I(N__14336));
    LocalMux I__2509 (
            .O(N__14336),
            .I(N__14332));
    InMux I__2508 (
            .O(N__14335),
            .I(N__14329));
    Odrv4 I__2507 (
            .O(N__14332),
            .I(TVP_HSYNC_buff));
    LocalMux I__2506 (
            .O(N__14329),
            .I(TVP_HSYNC_buff));
    InMux I__2505 (
            .O(N__14324),
            .I(N__14321));
    LocalMux I__2504 (
            .O(N__14321),
            .I(N__14318));
    Span4Mux_h I__2503 (
            .O(N__14318),
            .I(N__14315));
    Odrv4 I__2502 (
            .O(N__14315),
            .I(\transmit_module.n138 ));
    InMux I__2501 (
            .O(N__14312),
            .I(N__14309));
    LocalMux I__2500 (
            .O(N__14309),
            .I(N__14306));
    Span4Mux_h I__2499 (
            .O(N__14306),
            .I(N__14302));
    InMux I__2498 (
            .O(N__14305),
            .I(N__14299));
    Odrv4 I__2497 (
            .O(N__14302),
            .I(\transmit_module.video_signal_controller.n3382 ));
    LocalMux I__2496 (
            .O(N__14299),
            .I(\transmit_module.video_signal_controller.n3382 ));
    InMux I__2495 (
            .O(N__14294),
            .I(N__14291));
    LocalMux I__2494 (
            .O(N__14291),
            .I(\transmit_module.video_signal_controller.n3017 ));
    CascadeMux I__2493 (
            .O(N__14288),
            .I(N__14284));
    CascadeMux I__2492 (
            .O(N__14287),
            .I(N__14281));
    InMux I__2491 (
            .O(N__14284),
            .I(N__14278));
    InMux I__2490 (
            .O(N__14281),
            .I(N__14274));
    LocalMux I__2489 (
            .O(N__14278),
            .I(N__14270));
    InMux I__2488 (
            .O(N__14277),
            .I(N__14266));
    LocalMux I__2487 (
            .O(N__14274),
            .I(N__14263));
    InMux I__2486 (
            .O(N__14273),
            .I(N__14260));
    Span4Mux_h I__2485 (
            .O(N__14270),
            .I(N__14257));
    InMux I__2484 (
            .O(N__14269),
            .I(N__14254));
    LocalMux I__2483 (
            .O(N__14266),
            .I(N__14247));
    Span4Mux_v I__2482 (
            .O(N__14263),
            .I(N__14247));
    LocalMux I__2481 (
            .O(N__14260),
            .I(N__14247));
    Odrv4 I__2480 (
            .O(N__14257),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    LocalMux I__2479 (
            .O(N__14254),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    Odrv4 I__2478 (
            .O(N__14247),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    InMux I__2477 (
            .O(N__14240),
            .I(N__14237));
    LocalMux I__2476 (
            .O(N__14237),
            .I(\transmit_module.video_signal_controller.n7_adj_624 ));
    InMux I__2475 (
            .O(N__14234),
            .I(N__14231));
    LocalMux I__2474 (
            .O(N__14231),
            .I(N__14228));
    Odrv12 I__2473 (
            .O(N__14228),
            .I(\transmit_module.n132 ));
    InMux I__2472 (
            .O(N__14225),
            .I(N__14222));
    LocalMux I__2471 (
            .O(N__14222),
            .I(N__14219));
    Odrv12 I__2470 (
            .O(N__14219),
            .I(\transmit_module.ADDR_Y_COMPONENT_9 ));
    InMux I__2469 (
            .O(N__14216),
            .I(N__14213));
    LocalMux I__2468 (
            .O(N__14213),
            .I(N__14207));
    InMux I__2467 (
            .O(N__14212),
            .I(N__14204));
    InMux I__2466 (
            .O(N__14211),
            .I(N__14201));
    CascadeMux I__2465 (
            .O(N__14210),
            .I(N__14198));
    Span4Mux_h I__2464 (
            .O(N__14207),
            .I(N__14195));
    LocalMux I__2463 (
            .O(N__14204),
            .I(N__14190));
    LocalMux I__2462 (
            .O(N__14201),
            .I(N__14190));
    InMux I__2461 (
            .O(N__14198),
            .I(N__14187));
    Odrv4 I__2460 (
            .O(N__14195),
            .I(\transmit_module.TX_ADDR_9 ));
    Odrv4 I__2459 (
            .O(N__14190),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__2458 (
            .O(N__14187),
            .I(\transmit_module.TX_ADDR_9 ));
    InMux I__2457 (
            .O(N__14180),
            .I(N__14177));
    LocalMux I__2456 (
            .O(N__14177),
            .I(N__14173));
    InMux I__2455 (
            .O(N__14176),
            .I(N__14170));
    Odrv4 I__2454 (
            .O(N__14173),
            .I(\transmit_module.n107 ));
    LocalMux I__2453 (
            .O(N__14170),
            .I(\transmit_module.n107 ));
    InMux I__2452 (
            .O(N__14165),
            .I(N__14161));
    InMux I__2451 (
            .O(N__14164),
            .I(N__14158));
    LocalMux I__2450 (
            .O(N__14161),
            .I(N__14155));
    LocalMux I__2449 (
            .O(N__14158),
            .I(N__14152));
    Span4Mux_h I__2448 (
            .O(N__14155),
            .I(N__14149));
    Odrv4 I__2447 (
            .O(N__14152),
            .I(\transmit_module.n115 ));
    Odrv4 I__2446 (
            .O(N__14149),
            .I(\transmit_module.n115 ));
    InMux I__2445 (
            .O(N__14144),
            .I(N__14141));
    LocalMux I__2444 (
            .O(N__14141),
            .I(N__14138));
    Span4Mux_v I__2443 (
            .O(N__14138),
            .I(N__14135));
    Odrv4 I__2442 (
            .O(N__14135),
            .I(\transmit_module.n116 ));
    CascadeMux I__2441 (
            .O(N__14132),
            .I(\transmit_module.n116_cascade_ ));
    InMux I__2440 (
            .O(N__14129),
            .I(N__14126));
    LocalMux I__2439 (
            .O(N__14126),
            .I(N__14122));
    InMux I__2438 (
            .O(N__14125),
            .I(N__14119));
    Odrv12 I__2437 (
            .O(N__14122),
            .I(\transmit_module.n147 ));
    LocalMux I__2436 (
            .O(N__14119),
            .I(\transmit_module.n147 ));
    CascadeMux I__2435 (
            .O(N__14114),
            .I(N__14110));
    CascadeMux I__2434 (
            .O(N__14113),
            .I(N__14107));
    CascadeBuf I__2433 (
            .O(N__14110),
            .I(N__14104));
    CascadeBuf I__2432 (
            .O(N__14107),
            .I(N__14101));
    CascadeMux I__2431 (
            .O(N__14104),
            .I(N__14098));
    CascadeMux I__2430 (
            .O(N__14101),
            .I(N__14095));
    CascadeBuf I__2429 (
            .O(N__14098),
            .I(N__14092));
    CascadeBuf I__2428 (
            .O(N__14095),
            .I(N__14089));
    CascadeMux I__2427 (
            .O(N__14092),
            .I(N__14086));
    CascadeMux I__2426 (
            .O(N__14089),
            .I(N__14083));
    CascadeBuf I__2425 (
            .O(N__14086),
            .I(N__14080));
    CascadeBuf I__2424 (
            .O(N__14083),
            .I(N__14077));
    CascadeMux I__2423 (
            .O(N__14080),
            .I(N__14074));
    CascadeMux I__2422 (
            .O(N__14077),
            .I(N__14071));
    CascadeBuf I__2421 (
            .O(N__14074),
            .I(N__14068));
    CascadeBuf I__2420 (
            .O(N__14071),
            .I(N__14065));
    CascadeMux I__2419 (
            .O(N__14068),
            .I(N__14062));
    CascadeMux I__2418 (
            .O(N__14065),
            .I(N__14059));
    CascadeBuf I__2417 (
            .O(N__14062),
            .I(N__14056));
    CascadeBuf I__2416 (
            .O(N__14059),
            .I(N__14053));
    CascadeMux I__2415 (
            .O(N__14056),
            .I(N__14050));
    CascadeMux I__2414 (
            .O(N__14053),
            .I(N__14047));
    CascadeBuf I__2413 (
            .O(N__14050),
            .I(N__14044));
    CascadeBuf I__2412 (
            .O(N__14047),
            .I(N__14041));
    CascadeMux I__2411 (
            .O(N__14044),
            .I(N__14038));
    CascadeMux I__2410 (
            .O(N__14041),
            .I(N__14035));
    CascadeBuf I__2409 (
            .O(N__14038),
            .I(N__14032));
    CascadeBuf I__2408 (
            .O(N__14035),
            .I(N__14029));
    CascadeMux I__2407 (
            .O(N__14032),
            .I(N__14026));
    CascadeMux I__2406 (
            .O(N__14029),
            .I(N__14023));
    CascadeBuf I__2405 (
            .O(N__14026),
            .I(N__14020));
    CascadeBuf I__2404 (
            .O(N__14023),
            .I(N__14017));
    CascadeMux I__2403 (
            .O(N__14020),
            .I(N__14014));
    CascadeMux I__2402 (
            .O(N__14017),
            .I(N__14011));
    CascadeBuf I__2401 (
            .O(N__14014),
            .I(N__14008));
    CascadeBuf I__2400 (
            .O(N__14011),
            .I(N__14005));
    CascadeMux I__2399 (
            .O(N__14008),
            .I(N__14002));
    CascadeMux I__2398 (
            .O(N__14005),
            .I(N__13999));
    CascadeBuf I__2397 (
            .O(N__14002),
            .I(N__13996));
    CascadeBuf I__2396 (
            .O(N__13999),
            .I(N__13993));
    CascadeMux I__2395 (
            .O(N__13996),
            .I(N__13990));
    CascadeMux I__2394 (
            .O(N__13993),
            .I(N__13987));
    CascadeBuf I__2393 (
            .O(N__13990),
            .I(N__13984));
    CascadeBuf I__2392 (
            .O(N__13987),
            .I(N__13981));
    CascadeMux I__2391 (
            .O(N__13984),
            .I(N__13978));
    CascadeMux I__2390 (
            .O(N__13981),
            .I(N__13975));
    CascadeBuf I__2389 (
            .O(N__13978),
            .I(N__13972));
    CascadeBuf I__2388 (
            .O(N__13975),
            .I(N__13969));
    CascadeMux I__2387 (
            .O(N__13972),
            .I(N__13966));
    CascadeMux I__2386 (
            .O(N__13969),
            .I(N__13963));
    CascadeBuf I__2385 (
            .O(N__13966),
            .I(N__13960));
    CascadeBuf I__2384 (
            .O(N__13963),
            .I(N__13957));
    CascadeMux I__2383 (
            .O(N__13960),
            .I(N__13954));
    CascadeMux I__2382 (
            .O(N__13957),
            .I(N__13951));
    CascadeBuf I__2381 (
            .O(N__13954),
            .I(N__13948));
    CascadeBuf I__2380 (
            .O(N__13951),
            .I(N__13945));
    CascadeMux I__2379 (
            .O(N__13948),
            .I(N__13942));
    CascadeMux I__2378 (
            .O(N__13945),
            .I(N__13939));
    CascadeBuf I__2377 (
            .O(N__13942),
            .I(N__13936));
    CascadeBuf I__2376 (
            .O(N__13939),
            .I(N__13933));
    CascadeMux I__2375 (
            .O(N__13936),
            .I(N__13930));
    CascadeMux I__2374 (
            .O(N__13933),
            .I(N__13927));
    InMux I__2373 (
            .O(N__13930),
            .I(N__13924));
    InMux I__2372 (
            .O(N__13927),
            .I(N__13921));
    LocalMux I__2371 (
            .O(N__13924),
            .I(N__13918));
    LocalMux I__2370 (
            .O(N__13921),
            .I(N__13915));
    Span4Mux_h I__2369 (
            .O(N__13918),
            .I(N__13912));
    Span12Mux_h I__2368 (
            .O(N__13915),
            .I(N__13909));
    Sp12to4 I__2367 (
            .O(N__13912),
            .I(N__13906));
    Span12Mux_v I__2366 (
            .O(N__13909),
            .I(N__13903));
    Span12Mux_v I__2365 (
            .O(N__13906),
            .I(N__13900));
    Odrv12 I__2364 (
            .O(N__13903),
            .I(n28));
    Odrv12 I__2363 (
            .O(N__13900),
            .I(n28));
    InMux I__2362 (
            .O(N__13895),
            .I(N__13891));
    InMux I__2361 (
            .O(N__13894),
            .I(N__13888));
    LocalMux I__2360 (
            .O(N__13891),
            .I(\transmit_module.n106 ));
    LocalMux I__2359 (
            .O(N__13888),
            .I(\transmit_module.n106 ));
    InMux I__2358 (
            .O(N__13883),
            .I(N__13880));
    LocalMux I__2357 (
            .O(N__13880),
            .I(N__13877));
    Odrv4 I__2356 (
            .O(N__13877),
            .I(\transmit_module.n137 ));
    CascadeMux I__2355 (
            .O(N__13874),
            .I(N__13871));
    CascadeBuf I__2354 (
            .O(N__13871),
            .I(N__13867));
    CascadeMux I__2353 (
            .O(N__13870),
            .I(N__13864));
    CascadeMux I__2352 (
            .O(N__13867),
            .I(N__13861));
    CascadeBuf I__2351 (
            .O(N__13864),
            .I(N__13858));
    CascadeBuf I__2350 (
            .O(N__13861),
            .I(N__13855));
    CascadeMux I__2349 (
            .O(N__13858),
            .I(N__13852));
    CascadeMux I__2348 (
            .O(N__13855),
            .I(N__13849));
    CascadeBuf I__2347 (
            .O(N__13852),
            .I(N__13846));
    CascadeBuf I__2346 (
            .O(N__13849),
            .I(N__13843));
    CascadeMux I__2345 (
            .O(N__13846),
            .I(N__13840));
    CascadeMux I__2344 (
            .O(N__13843),
            .I(N__13837));
    CascadeBuf I__2343 (
            .O(N__13840),
            .I(N__13834));
    CascadeBuf I__2342 (
            .O(N__13837),
            .I(N__13831));
    CascadeMux I__2341 (
            .O(N__13834),
            .I(N__13828));
    CascadeMux I__2340 (
            .O(N__13831),
            .I(N__13825));
    CascadeBuf I__2339 (
            .O(N__13828),
            .I(N__13822));
    CascadeBuf I__2338 (
            .O(N__13825),
            .I(N__13819));
    CascadeMux I__2337 (
            .O(N__13822),
            .I(N__13816));
    CascadeMux I__2336 (
            .O(N__13819),
            .I(N__13813));
    CascadeBuf I__2335 (
            .O(N__13816),
            .I(N__13810));
    CascadeBuf I__2334 (
            .O(N__13813),
            .I(N__13807));
    CascadeMux I__2333 (
            .O(N__13810),
            .I(N__13804));
    CascadeMux I__2332 (
            .O(N__13807),
            .I(N__13801));
    CascadeBuf I__2331 (
            .O(N__13804),
            .I(N__13798));
    CascadeBuf I__2330 (
            .O(N__13801),
            .I(N__13795));
    CascadeMux I__2329 (
            .O(N__13798),
            .I(N__13792));
    CascadeMux I__2328 (
            .O(N__13795),
            .I(N__13789));
    CascadeBuf I__2327 (
            .O(N__13792),
            .I(N__13786));
    CascadeBuf I__2326 (
            .O(N__13789),
            .I(N__13783));
    CascadeMux I__2325 (
            .O(N__13786),
            .I(N__13780));
    CascadeMux I__2324 (
            .O(N__13783),
            .I(N__13777));
    CascadeBuf I__2323 (
            .O(N__13780),
            .I(N__13774));
    CascadeBuf I__2322 (
            .O(N__13777),
            .I(N__13771));
    CascadeMux I__2321 (
            .O(N__13774),
            .I(N__13768));
    CascadeMux I__2320 (
            .O(N__13771),
            .I(N__13765));
    CascadeBuf I__2319 (
            .O(N__13768),
            .I(N__13762));
    CascadeBuf I__2318 (
            .O(N__13765),
            .I(N__13759));
    CascadeMux I__2317 (
            .O(N__13762),
            .I(N__13756));
    CascadeMux I__2316 (
            .O(N__13759),
            .I(N__13753));
    CascadeBuf I__2315 (
            .O(N__13756),
            .I(N__13750));
    CascadeBuf I__2314 (
            .O(N__13753),
            .I(N__13747));
    CascadeMux I__2313 (
            .O(N__13750),
            .I(N__13744));
    CascadeMux I__2312 (
            .O(N__13747),
            .I(N__13741));
    CascadeBuf I__2311 (
            .O(N__13744),
            .I(N__13738));
    CascadeBuf I__2310 (
            .O(N__13741),
            .I(N__13735));
    CascadeMux I__2309 (
            .O(N__13738),
            .I(N__13732));
    CascadeMux I__2308 (
            .O(N__13735),
            .I(N__13729));
    CascadeBuf I__2307 (
            .O(N__13732),
            .I(N__13726));
    CascadeBuf I__2306 (
            .O(N__13729),
            .I(N__13723));
    CascadeMux I__2305 (
            .O(N__13726),
            .I(N__13720));
    CascadeMux I__2304 (
            .O(N__13723),
            .I(N__13717));
    CascadeBuf I__2303 (
            .O(N__13720),
            .I(N__13714));
    CascadeBuf I__2302 (
            .O(N__13717),
            .I(N__13711));
    CascadeMux I__2301 (
            .O(N__13714),
            .I(N__13708));
    CascadeMux I__2300 (
            .O(N__13711),
            .I(N__13705));
    CascadeBuf I__2299 (
            .O(N__13708),
            .I(N__13702));
    CascadeBuf I__2298 (
            .O(N__13705),
            .I(N__13699));
    CascadeMux I__2297 (
            .O(N__13702),
            .I(N__13696));
    CascadeMux I__2296 (
            .O(N__13699),
            .I(N__13693));
    CascadeBuf I__2295 (
            .O(N__13696),
            .I(N__13690));
    InMux I__2294 (
            .O(N__13693),
            .I(N__13687));
    CascadeMux I__2293 (
            .O(N__13690),
            .I(N__13684));
    LocalMux I__2292 (
            .O(N__13687),
            .I(N__13681));
    InMux I__2291 (
            .O(N__13684),
            .I(N__13678));
    Span4Mux_h I__2290 (
            .O(N__13681),
            .I(N__13675));
    LocalMux I__2289 (
            .O(N__13678),
            .I(N__13672));
    Sp12to4 I__2288 (
            .O(N__13675),
            .I(N__13669));
    Sp12to4 I__2287 (
            .O(N__13672),
            .I(N__13666));
    Span12Mux_h I__2286 (
            .O(N__13669),
            .I(N__13661));
    Span12Mux_s9_h I__2285 (
            .O(N__13666),
            .I(N__13661));
    Span12Mux_v I__2284 (
            .O(N__13661),
            .I(N__13658));
    Odrv12 I__2283 (
            .O(N__13658),
            .I(n18));
    InMux I__2282 (
            .O(N__13655),
            .I(N__13652));
    LocalMux I__2281 (
            .O(N__13652),
            .I(N__13649));
    Odrv4 I__2280 (
            .O(N__13649),
            .I(\transmit_module.n121 ));
    InMux I__2279 (
            .O(N__13646),
            .I(\transmit_module.n3172 ));
    InMux I__2278 (
            .O(N__13643),
            .I(N__13640));
    LocalMux I__2277 (
            .O(N__13640),
            .I(N__13637));
    Odrv4 I__2276 (
            .O(N__13637),
            .I(\transmit_module.n120 ));
    InMux I__2275 (
            .O(N__13634),
            .I(\transmit_module.n3173 ));
    InMux I__2274 (
            .O(N__13631),
            .I(\transmit_module.n3174 ));
    InMux I__2273 (
            .O(N__13628),
            .I(N__13625));
    LocalMux I__2272 (
            .O(N__13625),
            .I(N__13622));
    Span4Mux_h I__2271 (
            .O(N__13622),
            .I(N__13619));
    Odrv4 I__2270 (
            .O(N__13619),
            .I(\transmit_module.n119 ));
    InMux I__2269 (
            .O(N__13616),
            .I(N__13612));
    InMux I__2268 (
            .O(N__13615),
            .I(N__13609));
    LocalMux I__2267 (
            .O(N__13612),
            .I(\transmit_module.n112 ));
    LocalMux I__2266 (
            .O(N__13609),
            .I(\transmit_module.n112 ));
    InMux I__2265 (
            .O(N__13604),
            .I(N__13601));
    LocalMux I__2264 (
            .O(N__13601),
            .I(N__13597));
    InMux I__2263 (
            .O(N__13600),
            .I(N__13594));
    Span4Mux_h I__2262 (
            .O(N__13597),
            .I(N__13591));
    LocalMux I__2261 (
            .O(N__13594),
            .I(\transmit_module.n146 ));
    Odrv4 I__2260 (
            .O(N__13591),
            .I(\transmit_module.n146 ));
    InMux I__2259 (
            .O(N__13586),
            .I(N__13583));
    LocalMux I__2258 (
            .O(N__13583),
            .I(N__13580));
    Odrv12 I__2257 (
            .O(N__13580),
            .I(\sync_buffer.BUFFER_1_0 ));
    InMux I__2256 (
            .O(N__13577),
            .I(N__13574));
    LocalMux I__2255 (
            .O(N__13574),
            .I(N__13571));
    Odrv4 I__2254 (
            .O(N__13571),
            .I(RX_TX_SYNC_BUFF));
    InMux I__2253 (
            .O(N__13568),
            .I(N__13565));
    LocalMux I__2252 (
            .O(N__13565),
            .I(\transmit_module.n122 ));
    CascadeMux I__2251 (
            .O(N__13562),
            .I(\transmit_module.n137_cascade_ ));
    InMux I__2250 (
            .O(N__13559),
            .I(\transmit_module.n3163 ));
    InMux I__2249 (
            .O(N__13556),
            .I(\transmit_module.n3164 ));
    CascadeMux I__2248 (
            .O(N__13553),
            .I(N__13550));
    InMux I__2247 (
            .O(N__13550),
            .I(N__13547));
    LocalMux I__2246 (
            .O(N__13547),
            .I(N__13544));
    Odrv4 I__2245 (
            .O(N__13544),
            .I(\transmit_module.n128 ));
    InMux I__2244 (
            .O(N__13541),
            .I(\transmit_module.n3165 ));
    InMux I__2243 (
            .O(N__13538),
            .I(N__13535));
    LocalMux I__2242 (
            .O(N__13535),
            .I(N__13529));
    InMux I__2241 (
            .O(N__13534),
            .I(N__13526));
    InMux I__2240 (
            .O(N__13533),
            .I(N__13523));
    InMux I__2239 (
            .O(N__13532),
            .I(N__13520));
    Odrv4 I__2238 (
            .O(N__13529),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__2237 (
            .O(N__13526),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__2236 (
            .O(N__13523),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__2235 (
            .O(N__13520),
            .I(\transmit_module.TX_ADDR_5 ));
    CascadeMux I__2234 (
            .O(N__13511),
            .I(N__13508));
    InMux I__2233 (
            .O(N__13508),
            .I(N__13505));
    LocalMux I__2232 (
            .O(N__13505),
            .I(\transmit_module.n127 ));
    InMux I__2231 (
            .O(N__13502),
            .I(\transmit_module.n3166 ));
    InMux I__2230 (
            .O(N__13499),
            .I(N__13496));
    LocalMux I__2229 (
            .O(N__13496),
            .I(\transmit_module.n126 ));
    InMux I__2228 (
            .O(N__13493),
            .I(\transmit_module.n3167 ));
    InMux I__2227 (
            .O(N__13490),
            .I(N__13487));
    LocalMux I__2226 (
            .O(N__13487),
            .I(N__13483));
    CascadeMux I__2225 (
            .O(N__13486),
            .I(N__13479));
    Span4Mux_v I__2224 (
            .O(N__13483),
            .I(N__13475));
    InMux I__2223 (
            .O(N__13482),
            .I(N__13472));
    InMux I__2222 (
            .O(N__13479),
            .I(N__13469));
    InMux I__2221 (
            .O(N__13478),
            .I(N__13466));
    Odrv4 I__2220 (
            .O(N__13475),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__2219 (
            .O(N__13472),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__2218 (
            .O(N__13469),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__2217 (
            .O(N__13466),
            .I(\transmit_module.TX_ADDR_7 ));
    InMux I__2216 (
            .O(N__13457),
            .I(N__13454));
    LocalMux I__2215 (
            .O(N__13454),
            .I(\transmit_module.n125 ));
    InMux I__2214 (
            .O(N__13451),
            .I(\transmit_module.n3168 ));
    InMux I__2213 (
            .O(N__13448),
            .I(N__13445));
    LocalMux I__2212 (
            .O(N__13445),
            .I(N__13442));
    Odrv4 I__2211 (
            .O(N__13442),
            .I(\transmit_module.n124 ));
    InMux I__2210 (
            .O(N__13439),
            .I(bfn_14_16_0_));
    InMux I__2209 (
            .O(N__13436),
            .I(N__13433));
    LocalMux I__2208 (
            .O(N__13433),
            .I(N__13430));
    Span4Mux_v I__2207 (
            .O(N__13430),
            .I(N__13427));
    Odrv4 I__2206 (
            .O(N__13427),
            .I(\transmit_module.n123 ));
    InMux I__2205 (
            .O(N__13424),
            .I(\transmit_module.n3170 ));
    InMux I__2204 (
            .O(N__13421),
            .I(\transmit_module.n3171 ));
    SRMux I__2203 (
            .O(N__13418),
            .I(N__13415));
    LocalMux I__2202 (
            .O(N__13415),
            .I(N__13410));
    SRMux I__2201 (
            .O(N__13414),
            .I(N__13407));
    SRMux I__2200 (
            .O(N__13413),
            .I(N__13404));
    Span4Mux_s2_v I__2199 (
            .O(N__13410),
            .I(N__13396));
    LocalMux I__2198 (
            .O(N__13407),
            .I(N__13396));
    LocalMux I__2197 (
            .O(N__13404),
            .I(N__13396));
    SRMux I__2196 (
            .O(N__13403),
            .I(N__13393));
    Span4Mux_v I__2195 (
            .O(N__13396),
            .I(N__13390));
    LocalMux I__2194 (
            .O(N__13393),
            .I(N__13387));
    Sp12to4 I__2193 (
            .O(N__13390),
            .I(N__13384));
    Span4Mux_h I__2192 (
            .O(N__13387),
            .I(N__13381));
    Span12Mux_v I__2191 (
            .O(N__13384),
            .I(N__13378));
    Span4Mux_h I__2190 (
            .O(N__13381),
            .I(N__13375));
    Odrv12 I__2189 (
            .O(N__13378),
            .I(\line_buffer.n605 ));
    Odrv4 I__2188 (
            .O(N__13375),
            .I(\line_buffer.n605 ));
    InMux I__2187 (
            .O(N__13370),
            .I(N__13367));
    LocalMux I__2186 (
            .O(N__13367),
            .I(N__13364));
    Span4Mux_h I__2185 (
            .O(N__13364),
            .I(N__13361));
    Span4Mux_h I__2184 (
            .O(N__13361),
            .I(N__13358));
    Span4Mux_v I__2183 (
            .O(N__13358),
            .I(N__13355));
    Odrv4 I__2182 (
            .O(N__13355),
            .I(\line_buffer.n568 ));
    InMux I__2181 (
            .O(N__13352),
            .I(N__13349));
    LocalMux I__2180 (
            .O(N__13349),
            .I(N__13346));
    Span4Mux_h I__2179 (
            .O(N__13346),
            .I(N__13343));
    Span4Mux_h I__2178 (
            .O(N__13343),
            .I(N__13340));
    Odrv4 I__2177 (
            .O(N__13340),
            .I(\line_buffer.n560 ));
    InMux I__2176 (
            .O(N__13337),
            .I(N__13334));
    LocalMux I__2175 (
            .O(N__13334),
            .I(\sync_buffer.BUFFER_0_0 ));
    InMux I__2174 (
            .O(N__13331),
            .I(N__13328));
    LocalMux I__2173 (
            .O(N__13328),
            .I(N__13325));
    Odrv4 I__2172 (
            .O(N__13325),
            .I(\transmit_module.ADDR_Y_COMPONENT_6 ));
    InMux I__2171 (
            .O(N__13322),
            .I(N__13319));
    LocalMux I__2170 (
            .O(N__13319),
            .I(\transmit_module.n131 ));
    InMux I__2169 (
            .O(N__13316),
            .I(\transmit_module.n3162 ));
    CascadeMux I__2168 (
            .O(N__13313),
            .I(\receive_module.rx_counter.n5_cascade_ ));
    InMux I__2167 (
            .O(N__13310),
            .I(N__13306));
    InMux I__2166 (
            .O(N__13309),
            .I(N__13301));
    LocalMux I__2165 (
            .O(N__13306),
            .I(N__13298));
    InMux I__2164 (
            .O(N__13305),
            .I(N__13293));
    InMux I__2163 (
            .O(N__13304),
            .I(N__13293));
    LocalMux I__2162 (
            .O(N__13301),
            .I(\receive_module.rx_counter.Y_7 ));
    Odrv4 I__2161 (
            .O(N__13298),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__2160 (
            .O(N__13293),
            .I(\receive_module.rx_counter.Y_7 ));
    CascadeMux I__2159 (
            .O(N__13286),
            .I(\receive_module.rx_counter.n3455_cascade_ ));
    InMux I__2158 (
            .O(N__13283),
            .I(N__13280));
    LocalMux I__2157 (
            .O(N__13280),
            .I(N__13276));
    InMux I__2156 (
            .O(N__13279),
            .I(N__13273));
    Odrv4 I__2155 (
            .O(N__13276),
            .I(\receive_module.rx_counter.n3680 ));
    LocalMux I__2154 (
            .O(N__13273),
            .I(\receive_module.rx_counter.n3680 ));
    CascadeMux I__2153 (
            .O(N__13268),
            .I(N__13265));
    InMux I__2152 (
            .O(N__13265),
            .I(N__13259));
    InMux I__2151 (
            .O(N__13264),
            .I(N__13256));
    InMux I__2150 (
            .O(N__13263),
            .I(N__13253));
    InMux I__2149 (
            .O(N__13262),
            .I(N__13250));
    LocalMux I__2148 (
            .O(N__13259),
            .I(N__13247));
    LocalMux I__2147 (
            .O(N__13256),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__2146 (
            .O(N__13253),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__2145 (
            .O(N__13250),
            .I(\receive_module.rx_counter.Y_8 ));
    Odrv4 I__2144 (
            .O(N__13247),
            .I(\receive_module.rx_counter.Y_8 ));
    InMux I__2143 (
            .O(N__13238),
            .I(N__13235));
    LocalMux I__2142 (
            .O(N__13235),
            .I(\receive_module.rx_counter.n3481 ));
    CascadeMux I__2141 (
            .O(N__13232),
            .I(\receive_module.rx_counter.n4_adj_612_cascade_ ));
    InMux I__2140 (
            .O(N__13229),
            .I(N__13226));
    LocalMux I__2139 (
            .O(N__13226),
            .I(\receive_module.rx_counter.n54 ));
    InMux I__2138 (
            .O(N__13223),
            .I(N__13220));
    LocalMux I__2137 (
            .O(N__13220),
            .I(N__13214));
    InMux I__2136 (
            .O(N__13219),
            .I(N__13211));
    InMux I__2135 (
            .O(N__13218),
            .I(N__13206));
    InMux I__2134 (
            .O(N__13217),
            .I(N__13206));
    Odrv4 I__2133 (
            .O(N__13214),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__2132 (
            .O(N__13211),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__2131 (
            .O(N__13206),
            .I(\receive_module.rx_counter.Y_1 ));
    InMux I__2130 (
            .O(N__13199),
            .I(N__13195));
    CascadeMux I__2129 (
            .O(N__13198),
            .I(N__13190));
    LocalMux I__2128 (
            .O(N__13195),
            .I(N__13187));
    InMux I__2127 (
            .O(N__13194),
            .I(N__13184));
    InMux I__2126 (
            .O(N__13193),
            .I(N__13181));
    InMux I__2125 (
            .O(N__13190),
            .I(N__13178));
    Odrv4 I__2124 (
            .O(N__13187),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__2123 (
            .O(N__13184),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__2122 (
            .O(N__13181),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__2121 (
            .O(N__13178),
            .I(\receive_module.rx_counter.Y_0 ));
    InMux I__2120 (
            .O(N__13169),
            .I(N__13166));
    LocalMux I__2119 (
            .O(N__13166),
            .I(N__13160));
    InMux I__2118 (
            .O(N__13165),
            .I(N__13157));
    InMux I__2117 (
            .O(N__13164),
            .I(N__13152));
    InMux I__2116 (
            .O(N__13163),
            .I(N__13152));
    Odrv4 I__2115 (
            .O(N__13160),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__2114 (
            .O(N__13157),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__2113 (
            .O(N__13152),
            .I(\receive_module.rx_counter.Y_2 ));
    InMux I__2112 (
            .O(N__13145),
            .I(N__13142));
    LocalMux I__2111 (
            .O(N__13142),
            .I(\receive_module.rx_counter.n3453 ));
    InMux I__2110 (
            .O(N__13139),
            .I(N__13136));
    LocalMux I__2109 (
            .O(N__13136),
            .I(N__13130));
    InMux I__2108 (
            .O(N__13135),
            .I(N__13127));
    InMux I__2107 (
            .O(N__13134),
            .I(N__13122));
    InMux I__2106 (
            .O(N__13133),
            .I(N__13122));
    Odrv4 I__2105 (
            .O(N__13130),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__2104 (
            .O(N__13127),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__2103 (
            .O(N__13122),
            .I(\receive_module.rx_counter.Y_3 ));
    InMux I__2102 (
            .O(N__13115),
            .I(N__13111));
    InMux I__2101 (
            .O(N__13114),
            .I(N__13106));
    LocalMux I__2100 (
            .O(N__13111),
            .I(N__13103));
    InMux I__2099 (
            .O(N__13110),
            .I(N__13100));
    InMux I__2098 (
            .O(N__13109),
            .I(N__13097));
    LocalMux I__2097 (
            .O(N__13106),
            .I(\receive_module.rx_counter.Y_4 ));
    Odrv4 I__2096 (
            .O(N__13103),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__2095 (
            .O(N__13100),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__2094 (
            .O(N__13097),
            .I(\receive_module.rx_counter.Y_4 ));
    InMux I__2093 (
            .O(N__13088),
            .I(N__13085));
    LocalMux I__2092 (
            .O(N__13085),
            .I(\receive_module.rx_counter.n4 ));
    InMux I__2091 (
            .O(N__13082),
            .I(N__13079));
    LocalMux I__2090 (
            .O(N__13079),
            .I(RX_TX_SYNC));
    SRMux I__2089 (
            .O(N__13076),
            .I(N__13073));
    LocalMux I__2088 (
            .O(N__13073),
            .I(N__13068));
    SRMux I__2087 (
            .O(N__13072),
            .I(N__13065));
    SRMux I__2086 (
            .O(N__13071),
            .I(N__13062));
    Span4Mux_v I__2085 (
            .O(N__13068),
            .I(N__13054));
    LocalMux I__2084 (
            .O(N__13065),
            .I(N__13054));
    LocalMux I__2083 (
            .O(N__13062),
            .I(N__13054));
    SRMux I__2082 (
            .O(N__13061),
            .I(N__13051));
    Span4Mux_v I__2081 (
            .O(N__13054),
            .I(N__13048));
    LocalMux I__2080 (
            .O(N__13051),
            .I(N__13045));
    Span4Mux_h I__2079 (
            .O(N__13048),
            .I(N__13040));
    Span4Mux_h I__2078 (
            .O(N__13045),
            .I(N__13040));
    Span4Mux_h I__2077 (
            .O(N__13040),
            .I(N__13037));
    Span4Mux_h I__2076 (
            .O(N__13037),
            .I(N__13034));
    Span4Mux_v I__2075 (
            .O(N__13034),
            .I(N__13031));
    Odrv4 I__2074 (
            .O(N__13031),
            .I(\line_buffer.n477 ));
    SRMux I__2073 (
            .O(N__13028),
            .I(N__13025));
    LocalMux I__2072 (
            .O(N__13025),
            .I(N__13021));
    SRMux I__2071 (
            .O(N__13024),
            .I(N__13018));
    Span4Mux_v I__2070 (
            .O(N__13021),
            .I(N__13011));
    LocalMux I__2069 (
            .O(N__13018),
            .I(N__13011));
    SRMux I__2068 (
            .O(N__13017),
            .I(N__13008));
    SRMux I__2067 (
            .O(N__13016),
            .I(N__13005));
    Span4Mux_v I__2066 (
            .O(N__13011),
            .I(N__12998));
    LocalMux I__2065 (
            .O(N__13008),
            .I(N__12998));
    LocalMux I__2064 (
            .O(N__13005),
            .I(N__12998));
    Span4Mux_v I__2063 (
            .O(N__12998),
            .I(N__12995));
    Sp12to4 I__2062 (
            .O(N__12995),
            .I(N__12992));
    Odrv12 I__2061 (
            .O(N__12992),
            .I(\line_buffer.n541 ));
    InMux I__2060 (
            .O(N__12989),
            .I(N__12984));
    InMux I__2059 (
            .O(N__12988),
            .I(N__12981));
    InMux I__2058 (
            .O(N__12987),
            .I(N__12978));
    LocalMux I__2057 (
            .O(N__12984),
            .I(\receive_module.rx_counter.X_3 ));
    LocalMux I__2056 (
            .O(N__12981),
            .I(\receive_module.rx_counter.X_3 ));
    LocalMux I__2055 (
            .O(N__12978),
            .I(\receive_module.rx_counter.X_3 ));
    InMux I__2054 (
            .O(N__12971),
            .I(N__12966));
    InMux I__2053 (
            .O(N__12970),
            .I(N__12963));
    InMux I__2052 (
            .O(N__12969),
            .I(N__12960));
    LocalMux I__2051 (
            .O(N__12966),
            .I(\receive_module.rx_counter.X_5 ));
    LocalMux I__2050 (
            .O(N__12963),
            .I(\receive_module.rx_counter.X_5 ));
    LocalMux I__2049 (
            .O(N__12960),
            .I(\receive_module.rx_counter.X_5 ));
    InMux I__2048 (
            .O(N__12953),
            .I(N__12948));
    InMux I__2047 (
            .O(N__12952),
            .I(N__12945));
    InMux I__2046 (
            .O(N__12951),
            .I(N__12942));
    LocalMux I__2045 (
            .O(N__12948),
            .I(\receive_module.rx_counter.X_7 ));
    LocalMux I__2044 (
            .O(N__12945),
            .I(\receive_module.rx_counter.X_7 ));
    LocalMux I__2043 (
            .O(N__12942),
            .I(\receive_module.rx_counter.X_7 ));
    InMux I__2042 (
            .O(N__12935),
            .I(N__12932));
    LocalMux I__2041 (
            .O(N__12932),
            .I(\receive_module.rx_counter.n6 ));
    CascadeMux I__2040 (
            .O(N__12929),
            .I(\receive_module.rx_counter.n7_cascade_ ));
    InMux I__2039 (
            .O(N__12926),
            .I(N__12923));
    LocalMux I__2038 (
            .O(N__12923),
            .I(\receive_module.rx_counter.n3225 ));
    InMux I__2037 (
            .O(N__12920),
            .I(N__12917));
    LocalMux I__2036 (
            .O(N__12917),
            .I(\receive_module.rx_counter.old_HS ));
    CEMux I__2035 (
            .O(N__12914),
            .I(N__12910));
    CEMux I__2034 (
            .O(N__12913),
            .I(N__12907));
    LocalMux I__2033 (
            .O(N__12910),
            .I(\receive_module.rx_counter.n2081 ));
    LocalMux I__2032 (
            .O(N__12907),
            .I(\receive_module.rx_counter.n2081 ));
    SRMux I__2031 (
            .O(N__12902),
            .I(N__12897));
    SRMux I__2030 (
            .O(N__12901),
            .I(N__12894));
    SRMux I__2029 (
            .O(N__12900),
            .I(N__12891));
    LocalMux I__2028 (
            .O(N__12897),
            .I(N__12887));
    LocalMux I__2027 (
            .O(N__12894),
            .I(N__12882));
    LocalMux I__2026 (
            .O(N__12891),
            .I(N__12882));
    SRMux I__2025 (
            .O(N__12890),
            .I(N__12879));
    Span4Mux_v I__2024 (
            .O(N__12887),
            .I(N__12876));
    Span4Mux_v I__2023 (
            .O(N__12882),
            .I(N__12871));
    LocalMux I__2022 (
            .O(N__12879),
            .I(N__12871));
    Span4Mux_v I__2021 (
            .O(N__12876),
            .I(N__12866));
    Span4Mux_v I__2020 (
            .O(N__12871),
            .I(N__12866));
    Sp12to4 I__2019 (
            .O(N__12866),
            .I(N__12863));
    Odrv12 I__2018 (
            .O(N__12863),
            .I(\line_buffer.n573 ));
    InMux I__2017 (
            .O(N__12860),
            .I(N__12857));
    LocalMux I__2016 (
            .O(N__12857),
            .I(\receive_module.rx_counter.n3429 ));
    InMux I__2015 (
            .O(N__12854),
            .I(N__12849));
    InMux I__2014 (
            .O(N__12853),
            .I(N__12846));
    InMux I__2013 (
            .O(N__12852),
            .I(N__12843));
    LocalMux I__2012 (
            .O(N__12849),
            .I(\receive_module.rx_counter.X_8 ));
    LocalMux I__2011 (
            .O(N__12846),
            .I(\receive_module.rx_counter.X_8 ));
    LocalMux I__2010 (
            .O(N__12843),
            .I(\receive_module.rx_counter.X_8 ));
    CascadeMux I__2009 (
            .O(N__12836),
            .I(N__12832));
    InMux I__2008 (
            .O(N__12835),
            .I(N__12829));
    InMux I__2007 (
            .O(N__12832),
            .I(N__12826));
    LocalMux I__2006 (
            .O(N__12829),
            .I(\receive_module.rx_counter.X_9 ));
    LocalMux I__2005 (
            .O(N__12826),
            .I(\receive_module.rx_counter.X_9 ));
    InMux I__2004 (
            .O(N__12821),
            .I(N__12818));
    LocalMux I__2003 (
            .O(N__12818),
            .I(N__12815));
    Odrv4 I__2002 (
            .O(N__12815),
            .I(\receive_module.rx_counter.n39 ));
    InMux I__2001 (
            .O(N__12812),
            .I(N__12807));
    InMux I__2000 (
            .O(N__12811),
            .I(N__12804));
    InMux I__1999 (
            .O(N__12810),
            .I(N__12801));
    LocalMux I__1998 (
            .O(N__12807),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__1997 (
            .O(N__12804),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__1996 (
            .O(N__12801),
            .I(\receive_module.rx_counter.Y_6 ));
    InMux I__1995 (
            .O(N__12794),
            .I(N__12789));
    InMux I__1994 (
            .O(N__12793),
            .I(N__12786));
    InMux I__1993 (
            .O(N__12792),
            .I(N__12783));
    LocalMux I__1992 (
            .O(N__12789),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__1991 (
            .O(N__12786),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__1990 (
            .O(N__12783),
            .I(\receive_module.rx_counter.Y_5 ));
    InMux I__1989 (
            .O(N__12776),
            .I(N__12773));
    LocalMux I__1988 (
            .O(N__12773),
            .I(N__12770));
    Span4Mux_h I__1987 (
            .O(N__12770),
            .I(N__12767));
    Span4Mux_h I__1986 (
            .O(N__12767),
            .I(N__12764));
    Odrv4 I__1985 (
            .O(N__12764),
            .I(\line_buffer.n571 ));
    InMux I__1984 (
            .O(N__12761),
            .I(N__12758));
    LocalMux I__1983 (
            .O(N__12758),
            .I(N__12755));
    Span12Mux_v I__1982 (
            .O(N__12755),
            .I(N__12752));
    Span12Mux_v I__1981 (
            .O(N__12752),
            .I(N__12749));
    Span12Mux_h I__1980 (
            .O(N__12749),
            .I(N__12746));
    Odrv12 I__1979 (
            .O(N__12746),
            .I(\line_buffer.n563 ));
    InMux I__1978 (
            .O(N__12743),
            .I(N__12740));
    LocalMux I__1977 (
            .O(N__12740),
            .I(\line_buffer.n3534 ));
    InMux I__1976 (
            .O(N__12737),
            .I(N__12734));
    LocalMux I__1975 (
            .O(N__12734),
            .I(N__12731));
    Odrv4 I__1974 (
            .O(N__12731),
            .I(TX_DATA_7));
    IoInMux I__1973 (
            .O(N__12728),
            .I(N__12723));
    IoInMux I__1972 (
            .O(N__12727),
            .I(N__12720));
    IoInMux I__1971 (
            .O(N__12726),
            .I(N__12717));
    LocalMux I__1970 (
            .O(N__12723),
            .I(N__12714));
    LocalMux I__1969 (
            .O(N__12720),
            .I(N__12711));
    LocalMux I__1968 (
            .O(N__12717),
            .I(N__12708));
    IoSpan4Mux I__1967 (
            .O(N__12714),
            .I(N__12705));
    IoSpan4Mux I__1966 (
            .O(N__12711),
            .I(N__12702));
    Span12Mux_s8_v I__1965 (
            .O(N__12708),
            .I(N__12699));
    Sp12to4 I__1964 (
            .O(N__12705),
            .I(N__12696));
    Span4Mux_s2_v I__1963 (
            .O(N__12702),
            .I(N__12693));
    Span12Mux_h I__1962 (
            .O(N__12699),
            .I(N__12690));
    Span12Mux_h I__1961 (
            .O(N__12696),
            .I(N__12687));
    Sp12to4 I__1960 (
            .O(N__12693),
            .I(N__12684));
    Odrv12 I__1959 (
            .O(N__12690),
            .I(ADV_B_c));
    Odrv12 I__1958 (
            .O(N__12687),
            .I(ADV_B_c));
    Odrv12 I__1957 (
            .O(N__12684),
            .I(ADV_B_c));
    InMux I__1956 (
            .O(N__12677),
            .I(N__12674));
    LocalMux I__1955 (
            .O(N__12674),
            .I(N__12671));
    Span12Mux_h I__1954 (
            .O(N__12671),
            .I(N__12668));
    Odrv12 I__1953 (
            .O(N__12668),
            .I(\line_buffer.n474 ));
    InMux I__1952 (
            .O(N__12665),
            .I(N__12662));
    LocalMux I__1951 (
            .O(N__12662),
            .I(N__12659));
    Span4Mux_h I__1950 (
            .O(N__12659),
            .I(N__12656));
    Span4Mux_h I__1949 (
            .O(N__12656),
            .I(N__12653));
    Odrv4 I__1948 (
            .O(N__12653),
            .I(\line_buffer.n466 ));
    InMux I__1947 (
            .O(N__12650),
            .I(N__12647));
    LocalMux I__1946 (
            .O(N__12647),
            .I(N__12644));
    Odrv12 I__1945 (
            .O(N__12644),
            .I(\line_buffer.n3533 ));
    SRMux I__1944 (
            .O(N__12641),
            .I(N__12636));
    SRMux I__1943 (
            .O(N__12640),
            .I(N__12633));
    SRMux I__1942 (
            .O(N__12639),
            .I(N__12630));
    LocalMux I__1941 (
            .O(N__12636),
            .I(N__12627));
    LocalMux I__1940 (
            .O(N__12633),
            .I(N__12623));
    LocalMux I__1939 (
            .O(N__12630),
            .I(N__12620));
    Span4Mux_h I__1938 (
            .O(N__12627),
            .I(N__12617));
    SRMux I__1937 (
            .O(N__12626),
            .I(N__12614));
    Span4Mux_v I__1936 (
            .O(N__12623),
            .I(N__12611));
    Span4Mux_h I__1935 (
            .O(N__12620),
            .I(N__12608));
    Span4Mux_v I__1934 (
            .O(N__12617),
            .I(N__12603));
    LocalMux I__1933 (
            .O(N__12614),
            .I(N__12603));
    Sp12to4 I__1932 (
            .O(N__12611),
            .I(N__12600));
    Span4Mux_h I__1931 (
            .O(N__12608),
            .I(N__12597));
    Span4Mux_h I__1930 (
            .O(N__12603),
            .I(N__12594));
    Span12Mux_v I__1929 (
            .O(N__12600),
            .I(N__12591));
    Span4Mux_v I__1928 (
            .O(N__12597),
            .I(N__12588));
    Span4Mux_h I__1927 (
            .O(N__12594),
            .I(N__12585));
    Odrv12 I__1926 (
            .O(N__12591),
            .I(\line_buffer.n542 ));
    Odrv4 I__1925 (
            .O(N__12588),
            .I(\line_buffer.n542 ));
    Odrv4 I__1924 (
            .O(N__12585),
            .I(\line_buffer.n542 ));
    InMux I__1923 (
            .O(N__12578),
            .I(N__12574));
    InMux I__1922 (
            .O(N__12577),
            .I(N__12571));
    LocalMux I__1921 (
            .O(N__12574),
            .I(\receive_module.rx_counter.X_1 ));
    LocalMux I__1920 (
            .O(N__12571),
            .I(\receive_module.rx_counter.X_1 ));
    InMux I__1919 (
            .O(N__12566),
            .I(N__12562));
    InMux I__1918 (
            .O(N__12565),
            .I(N__12559));
    LocalMux I__1917 (
            .O(N__12562),
            .I(\receive_module.rx_counter.X_0 ));
    LocalMux I__1916 (
            .O(N__12559),
            .I(\receive_module.rx_counter.X_0 ));
    InMux I__1915 (
            .O(N__12554),
            .I(N__12550));
    InMux I__1914 (
            .O(N__12553),
            .I(N__12547));
    LocalMux I__1913 (
            .O(N__12550),
            .I(\receive_module.rx_counter.X_2 ));
    LocalMux I__1912 (
            .O(N__12547),
            .I(\receive_module.rx_counter.X_2 ));
    CascadeMux I__1911 (
            .O(N__12542),
            .I(\receive_module.rx_counter.n3225_cascade_ ));
    CascadeMux I__1910 (
            .O(N__12539),
            .I(\receive_module.rx_counter.n3458_cascade_ ));
    InMux I__1909 (
            .O(N__12536),
            .I(N__12531));
    InMux I__1908 (
            .O(N__12535),
            .I(N__12526));
    InMux I__1907 (
            .O(N__12534),
            .I(N__12526));
    LocalMux I__1906 (
            .O(N__12531),
            .I(\receive_module.rx_counter.X_4 ));
    LocalMux I__1905 (
            .O(N__12526),
            .I(\receive_module.rx_counter.X_4 ));
    InMux I__1904 (
            .O(N__12521),
            .I(N__12516));
    InMux I__1903 (
            .O(N__12520),
            .I(N__12511));
    InMux I__1902 (
            .O(N__12519),
            .I(N__12511));
    LocalMux I__1901 (
            .O(N__12516),
            .I(\receive_module.rx_counter.X_6 ));
    LocalMux I__1900 (
            .O(N__12511),
            .I(\receive_module.rx_counter.X_6 ));
    SRMux I__1899 (
            .O(N__12506),
            .I(N__12503));
    LocalMux I__1898 (
            .O(N__12503),
            .I(N__12499));
    SRMux I__1897 (
            .O(N__12502),
            .I(N__12496));
    Span4Mux_h I__1896 (
            .O(N__12499),
            .I(N__12493));
    LocalMux I__1895 (
            .O(N__12496),
            .I(N__12490));
    Odrv4 I__1894 (
            .O(N__12493),
            .I(\receive_module.rx_counter.n3 ));
    Odrv12 I__1893 (
            .O(N__12490),
            .I(\receive_module.rx_counter.n3 ));
    InMux I__1892 (
            .O(N__12485),
            .I(N__12480));
    InMux I__1891 (
            .O(N__12484),
            .I(N__12477));
    CascadeMux I__1890 (
            .O(N__12483),
            .I(N__12474));
    LocalMux I__1889 (
            .O(N__12480),
            .I(N__12468));
    LocalMux I__1888 (
            .O(N__12477),
            .I(N__12468));
    InMux I__1887 (
            .O(N__12474),
            .I(N__12463));
    InMux I__1886 (
            .O(N__12473),
            .I(N__12463));
    Odrv4 I__1885 (
            .O(N__12468),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__1884 (
            .O(N__12463),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    InMux I__1883 (
            .O(N__12458),
            .I(N__12452));
    InMux I__1882 (
            .O(N__12457),
            .I(N__12449));
    InMux I__1881 (
            .O(N__12456),
            .I(N__12444));
    InMux I__1880 (
            .O(N__12455),
            .I(N__12444));
    LocalMux I__1879 (
            .O(N__12452),
            .I(N__12439));
    LocalMux I__1878 (
            .O(N__12449),
            .I(N__12439));
    LocalMux I__1877 (
            .O(N__12444),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    Odrv4 I__1876 (
            .O(N__12439),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    InMux I__1875 (
            .O(N__12434),
            .I(N__12431));
    LocalMux I__1874 (
            .O(N__12431),
            .I(\transmit_module.video_signal_controller.n3679 ));
    InMux I__1873 (
            .O(N__12428),
            .I(N__12424));
    InMux I__1872 (
            .O(N__12427),
            .I(N__12421));
    LocalMux I__1871 (
            .O(N__12424),
            .I(\transmit_module.n108 ));
    LocalMux I__1870 (
            .O(N__12421),
            .I(\transmit_module.n108 ));
    InMux I__1869 (
            .O(N__12416),
            .I(N__12412));
    InMux I__1868 (
            .O(N__12415),
            .I(N__12409));
    LocalMux I__1867 (
            .O(N__12412),
            .I(N__12403));
    LocalMux I__1866 (
            .O(N__12409),
            .I(N__12400));
    InMux I__1865 (
            .O(N__12408),
            .I(N__12397));
    InMux I__1864 (
            .O(N__12407),
            .I(N__12394));
    InMux I__1863 (
            .O(N__12406),
            .I(N__12391));
    Span4Mux_v I__1862 (
            .O(N__12403),
            .I(N__12384));
    Span4Mux_v I__1861 (
            .O(N__12400),
            .I(N__12384));
    LocalMux I__1860 (
            .O(N__12397),
            .I(N__12384));
    LocalMux I__1859 (
            .O(N__12394),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    LocalMux I__1858 (
            .O(N__12391),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__1857 (
            .O(N__12384),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    InMux I__1856 (
            .O(N__12377),
            .I(N__12374));
    LocalMux I__1855 (
            .O(N__12374),
            .I(\transmit_module.video_signal_controller.n6_adj_623 ));
    InMux I__1854 (
            .O(N__12371),
            .I(N__12367));
    InMux I__1853 (
            .O(N__12370),
            .I(N__12364));
    LocalMux I__1852 (
            .O(N__12367),
            .I(\transmit_module.n139 ));
    LocalMux I__1851 (
            .O(N__12364),
            .I(\transmit_module.n139 ));
    CascadeMux I__1850 (
            .O(N__12359),
            .I(\transmit_module.n138_cascade_ ));
    CascadeMux I__1849 (
            .O(N__12356),
            .I(N__12352));
    CascadeMux I__1848 (
            .O(N__12355),
            .I(N__12349));
    CascadeBuf I__1847 (
            .O(N__12352),
            .I(N__12346));
    CascadeBuf I__1846 (
            .O(N__12349),
            .I(N__12343));
    CascadeMux I__1845 (
            .O(N__12346),
            .I(N__12340));
    CascadeMux I__1844 (
            .O(N__12343),
            .I(N__12337));
    CascadeBuf I__1843 (
            .O(N__12340),
            .I(N__12334));
    CascadeBuf I__1842 (
            .O(N__12337),
            .I(N__12331));
    CascadeMux I__1841 (
            .O(N__12334),
            .I(N__12328));
    CascadeMux I__1840 (
            .O(N__12331),
            .I(N__12325));
    CascadeBuf I__1839 (
            .O(N__12328),
            .I(N__12322));
    CascadeBuf I__1838 (
            .O(N__12325),
            .I(N__12319));
    CascadeMux I__1837 (
            .O(N__12322),
            .I(N__12316));
    CascadeMux I__1836 (
            .O(N__12319),
            .I(N__12313));
    CascadeBuf I__1835 (
            .O(N__12316),
            .I(N__12310));
    CascadeBuf I__1834 (
            .O(N__12313),
            .I(N__12307));
    CascadeMux I__1833 (
            .O(N__12310),
            .I(N__12304));
    CascadeMux I__1832 (
            .O(N__12307),
            .I(N__12301));
    CascadeBuf I__1831 (
            .O(N__12304),
            .I(N__12298));
    CascadeBuf I__1830 (
            .O(N__12301),
            .I(N__12295));
    CascadeMux I__1829 (
            .O(N__12298),
            .I(N__12292));
    CascadeMux I__1828 (
            .O(N__12295),
            .I(N__12289));
    CascadeBuf I__1827 (
            .O(N__12292),
            .I(N__12286));
    CascadeBuf I__1826 (
            .O(N__12289),
            .I(N__12283));
    CascadeMux I__1825 (
            .O(N__12286),
            .I(N__12280));
    CascadeMux I__1824 (
            .O(N__12283),
            .I(N__12277));
    CascadeBuf I__1823 (
            .O(N__12280),
            .I(N__12274));
    CascadeBuf I__1822 (
            .O(N__12277),
            .I(N__12271));
    CascadeMux I__1821 (
            .O(N__12274),
            .I(N__12268));
    CascadeMux I__1820 (
            .O(N__12271),
            .I(N__12265));
    CascadeBuf I__1819 (
            .O(N__12268),
            .I(N__12262));
    CascadeBuf I__1818 (
            .O(N__12265),
            .I(N__12259));
    CascadeMux I__1817 (
            .O(N__12262),
            .I(N__12256));
    CascadeMux I__1816 (
            .O(N__12259),
            .I(N__12253));
    CascadeBuf I__1815 (
            .O(N__12256),
            .I(N__12250));
    CascadeBuf I__1814 (
            .O(N__12253),
            .I(N__12247));
    CascadeMux I__1813 (
            .O(N__12250),
            .I(N__12244));
    CascadeMux I__1812 (
            .O(N__12247),
            .I(N__12241));
    CascadeBuf I__1811 (
            .O(N__12244),
            .I(N__12238));
    CascadeBuf I__1810 (
            .O(N__12241),
            .I(N__12235));
    CascadeMux I__1809 (
            .O(N__12238),
            .I(N__12232));
    CascadeMux I__1808 (
            .O(N__12235),
            .I(N__12229));
    CascadeBuf I__1807 (
            .O(N__12232),
            .I(N__12226));
    CascadeBuf I__1806 (
            .O(N__12229),
            .I(N__12223));
    CascadeMux I__1805 (
            .O(N__12226),
            .I(N__12220));
    CascadeMux I__1804 (
            .O(N__12223),
            .I(N__12217));
    CascadeBuf I__1803 (
            .O(N__12220),
            .I(N__12214));
    CascadeBuf I__1802 (
            .O(N__12217),
            .I(N__12211));
    CascadeMux I__1801 (
            .O(N__12214),
            .I(N__12208));
    CascadeMux I__1800 (
            .O(N__12211),
            .I(N__12205));
    CascadeBuf I__1799 (
            .O(N__12208),
            .I(N__12202));
    CascadeBuf I__1798 (
            .O(N__12205),
            .I(N__12199));
    CascadeMux I__1797 (
            .O(N__12202),
            .I(N__12196));
    CascadeMux I__1796 (
            .O(N__12199),
            .I(N__12193));
    CascadeBuf I__1795 (
            .O(N__12196),
            .I(N__12190));
    CascadeBuf I__1794 (
            .O(N__12193),
            .I(N__12187));
    CascadeMux I__1793 (
            .O(N__12190),
            .I(N__12184));
    CascadeMux I__1792 (
            .O(N__12187),
            .I(N__12181));
    CascadeBuf I__1791 (
            .O(N__12184),
            .I(N__12178));
    CascadeBuf I__1790 (
            .O(N__12181),
            .I(N__12175));
    CascadeMux I__1789 (
            .O(N__12178),
            .I(N__12172));
    CascadeMux I__1788 (
            .O(N__12175),
            .I(N__12169));
    InMux I__1787 (
            .O(N__12172),
            .I(N__12166));
    InMux I__1786 (
            .O(N__12169),
            .I(N__12163));
    LocalMux I__1785 (
            .O(N__12166),
            .I(N__12160));
    LocalMux I__1784 (
            .O(N__12163),
            .I(N__12157));
    Span12Mux_s7_v I__1783 (
            .O(N__12160),
            .I(N__12154));
    Span12Mux_h I__1782 (
            .O(N__12157),
            .I(N__12151));
    Span12Mux_h I__1781 (
            .O(N__12154),
            .I(N__12148));
    Span12Mux_v I__1780 (
            .O(N__12151),
            .I(N__12145));
    Odrv12 I__1779 (
            .O(N__12148),
            .I(n19));
    Odrv12 I__1778 (
            .O(N__12145),
            .I(n19));
    InMux I__1777 (
            .O(N__12140),
            .I(N__12137));
    LocalMux I__1776 (
            .O(N__12137),
            .I(N__12134));
    Odrv12 I__1775 (
            .O(N__12134),
            .I(\line_buffer.n3531 ));
    InMux I__1774 (
            .O(N__12131),
            .I(N__12128));
    LocalMux I__1773 (
            .O(N__12128),
            .I(N__12125));
    Span4Mux_v I__1772 (
            .O(N__12125),
            .I(N__12122));
    Odrv4 I__1771 (
            .O(N__12122),
            .I(\line_buffer.n3530 ));
    InMux I__1770 (
            .O(N__12119),
            .I(N__12116));
    LocalMux I__1769 (
            .O(N__12116),
            .I(\line_buffer.n3620 ));
    InMux I__1768 (
            .O(N__12113),
            .I(N__12110));
    LocalMux I__1767 (
            .O(N__12110),
            .I(\transmit_module.n142 ));
    CascadeMux I__1766 (
            .O(N__12107),
            .I(\transmit_module.n142_cascade_ ));
    InMux I__1765 (
            .O(N__12104),
            .I(N__12098));
    InMux I__1764 (
            .O(N__12103),
            .I(N__12098));
    LocalMux I__1763 (
            .O(N__12098),
            .I(\transmit_module.n111 ));
    CascadeMux I__1762 (
            .O(N__12095),
            .I(N__12092));
    CascadeBuf I__1761 (
            .O(N__12092),
            .I(N__12088));
    CascadeMux I__1760 (
            .O(N__12091),
            .I(N__12085));
    CascadeMux I__1759 (
            .O(N__12088),
            .I(N__12082));
    CascadeBuf I__1758 (
            .O(N__12085),
            .I(N__12079));
    CascadeBuf I__1757 (
            .O(N__12082),
            .I(N__12076));
    CascadeMux I__1756 (
            .O(N__12079),
            .I(N__12073));
    CascadeMux I__1755 (
            .O(N__12076),
            .I(N__12070));
    CascadeBuf I__1754 (
            .O(N__12073),
            .I(N__12067));
    CascadeBuf I__1753 (
            .O(N__12070),
            .I(N__12064));
    CascadeMux I__1752 (
            .O(N__12067),
            .I(N__12061));
    CascadeMux I__1751 (
            .O(N__12064),
            .I(N__12058));
    CascadeBuf I__1750 (
            .O(N__12061),
            .I(N__12055));
    CascadeBuf I__1749 (
            .O(N__12058),
            .I(N__12052));
    CascadeMux I__1748 (
            .O(N__12055),
            .I(N__12049));
    CascadeMux I__1747 (
            .O(N__12052),
            .I(N__12046));
    CascadeBuf I__1746 (
            .O(N__12049),
            .I(N__12043));
    CascadeBuf I__1745 (
            .O(N__12046),
            .I(N__12040));
    CascadeMux I__1744 (
            .O(N__12043),
            .I(N__12037));
    CascadeMux I__1743 (
            .O(N__12040),
            .I(N__12034));
    CascadeBuf I__1742 (
            .O(N__12037),
            .I(N__12031));
    CascadeBuf I__1741 (
            .O(N__12034),
            .I(N__12028));
    CascadeMux I__1740 (
            .O(N__12031),
            .I(N__12025));
    CascadeMux I__1739 (
            .O(N__12028),
            .I(N__12022));
    CascadeBuf I__1738 (
            .O(N__12025),
            .I(N__12019));
    CascadeBuf I__1737 (
            .O(N__12022),
            .I(N__12016));
    CascadeMux I__1736 (
            .O(N__12019),
            .I(N__12013));
    CascadeMux I__1735 (
            .O(N__12016),
            .I(N__12010));
    CascadeBuf I__1734 (
            .O(N__12013),
            .I(N__12007));
    CascadeBuf I__1733 (
            .O(N__12010),
            .I(N__12004));
    CascadeMux I__1732 (
            .O(N__12007),
            .I(N__12001));
    CascadeMux I__1731 (
            .O(N__12004),
            .I(N__11998));
    CascadeBuf I__1730 (
            .O(N__12001),
            .I(N__11995));
    CascadeBuf I__1729 (
            .O(N__11998),
            .I(N__11992));
    CascadeMux I__1728 (
            .O(N__11995),
            .I(N__11989));
    CascadeMux I__1727 (
            .O(N__11992),
            .I(N__11986));
    CascadeBuf I__1726 (
            .O(N__11989),
            .I(N__11983));
    CascadeBuf I__1725 (
            .O(N__11986),
            .I(N__11980));
    CascadeMux I__1724 (
            .O(N__11983),
            .I(N__11977));
    CascadeMux I__1723 (
            .O(N__11980),
            .I(N__11974));
    CascadeBuf I__1722 (
            .O(N__11977),
            .I(N__11971));
    CascadeBuf I__1721 (
            .O(N__11974),
            .I(N__11968));
    CascadeMux I__1720 (
            .O(N__11971),
            .I(N__11965));
    CascadeMux I__1719 (
            .O(N__11968),
            .I(N__11962));
    CascadeBuf I__1718 (
            .O(N__11965),
            .I(N__11959));
    CascadeBuf I__1717 (
            .O(N__11962),
            .I(N__11956));
    CascadeMux I__1716 (
            .O(N__11959),
            .I(N__11953));
    CascadeMux I__1715 (
            .O(N__11956),
            .I(N__11950));
    CascadeBuf I__1714 (
            .O(N__11953),
            .I(N__11947));
    CascadeBuf I__1713 (
            .O(N__11950),
            .I(N__11944));
    CascadeMux I__1712 (
            .O(N__11947),
            .I(N__11941));
    CascadeMux I__1711 (
            .O(N__11944),
            .I(N__11938));
    CascadeBuf I__1710 (
            .O(N__11941),
            .I(N__11935));
    CascadeBuf I__1709 (
            .O(N__11938),
            .I(N__11932));
    CascadeMux I__1708 (
            .O(N__11935),
            .I(N__11929));
    CascadeMux I__1707 (
            .O(N__11932),
            .I(N__11926));
    CascadeBuf I__1706 (
            .O(N__11929),
            .I(N__11923));
    CascadeBuf I__1705 (
            .O(N__11926),
            .I(N__11920));
    CascadeMux I__1704 (
            .O(N__11923),
            .I(N__11917));
    CascadeMux I__1703 (
            .O(N__11920),
            .I(N__11914));
    CascadeBuf I__1702 (
            .O(N__11917),
            .I(N__11911));
    InMux I__1701 (
            .O(N__11914),
            .I(N__11908));
    CascadeMux I__1700 (
            .O(N__11911),
            .I(N__11905));
    LocalMux I__1699 (
            .O(N__11908),
            .I(N__11902));
    InMux I__1698 (
            .O(N__11905),
            .I(N__11899));
    Span4Mux_v I__1697 (
            .O(N__11902),
            .I(N__11896));
    LocalMux I__1696 (
            .O(N__11899),
            .I(N__11893));
    Span4Mux_v I__1695 (
            .O(N__11896),
            .I(N__11890));
    Span12Mux_s9_v I__1694 (
            .O(N__11893),
            .I(N__11887));
    Span4Mux_v I__1693 (
            .O(N__11890),
            .I(N__11884));
    Span12Mux_h I__1692 (
            .O(N__11887),
            .I(N__11881));
    Span4Mux_h I__1691 (
            .O(N__11884),
            .I(N__11878));
    Odrv12 I__1690 (
            .O(N__11881),
            .I(n23));
    Odrv4 I__1689 (
            .O(N__11878),
            .I(n23));
    InMux I__1688 (
            .O(N__11873),
            .I(N__11869));
    InMux I__1687 (
            .O(N__11872),
            .I(N__11866));
    LocalMux I__1686 (
            .O(N__11869),
            .I(\transmit_module.video_signal_controller.n3366 ));
    LocalMux I__1685 (
            .O(N__11866),
            .I(\transmit_module.video_signal_controller.n3366 ));
    CascadeMux I__1684 (
            .O(N__11861),
            .I(N__11857));
    InMux I__1683 (
            .O(N__11860),
            .I(N__11853));
    InMux I__1682 (
            .O(N__11857),
            .I(N__11850));
    InMux I__1681 (
            .O(N__11856),
            .I(N__11847));
    LocalMux I__1680 (
            .O(N__11853),
            .I(N__11843));
    LocalMux I__1679 (
            .O(N__11850),
            .I(N__11840));
    LocalMux I__1678 (
            .O(N__11847),
            .I(N__11837));
    InMux I__1677 (
            .O(N__11846),
            .I(N__11834));
    Span4Mux_v I__1676 (
            .O(N__11843),
            .I(N__11829));
    Span4Mux_v I__1675 (
            .O(N__11840),
            .I(N__11829));
    Span4Mux_h I__1674 (
            .O(N__11837),
            .I(N__11826));
    LocalMux I__1673 (
            .O(N__11834),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    Odrv4 I__1672 (
            .O(N__11829),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    Odrv4 I__1671 (
            .O(N__11826),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    InMux I__1670 (
            .O(N__11819),
            .I(N__11815));
    InMux I__1669 (
            .O(N__11818),
            .I(N__11812));
    LocalMux I__1668 (
            .O(N__11815),
            .I(N__11809));
    LocalMux I__1667 (
            .O(N__11812),
            .I(\transmit_module.video_signal_controller.n2017 ));
    Odrv4 I__1666 (
            .O(N__11809),
            .I(\transmit_module.video_signal_controller.n2017 ));
    CascadeMux I__1665 (
            .O(N__11804),
            .I(\transmit_module.video_signal_controller.n3007_cascade_ ));
    InMux I__1664 (
            .O(N__11801),
            .I(N__11797));
    InMux I__1663 (
            .O(N__11800),
            .I(N__11794));
    LocalMux I__1662 (
            .O(N__11797),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_588 ));
    LocalMux I__1661 (
            .O(N__11794),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_588 ));
    InMux I__1660 (
            .O(N__11789),
            .I(N__11786));
    LocalMux I__1659 (
            .O(N__11786),
            .I(\transmit_module.n143 ));
    CascadeMux I__1658 (
            .O(N__11783),
            .I(\transmit_module.n143_cascade_ ));
    CascadeMux I__1657 (
            .O(N__11780),
            .I(N__11776));
    CascadeMux I__1656 (
            .O(N__11779),
            .I(N__11773));
    CascadeBuf I__1655 (
            .O(N__11776),
            .I(N__11770));
    CascadeBuf I__1654 (
            .O(N__11773),
            .I(N__11767));
    CascadeMux I__1653 (
            .O(N__11770),
            .I(N__11764));
    CascadeMux I__1652 (
            .O(N__11767),
            .I(N__11761));
    CascadeBuf I__1651 (
            .O(N__11764),
            .I(N__11758));
    CascadeBuf I__1650 (
            .O(N__11761),
            .I(N__11755));
    CascadeMux I__1649 (
            .O(N__11758),
            .I(N__11752));
    CascadeMux I__1648 (
            .O(N__11755),
            .I(N__11749));
    CascadeBuf I__1647 (
            .O(N__11752),
            .I(N__11746));
    CascadeBuf I__1646 (
            .O(N__11749),
            .I(N__11743));
    CascadeMux I__1645 (
            .O(N__11746),
            .I(N__11740));
    CascadeMux I__1644 (
            .O(N__11743),
            .I(N__11737));
    CascadeBuf I__1643 (
            .O(N__11740),
            .I(N__11734));
    CascadeBuf I__1642 (
            .O(N__11737),
            .I(N__11731));
    CascadeMux I__1641 (
            .O(N__11734),
            .I(N__11728));
    CascadeMux I__1640 (
            .O(N__11731),
            .I(N__11725));
    CascadeBuf I__1639 (
            .O(N__11728),
            .I(N__11722));
    CascadeBuf I__1638 (
            .O(N__11725),
            .I(N__11719));
    CascadeMux I__1637 (
            .O(N__11722),
            .I(N__11716));
    CascadeMux I__1636 (
            .O(N__11719),
            .I(N__11713));
    CascadeBuf I__1635 (
            .O(N__11716),
            .I(N__11710));
    CascadeBuf I__1634 (
            .O(N__11713),
            .I(N__11707));
    CascadeMux I__1633 (
            .O(N__11710),
            .I(N__11704));
    CascadeMux I__1632 (
            .O(N__11707),
            .I(N__11701));
    CascadeBuf I__1631 (
            .O(N__11704),
            .I(N__11698));
    CascadeBuf I__1630 (
            .O(N__11701),
            .I(N__11695));
    CascadeMux I__1629 (
            .O(N__11698),
            .I(N__11692));
    CascadeMux I__1628 (
            .O(N__11695),
            .I(N__11689));
    CascadeBuf I__1627 (
            .O(N__11692),
            .I(N__11686));
    CascadeBuf I__1626 (
            .O(N__11689),
            .I(N__11683));
    CascadeMux I__1625 (
            .O(N__11686),
            .I(N__11680));
    CascadeMux I__1624 (
            .O(N__11683),
            .I(N__11677));
    CascadeBuf I__1623 (
            .O(N__11680),
            .I(N__11674));
    CascadeBuf I__1622 (
            .O(N__11677),
            .I(N__11671));
    CascadeMux I__1621 (
            .O(N__11674),
            .I(N__11668));
    CascadeMux I__1620 (
            .O(N__11671),
            .I(N__11665));
    CascadeBuf I__1619 (
            .O(N__11668),
            .I(N__11662));
    CascadeBuf I__1618 (
            .O(N__11665),
            .I(N__11659));
    CascadeMux I__1617 (
            .O(N__11662),
            .I(N__11656));
    CascadeMux I__1616 (
            .O(N__11659),
            .I(N__11653));
    CascadeBuf I__1615 (
            .O(N__11656),
            .I(N__11650));
    CascadeBuf I__1614 (
            .O(N__11653),
            .I(N__11647));
    CascadeMux I__1613 (
            .O(N__11650),
            .I(N__11644));
    CascadeMux I__1612 (
            .O(N__11647),
            .I(N__11641));
    CascadeBuf I__1611 (
            .O(N__11644),
            .I(N__11638));
    CascadeBuf I__1610 (
            .O(N__11641),
            .I(N__11635));
    CascadeMux I__1609 (
            .O(N__11638),
            .I(N__11632));
    CascadeMux I__1608 (
            .O(N__11635),
            .I(N__11629));
    CascadeBuf I__1607 (
            .O(N__11632),
            .I(N__11626));
    CascadeBuf I__1606 (
            .O(N__11629),
            .I(N__11623));
    CascadeMux I__1605 (
            .O(N__11626),
            .I(N__11620));
    CascadeMux I__1604 (
            .O(N__11623),
            .I(N__11617));
    CascadeBuf I__1603 (
            .O(N__11620),
            .I(N__11614));
    CascadeBuf I__1602 (
            .O(N__11617),
            .I(N__11611));
    CascadeMux I__1601 (
            .O(N__11614),
            .I(N__11608));
    CascadeMux I__1600 (
            .O(N__11611),
            .I(N__11605));
    CascadeBuf I__1599 (
            .O(N__11608),
            .I(N__11602));
    CascadeBuf I__1598 (
            .O(N__11605),
            .I(N__11599));
    CascadeMux I__1597 (
            .O(N__11602),
            .I(N__11596));
    CascadeMux I__1596 (
            .O(N__11599),
            .I(N__11593));
    InMux I__1595 (
            .O(N__11596),
            .I(N__11590));
    InMux I__1594 (
            .O(N__11593),
            .I(N__11587));
    LocalMux I__1593 (
            .O(N__11590),
            .I(N__11584));
    LocalMux I__1592 (
            .O(N__11587),
            .I(N__11581));
    Span4Mux_v I__1591 (
            .O(N__11584),
            .I(N__11578));
    Span4Mux_v I__1590 (
            .O(N__11581),
            .I(N__11575));
    Span4Mux_v I__1589 (
            .O(N__11578),
            .I(N__11572));
    Sp12to4 I__1588 (
            .O(N__11575),
            .I(N__11569));
    Span4Mux_v I__1587 (
            .O(N__11572),
            .I(N__11566));
    Span12Mux_v I__1586 (
            .O(N__11569),
            .I(N__11563));
    Span4Mux_h I__1585 (
            .O(N__11566),
            .I(N__11560));
    Odrv12 I__1584 (
            .O(N__11563),
            .I(n24));
    Odrv4 I__1583 (
            .O(N__11560),
            .I(n24));
    InMux I__1582 (
            .O(N__11555),
            .I(N__11549));
    InMux I__1581 (
            .O(N__11554),
            .I(N__11549));
    LocalMux I__1580 (
            .O(N__11549),
            .I(N__11545));
    InMux I__1579 (
            .O(N__11548),
            .I(N__11540));
    Span4Mux_h I__1578 (
            .O(N__11545),
            .I(N__11537));
    InMux I__1577 (
            .O(N__11544),
            .I(N__11534));
    InMux I__1576 (
            .O(N__11543),
            .I(N__11531));
    LocalMux I__1575 (
            .O(N__11540),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    Odrv4 I__1574 (
            .O(N__11537),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__1573 (
            .O(N__11534),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__1572 (
            .O(N__11531),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    InMux I__1571 (
            .O(N__11522),
            .I(N__11519));
    LocalMux I__1570 (
            .O(N__11519),
            .I(\transmit_module.video_signal_controller.n3007 ));
    CascadeMux I__1569 (
            .O(N__11516),
            .I(\transmit_module.n141_cascade_ ));
    CascadeMux I__1568 (
            .O(N__11513),
            .I(N__11510));
    CascadeBuf I__1567 (
            .O(N__11510),
            .I(N__11507));
    CascadeMux I__1566 (
            .O(N__11507),
            .I(N__11504));
    CascadeBuf I__1565 (
            .O(N__11504),
            .I(N__11500));
    CascadeMux I__1564 (
            .O(N__11503),
            .I(N__11497));
    CascadeMux I__1563 (
            .O(N__11500),
            .I(N__11494));
    CascadeBuf I__1562 (
            .O(N__11497),
            .I(N__11491));
    CascadeBuf I__1561 (
            .O(N__11494),
            .I(N__11488));
    CascadeMux I__1560 (
            .O(N__11491),
            .I(N__11485));
    CascadeMux I__1559 (
            .O(N__11488),
            .I(N__11482));
    CascadeBuf I__1558 (
            .O(N__11485),
            .I(N__11479));
    CascadeBuf I__1557 (
            .O(N__11482),
            .I(N__11476));
    CascadeMux I__1556 (
            .O(N__11479),
            .I(N__11473));
    CascadeMux I__1555 (
            .O(N__11476),
            .I(N__11470));
    CascadeBuf I__1554 (
            .O(N__11473),
            .I(N__11467));
    CascadeBuf I__1553 (
            .O(N__11470),
            .I(N__11464));
    CascadeMux I__1552 (
            .O(N__11467),
            .I(N__11461));
    CascadeMux I__1551 (
            .O(N__11464),
            .I(N__11458));
    CascadeBuf I__1550 (
            .O(N__11461),
            .I(N__11455));
    CascadeBuf I__1549 (
            .O(N__11458),
            .I(N__11452));
    CascadeMux I__1548 (
            .O(N__11455),
            .I(N__11449));
    CascadeMux I__1547 (
            .O(N__11452),
            .I(N__11446));
    CascadeBuf I__1546 (
            .O(N__11449),
            .I(N__11443));
    CascadeBuf I__1545 (
            .O(N__11446),
            .I(N__11440));
    CascadeMux I__1544 (
            .O(N__11443),
            .I(N__11437));
    CascadeMux I__1543 (
            .O(N__11440),
            .I(N__11434));
    CascadeBuf I__1542 (
            .O(N__11437),
            .I(N__11431));
    CascadeBuf I__1541 (
            .O(N__11434),
            .I(N__11428));
    CascadeMux I__1540 (
            .O(N__11431),
            .I(N__11425));
    CascadeMux I__1539 (
            .O(N__11428),
            .I(N__11422));
    CascadeBuf I__1538 (
            .O(N__11425),
            .I(N__11419));
    CascadeBuf I__1537 (
            .O(N__11422),
            .I(N__11416));
    CascadeMux I__1536 (
            .O(N__11419),
            .I(N__11413));
    CascadeMux I__1535 (
            .O(N__11416),
            .I(N__11410));
    CascadeBuf I__1534 (
            .O(N__11413),
            .I(N__11407));
    CascadeBuf I__1533 (
            .O(N__11410),
            .I(N__11404));
    CascadeMux I__1532 (
            .O(N__11407),
            .I(N__11401));
    CascadeMux I__1531 (
            .O(N__11404),
            .I(N__11398));
    CascadeBuf I__1530 (
            .O(N__11401),
            .I(N__11395));
    CascadeBuf I__1529 (
            .O(N__11398),
            .I(N__11392));
    CascadeMux I__1528 (
            .O(N__11395),
            .I(N__11389));
    CascadeMux I__1527 (
            .O(N__11392),
            .I(N__11386));
    CascadeBuf I__1526 (
            .O(N__11389),
            .I(N__11383));
    CascadeBuf I__1525 (
            .O(N__11386),
            .I(N__11380));
    CascadeMux I__1524 (
            .O(N__11383),
            .I(N__11377));
    CascadeMux I__1523 (
            .O(N__11380),
            .I(N__11374));
    CascadeBuf I__1522 (
            .O(N__11377),
            .I(N__11371));
    CascadeBuf I__1521 (
            .O(N__11374),
            .I(N__11368));
    CascadeMux I__1520 (
            .O(N__11371),
            .I(N__11365));
    CascadeMux I__1519 (
            .O(N__11368),
            .I(N__11362));
    CascadeBuf I__1518 (
            .O(N__11365),
            .I(N__11359));
    CascadeBuf I__1517 (
            .O(N__11362),
            .I(N__11356));
    CascadeMux I__1516 (
            .O(N__11359),
            .I(N__11353));
    CascadeMux I__1515 (
            .O(N__11356),
            .I(N__11350));
    CascadeBuf I__1514 (
            .O(N__11353),
            .I(N__11347));
    CascadeBuf I__1513 (
            .O(N__11350),
            .I(N__11344));
    CascadeMux I__1512 (
            .O(N__11347),
            .I(N__11341));
    CascadeMux I__1511 (
            .O(N__11344),
            .I(N__11338));
    CascadeBuf I__1510 (
            .O(N__11341),
            .I(N__11335));
    InMux I__1509 (
            .O(N__11338),
            .I(N__11332));
    CascadeMux I__1508 (
            .O(N__11335),
            .I(N__11329));
    LocalMux I__1507 (
            .O(N__11332),
            .I(N__11326));
    CascadeBuf I__1506 (
            .O(N__11329),
            .I(N__11323));
    Span4Mux_v I__1505 (
            .O(N__11326),
            .I(N__11320));
    CascadeMux I__1504 (
            .O(N__11323),
            .I(N__11317));
    Span4Mux_v I__1503 (
            .O(N__11320),
            .I(N__11314));
    InMux I__1502 (
            .O(N__11317),
            .I(N__11311));
    Span4Mux_h I__1501 (
            .O(N__11314),
            .I(N__11308));
    LocalMux I__1500 (
            .O(N__11311),
            .I(N__11305));
    Span4Mux_h I__1499 (
            .O(N__11308),
            .I(N__11302));
    Span4Mux_v I__1498 (
            .O(N__11305),
            .I(N__11299));
    Span4Mux_h I__1497 (
            .O(N__11302),
            .I(N__11296));
    Span4Mux_h I__1496 (
            .O(N__11299),
            .I(N__11293));
    Sp12to4 I__1495 (
            .O(N__11296),
            .I(N__11288));
    Sp12to4 I__1494 (
            .O(N__11293),
            .I(N__11288));
    Odrv12 I__1493 (
            .O(N__11288),
            .I(n22));
    InMux I__1492 (
            .O(N__11285),
            .I(N__11278));
    InMux I__1491 (
            .O(N__11284),
            .I(N__11278));
    CascadeMux I__1490 (
            .O(N__11283),
            .I(N__11275));
    LocalMux I__1489 (
            .O(N__11278),
            .I(N__11271));
    InMux I__1488 (
            .O(N__11275),
            .I(N__11266));
    InMux I__1487 (
            .O(N__11274),
            .I(N__11266));
    Odrv4 I__1486 (
            .O(N__11271),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    LocalMux I__1485 (
            .O(N__11266),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    InMux I__1484 (
            .O(N__11261),
            .I(N__11258));
    LocalMux I__1483 (
            .O(N__11258),
            .I(\transmit_module.n140 ));
    CascadeMux I__1482 (
            .O(N__11255),
            .I(\transmit_module.n140_cascade_ ));
    InMux I__1481 (
            .O(N__11252),
            .I(N__11246));
    InMux I__1480 (
            .O(N__11251),
            .I(N__11246));
    LocalMux I__1479 (
            .O(N__11246),
            .I(\transmit_module.n109 ));
    CascadeMux I__1478 (
            .O(N__11243),
            .I(N__11240));
    CascadeBuf I__1477 (
            .O(N__11240),
            .I(N__11236));
    CascadeMux I__1476 (
            .O(N__11239),
            .I(N__11233));
    CascadeMux I__1475 (
            .O(N__11236),
            .I(N__11230));
    CascadeBuf I__1474 (
            .O(N__11233),
            .I(N__11227));
    CascadeBuf I__1473 (
            .O(N__11230),
            .I(N__11224));
    CascadeMux I__1472 (
            .O(N__11227),
            .I(N__11221));
    CascadeMux I__1471 (
            .O(N__11224),
            .I(N__11218));
    CascadeBuf I__1470 (
            .O(N__11221),
            .I(N__11215));
    CascadeBuf I__1469 (
            .O(N__11218),
            .I(N__11212));
    CascadeMux I__1468 (
            .O(N__11215),
            .I(N__11209));
    CascadeMux I__1467 (
            .O(N__11212),
            .I(N__11206));
    CascadeBuf I__1466 (
            .O(N__11209),
            .I(N__11203));
    CascadeBuf I__1465 (
            .O(N__11206),
            .I(N__11200));
    CascadeMux I__1464 (
            .O(N__11203),
            .I(N__11197));
    CascadeMux I__1463 (
            .O(N__11200),
            .I(N__11194));
    CascadeBuf I__1462 (
            .O(N__11197),
            .I(N__11191));
    CascadeBuf I__1461 (
            .O(N__11194),
            .I(N__11188));
    CascadeMux I__1460 (
            .O(N__11191),
            .I(N__11185));
    CascadeMux I__1459 (
            .O(N__11188),
            .I(N__11182));
    CascadeBuf I__1458 (
            .O(N__11185),
            .I(N__11179));
    CascadeBuf I__1457 (
            .O(N__11182),
            .I(N__11176));
    CascadeMux I__1456 (
            .O(N__11179),
            .I(N__11173));
    CascadeMux I__1455 (
            .O(N__11176),
            .I(N__11170));
    CascadeBuf I__1454 (
            .O(N__11173),
            .I(N__11167));
    CascadeBuf I__1453 (
            .O(N__11170),
            .I(N__11164));
    CascadeMux I__1452 (
            .O(N__11167),
            .I(N__11161));
    CascadeMux I__1451 (
            .O(N__11164),
            .I(N__11158));
    CascadeBuf I__1450 (
            .O(N__11161),
            .I(N__11155));
    CascadeBuf I__1449 (
            .O(N__11158),
            .I(N__11152));
    CascadeMux I__1448 (
            .O(N__11155),
            .I(N__11149));
    CascadeMux I__1447 (
            .O(N__11152),
            .I(N__11146));
    CascadeBuf I__1446 (
            .O(N__11149),
            .I(N__11143));
    CascadeBuf I__1445 (
            .O(N__11146),
            .I(N__11140));
    CascadeMux I__1444 (
            .O(N__11143),
            .I(N__11137));
    CascadeMux I__1443 (
            .O(N__11140),
            .I(N__11134));
    CascadeBuf I__1442 (
            .O(N__11137),
            .I(N__11131));
    CascadeBuf I__1441 (
            .O(N__11134),
            .I(N__11128));
    CascadeMux I__1440 (
            .O(N__11131),
            .I(N__11125));
    CascadeMux I__1439 (
            .O(N__11128),
            .I(N__11122));
    CascadeBuf I__1438 (
            .O(N__11125),
            .I(N__11119));
    CascadeBuf I__1437 (
            .O(N__11122),
            .I(N__11116));
    CascadeMux I__1436 (
            .O(N__11119),
            .I(N__11113));
    CascadeMux I__1435 (
            .O(N__11116),
            .I(N__11110));
    CascadeBuf I__1434 (
            .O(N__11113),
            .I(N__11107));
    CascadeBuf I__1433 (
            .O(N__11110),
            .I(N__11104));
    CascadeMux I__1432 (
            .O(N__11107),
            .I(N__11101));
    CascadeMux I__1431 (
            .O(N__11104),
            .I(N__11098));
    CascadeBuf I__1430 (
            .O(N__11101),
            .I(N__11095));
    CascadeBuf I__1429 (
            .O(N__11098),
            .I(N__11092));
    CascadeMux I__1428 (
            .O(N__11095),
            .I(N__11089));
    CascadeMux I__1427 (
            .O(N__11092),
            .I(N__11086));
    CascadeBuf I__1426 (
            .O(N__11089),
            .I(N__11083));
    CascadeBuf I__1425 (
            .O(N__11086),
            .I(N__11080));
    CascadeMux I__1424 (
            .O(N__11083),
            .I(N__11077));
    CascadeMux I__1423 (
            .O(N__11080),
            .I(N__11074));
    CascadeBuf I__1422 (
            .O(N__11077),
            .I(N__11071));
    CascadeBuf I__1421 (
            .O(N__11074),
            .I(N__11068));
    CascadeMux I__1420 (
            .O(N__11071),
            .I(N__11065));
    CascadeMux I__1419 (
            .O(N__11068),
            .I(N__11062));
    CascadeBuf I__1418 (
            .O(N__11065),
            .I(N__11059));
    InMux I__1417 (
            .O(N__11062),
            .I(N__11056));
    CascadeMux I__1416 (
            .O(N__11059),
            .I(N__11053));
    LocalMux I__1415 (
            .O(N__11056),
            .I(N__11050));
    InMux I__1414 (
            .O(N__11053),
            .I(N__11047));
    Span4Mux_s2_v I__1413 (
            .O(N__11050),
            .I(N__11044));
    LocalMux I__1412 (
            .O(N__11047),
            .I(N__11041));
    Span4Mux_v I__1411 (
            .O(N__11044),
            .I(N__11038));
    Sp12to4 I__1410 (
            .O(N__11041),
            .I(N__11035));
    Span4Mux_v I__1409 (
            .O(N__11038),
            .I(N__11032));
    Span12Mux_s11_v I__1408 (
            .O(N__11035),
            .I(N__11029));
    Span4Mux_v I__1407 (
            .O(N__11032),
            .I(N__11026));
    Span12Mux_h I__1406 (
            .O(N__11029),
            .I(N__11023));
    Span4Mux_h I__1405 (
            .O(N__11026),
            .I(N__11020));
    Odrv12 I__1404 (
            .O(N__11023),
            .I(n21));
    Odrv4 I__1403 (
            .O(N__11020),
            .I(n21));
    InMux I__1402 (
            .O(N__11015),
            .I(N__11010));
    InMux I__1401 (
            .O(N__11014),
            .I(N__11006));
    InMux I__1400 (
            .O(N__11013),
            .I(N__11003));
    LocalMux I__1399 (
            .O(N__11010),
            .I(N__11000));
    InMux I__1398 (
            .O(N__11009),
            .I(N__10997));
    LocalMux I__1397 (
            .O(N__11006),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1396 (
            .O(N__11003),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    Odrv4 I__1395 (
            .O(N__11000),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1394 (
            .O(N__10997),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    InMux I__1393 (
            .O(N__10988),
            .I(N__10985));
    LocalMux I__1392 (
            .O(N__10985),
            .I(N__10982));
    Odrv4 I__1391 (
            .O(N__10982),
            .I(\transmit_module.video_signal_controller.n3520 ));
    CascadeMux I__1390 (
            .O(N__10979),
            .I(N__10976));
    InMux I__1389 (
            .O(N__10976),
            .I(N__10972));
    InMux I__1388 (
            .O(N__10975),
            .I(N__10969));
    LocalMux I__1387 (
            .O(N__10972),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    LocalMux I__1386 (
            .O(N__10969),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    InMux I__1385 (
            .O(N__10964),
            .I(N__10959));
    InMux I__1384 (
            .O(N__10963),
            .I(N__10955));
    InMux I__1383 (
            .O(N__10962),
            .I(N__10952));
    LocalMux I__1382 (
            .O(N__10959),
            .I(N__10949));
    InMux I__1381 (
            .O(N__10958),
            .I(N__10946));
    LocalMux I__1380 (
            .O(N__10955),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1379 (
            .O(N__10952),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    Odrv4 I__1378 (
            .O(N__10949),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1377 (
            .O(N__10946),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    CascadeMux I__1376 (
            .O(N__10937),
            .I(N__10934));
    InMux I__1375 (
            .O(N__10934),
            .I(N__10931));
    LocalMux I__1374 (
            .O(N__10931),
            .I(N__10928));
    Odrv4 I__1373 (
            .O(N__10928),
            .I(\transmit_module.video_signal_controller.n2958 ));
    CascadeMux I__1372 (
            .O(N__10925),
            .I(N__10922));
    InMux I__1371 (
            .O(N__10922),
            .I(N__10919));
    LocalMux I__1370 (
            .O(N__10919),
            .I(N__10916));
    Span4Mux_h I__1369 (
            .O(N__10916),
            .I(N__10913));
    Odrv4 I__1368 (
            .O(N__10913),
            .I(\transmit_module.video_signal_controller.n2975 ));
    InMux I__1367 (
            .O(N__10910),
            .I(N__10907));
    LocalMux I__1366 (
            .O(N__10907),
            .I(\receive_module.rx_counter.n10 ));
    CascadeMux I__1365 (
            .O(N__10904),
            .I(\receive_module.rx_counter.n14_cascade_ ));
    InMux I__1364 (
            .O(N__10901),
            .I(N__10898));
    LocalMux I__1363 (
            .O(N__10898),
            .I(N__10895));
    Span4Mux_v I__1362 (
            .O(N__10895),
            .I(N__10892));
    Span4Mux_h I__1361 (
            .O(N__10892),
            .I(N__10889));
    Odrv4 I__1360 (
            .O(N__10889),
            .I(\line_buffer.n539 ));
    InMux I__1359 (
            .O(N__10886),
            .I(N__10883));
    LocalMux I__1358 (
            .O(N__10883),
            .I(N__10880));
    Span12Mux_v I__1357 (
            .O(N__10880),
            .I(N__10877));
    Span12Mux_h I__1356 (
            .O(N__10877),
            .I(N__10874));
    Odrv12 I__1355 (
            .O(N__10874),
            .I(\line_buffer.n531 ));
    InMux I__1354 (
            .O(N__10871),
            .I(N__10865));
    InMux I__1353 (
            .O(N__10870),
            .I(N__10865));
    LocalMux I__1352 (
            .O(N__10865),
            .I(N__10862));
    Span4Mux_h I__1351 (
            .O(N__10862),
            .I(N__10857));
    InMux I__1350 (
            .O(N__10861),
            .I(N__10852));
    InMux I__1349 (
            .O(N__10860),
            .I(N__10852));
    Odrv4 I__1348 (
            .O(N__10857),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__1347 (
            .O(N__10852),
            .I(\transmit_module.old_VGA_HS ));
    InMux I__1346 (
            .O(N__10847),
            .I(N__10844));
    LocalMux I__1345 (
            .O(N__10844),
            .I(N__10841));
    Odrv4 I__1344 (
            .O(N__10841),
            .I(\transmit_module.ADDR_Y_COMPONENT_7 ));
    InMux I__1343 (
            .O(N__10838),
            .I(N__10835));
    LocalMux I__1342 (
            .O(N__10835),
            .I(N__10832));
    Odrv4 I__1341 (
            .O(N__10832),
            .I(\transmit_module.video_signal_controller.n7 ));
    IoInMux I__1340 (
            .O(N__10829),
            .I(N__10826));
    LocalMux I__1339 (
            .O(N__10826),
            .I(N__10823));
    IoSpan4Mux I__1338 (
            .O(N__10823),
            .I(N__10820));
    Sp12to4 I__1337 (
            .O(N__10820),
            .I(N__10815));
    InMux I__1336 (
            .O(N__10819),
            .I(N__10810));
    InMux I__1335 (
            .O(N__10818),
            .I(N__10810));
    Span12Mux_h I__1334 (
            .O(N__10815),
            .I(N__10804));
    LocalMux I__1333 (
            .O(N__10810),
            .I(N__10801));
    InMux I__1332 (
            .O(N__10809),
            .I(N__10794));
    InMux I__1331 (
            .O(N__10808),
            .I(N__10794));
    InMux I__1330 (
            .O(N__10807),
            .I(N__10794));
    Odrv12 I__1329 (
            .O(N__10804),
            .I(ADV_HSYNC_c));
    Odrv4 I__1328 (
            .O(N__10801),
            .I(ADV_HSYNC_c));
    LocalMux I__1327 (
            .O(N__10794),
            .I(ADV_HSYNC_c));
    InMux I__1326 (
            .O(N__10787),
            .I(\receive_module.rx_counter.n3175 ));
    InMux I__1325 (
            .O(N__10784),
            .I(\receive_module.rx_counter.n3176 ));
    InMux I__1324 (
            .O(N__10781),
            .I(\receive_module.rx_counter.n3177 ));
    InMux I__1323 (
            .O(N__10778),
            .I(\receive_module.rx_counter.n3178 ));
    InMux I__1322 (
            .O(N__10775),
            .I(\receive_module.rx_counter.n3179 ));
    InMux I__1321 (
            .O(N__10772),
            .I(\receive_module.rx_counter.n3180 ));
    InMux I__1320 (
            .O(N__10769),
            .I(\receive_module.rx_counter.n3181 ));
    InMux I__1319 (
            .O(N__10766),
            .I(bfn_13_12_0_));
    InMux I__1318 (
            .O(N__10763),
            .I(\receive_module.rx_counter.n3211 ));
    InMux I__1317 (
            .O(N__10760),
            .I(\receive_module.rx_counter.n3212 ));
    InMux I__1316 (
            .O(N__10757),
            .I(\receive_module.rx_counter.n3213 ));
    InMux I__1315 (
            .O(N__10754),
            .I(\receive_module.rx_counter.n3214 ));
    InMux I__1314 (
            .O(N__10751),
            .I(\receive_module.rx_counter.n3215 ));
    InMux I__1313 (
            .O(N__10748),
            .I(\receive_module.rx_counter.n3216 ));
    InMux I__1312 (
            .O(N__10745),
            .I(bfn_13_10_0_));
    InMux I__1311 (
            .O(N__10742),
            .I(\receive_module.rx_counter.n3218 ));
    InMux I__1310 (
            .O(N__10739),
            .I(bfn_13_11_0_));
    InMux I__1309 (
            .O(N__10736),
            .I(N__10732));
    InMux I__1308 (
            .O(N__10735),
            .I(N__10729));
    LocalMux I__1307 (
            .O(N__10732),
            .I(N__10725));
    LocalMux I__1306 (
            .O(N__10729),
            .I(N__10721));
    InMux I__1305 (
            .O(N__10728),
            .I(N__10718));
    Span4Mux_v I__1304 (
            .O(N__10725),
            .I(N__10712));
    InMux I__1303 (
            .O(N__10724),
            .I(N__10709));
    Sp12to4 I__1302 (
            .O(N__10721),
            .I(N__10703));
    LocalMux I__1301 (
            .O(N__10718),
            .I(N__10703));
    InMux I__1300 (
            .O(N__10717),
            .I(N__10700));
    InMux I__1299 (
            .O(N__10716),
            .I(N__10697));
    InMux I__1298 (
            .O(N__10715),
            .I(N__10694));
    Span4Mux_v I__1297 (
            .O(N__10712),
            .I(N__10689));
    LocalMux I__1296 (
            .O(N__10709),
            .I(N__10689));
    InMux I__1295 (
            .O(N__10708),
            .I(N__10686));
    Span12Mux_s9_v I__1294 (
            .O(N__10703),
            .I(N__10679));
    LocalMux I__1293 (
            .O(N__10700),
            .I(N__10679));
    LocalMux I__1292 (
            .O(N__10697),
            .I(N__10679));
    LocalMux I__1291 (
            .O(N__10694),
            .I(N__10676));
    Span4Mux_v I__1290 (
            .O(N__10689),
            .I(N__10673));
    LocalMux I__1289 (
            .O(N__10686),
            .I(N__10670));
    Span12Mux_v I__1288 (
            .O(N__10679),
            .I(N__10665));
    Span12Mux_s10_v I__1287 (
            .O(N__10676),
            .I(N__10665));
    Span4Mux_v I__1286 (
            .O(N__10673),
            .I(N__10660));
    Span4Mux_h I__1285 (
            .O(N__10670),
            .I(N__10660));
    Span12Mux_h I__1284 (
            .O(N__10665),
            .I(N__10657));
    Span4Mux_h I__1283 (
            .O(N__10660),
            .I(N__10654));
    Odrv12 I__1282 (
            .O(N__10657),
            .I(RX_DATA_0));
    Odrv4 I__1281 (
            .O(N__10654),
            .I(RX_DATA_0));
    InMux I__1280 (
            .O(N__10649),
            .I(N__10646));
    LocalMux I__1279 (
            .O(N__10646),
            .I(N__10643));
    Span4Mux_h I__1278 (
            .O(N__10643),
            .I(N__10640));
    Span4Mux_v I__1277 (
            .O(N__10640),
            .I(N__10637));
    Odrv4 I__1276 (
            .O(N__10637),
            .I(TVP_VIDEO_c_4));
    InMux I__1275 (
            .O(N__10634),
            .I(N__10631));
    LocalMux I__1274 (
            .O(N__10631),
            .I(\tvp_video_buffer.BUFFER_0_4 ));
    InMux I__1273 (
            .O(N__10628),
            .I(N__10625));
    LocalMux I__1272 (
            .O(N__10625),
            .I(N__10622));
    Span12Mux_h I__1271 (
            .O(N__10622),
            .I(N__10619));
    Odrv12 I__1270 (
            .O(N__10619),
            .I(TVP_VIDEO_c_8));
    InMux I__1269 (
            .O(N__10616),
            .I(N__10613));
    LocalMux I__1268 (
            .O(N__10613),
            .I(\tvp_video_buffer.BUFFER_1_3 ));
    InMux I__1267 (
            .O(N__10610),
            .I(N__10606));
    InMux I__1266 (
            .O(N__10609),
            .I(N__10603));
    LocalMux I__1265 (
            .O(N__10606),
            .I(N__10596));
    LocalMux I__1264 (
            .O(N__10603),
            .I(N__10591));
    InMux I__1263 (
            .O(N__10602),
            .I(N__10588));
    InMux I__1262 (
            .O(N__10601),
            .I(N__10585));
    InMux I__1261 (
            .O(N__10600),
            .I(N__10582));
    InMux I__1260 (
            .O(N__10599),
            .I(N__10579));
    Span4Mux_v I__1259 (
            .O(N__10596),
            .I(N__10576));
    InMux I__1258 (
            .O(N__10595),
            .I(N__10573));
    InMux I__1257 (
            .O(N__10594),
            .I(N__10570));
    Sp12to4 I__1256 (
            .O(N__10591),
            .I(N__10565));
    LocalMux I__1255 (
            .O(N__10588),
            .I(N__10565));
    LocalMux I__1254 (
            .O(N__10585),
            .I(N__10560));
    LocalMux I__1253 (
            .O(N__10582),
            .I(N__10560));
    LocalMux I__1252 (
            .O(N__10579),
            .I(N__10557));
    Span4Mux_v I__1251 (
            .O(N__10576),
            .I(N__10552));
    LocalMux I__1250 (
            .O(N__10573),
            .I(N__10552));
    LocalMux I__1249 (
            .O(N__10570),
            .I(N__10549));
    Span12Mux_v I__1248 (
            .O(N__10565),
            .I(N__10546));
    Span12Mux_v I__1247 (
            .O(N__10560),
            .I(N__10541));
    Span12Mux_s5_v I__1246 (
            .O(N__10557),
            .I(N__10541));
    Span4Mux_v I__1245 (
            .O(N__10552),
            .I(N__10536));
    Span4Mux_v I__1244 (
            .O(N__10549),
            .I(N__10536));
    Span12Mux_h I__1243 (
            .O(N__10546),
            .I(N__10531));
    Span12Mux_h I__1242 (
            .O(N__10541),
            .I(N__10531));
    Span4Mux_h I__1241 (
            .O(N__10536),
            .I(N__10528));
    Odrv12 I__1240 (
            .O(N__10531),
            .I(RX_DATA_1));
    Odrv4 I__1239 (
            .O(N__10528),
            .I(RX_DATA_1));
    InMux I__1238 (
            .O(N__10523),
            .I(N__10520));
    LocalMux I__1237 (
            .O(N__10520),
            .I(\tvp_video_buffer.BUFFER_1_4 ));
    InMux I__1236 (
            .O(N__10517),
            .I(N__10514));
    LocalMux I__1235 (
            .O(N__10514),
            .I(N__10510));
    InMux I__1234 (
            .O(N__10513),
            .I(N__10507));
    Span4Mux_s2_v I__1233 (
            .O(N__10510),
            .I(N__10504));
    LocalMux I__1232 (
            .O(N__10507),
            .I(N__10501));
    Span4Mux_v I__1231 (
            .O(N__10504),
            .I(N__10497));
    Span4Mux_v I__1230 (
            .O(N__10501),
            .I(N__10493));
    InMux I__1229 (
            .O(N__10500),
            .I(N__10490));
    Span4Mux_v I__1228 (
            .O(N__10497),
            .I(N__10486));
    InMux I__1227 (
            .O(N__10496),
            .I(N__10483));
    Span4Mux_v I__1226 (
            .O(N__10493),
            .I(N__10477));
    LocalMux I__1225 (
            .O(N__10490),
            .I(N__10477));
    InMux I__1224 (
            .O(N__10489),
            .I(N__10472));
    Span4Mux_v I__1223 (
            .O(N__10486),
            .I(N__10467));
    LocalMux I__1222 (
            .O(N__10483),
            .I(N__10467));
    InMux I__1221 (
            .O(N__10482),
            .I(N__10464));
    Span4Mux_v I__1220 (
            .O(N__10477),
            .I(N__10461));
    InMux I__1219 (
            .O(N__10476),
            .I(N__10458));
    InMux I__1218 (
            .O(N__10475),
            .I(N__10455));
    LocalMux I__1217 (
            .O(N__10472),
            .I(N__10452));
    Span4Mux_v I__1216 (
            .O(N__10467),
            .I(N__10449));
    LocalMux I__1215 (
            .O(N__10464),
            .I(N__10446));
    Sp12to4 I__1214 (
            .O(N__10461),
            .I(N__10439));
    LocalMux I__1213 (
            .O(N__10458),
            .I(N__10439));
    LocalMux I__1212 (
            .O(N__10455),
            .I(N__10439));
    Span4Mux_v I__1211 (
            .O(N__10452),
            .I(N__10436));
    Span4Mux_v I__1210 (
            .O(N__10449),
            .I(N__10431));
    Span4Mux_h I__1209 (
            .O(N__10446),
            .I(N__10431));
    Span12Mux_v I__1208 (
            .O(N__10439),
            .I(N__10428));
    Span4Mux_h I__1207 (
            .O(N__10436),
            .I(N__10423));
    Span4Mux_h I__1206 (
            .O(N__10431),
            .I(N__10423));
    Odrv12 I__1205 (
            .O(N__10428),
            .I(RX_DATA_2));
    Odrv4 I__1204 (
            .O(N__10423),
            .I(RX_DATA_2));
    InMux I__1203 (
            .O(N__10418),
            .I(N__10415));
    LocalMux I__1202 (
            .O(N__10415),
            .I(\tvp_video_buffer.BUFFER_0_8 ));
    InMux I__1201 (
            .O(N__10412),
            .I(N__10409));
    LocalMux I__1200 (
            .O(N__10409),
            .I(\tvp_video_buffer.BUFFER_1_8 ));
    InMux I__1199 (
            .O(N__10406),
            .I(bfn_13_9_0_));
    InMux I__1198 (
            .O(N__10403),
            .I(\receive_module.rx_counter.n3210 ));
    CascadeMux I__1197 (
            .O(N__10400),
            .I(N__10396));
    InMux I__1196 (
            .O(N__10399),
            .I(N__10391));
    InMux I__1195 (
            .O(N__10396),
            .I(N__10384));
    InMux I__1194 (
            .O(N__10395),
            .I(N__10384));
    InMux I__1193 (
            .O(N__10394),
            .I(N__10384));
    LocalMux I__1192 (
            .O(N__10391),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__1191 (
            .O(N__10384),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    InMux I__1190 (
            .O(N__10379),
            .I(N__10373));
    InMux I__1189 (
            .O(N__10378),
            .I(N__10366));
    InMux I__1188 (
            .O(N__10377),
            .I(N__10366));
    InMux I__1187 (
            .O(N__10376),
            .I(N__10366));
    LocalMux I__1186 (
            .O(N__10373),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__1185 (
            .O(N__10366),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    InMux I__1184 (
            .O(N__10361),
            .I(N__10358));
    LocalMux I__1183 (
            .O(N__10358),
            .I(N__10352));
    InMux I__1182 (
            .O(N__10357),
            .I(N__10349));
    InMux I__1181 (
            .O(N__10356),
            .I(N__10344));
    InMux I__1180 (
            .O(N__10355),
            .I(N__10344));
    Span4Mux_h I__1179 (
            .O(N__10352),
            .I(N__10341));
    LocalMux I__1178 (
            .O(N__10349),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1177 (
            .O(N__10344),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    Odrv4 I__1176 (
            .O(N__10341),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    CascadeMux I__1175 (
            .O(N__10334),
            .I(\transmit_module.video_signal_controller.n3482_cascade_ ));
    InMux I__1174 (
            .O(N__10331),
            .I(N__10328));
    LocalMux I__1173 (
            .O(N__10328),
            .I(N__10322));
    InMux I__1172 (
            .O(N__10327),
            .I(N__10319));
    InMux I__1171 (
            .O(N__10326),
            .I(N__10314));
    InMux I__1170 (
            .O(N__10325),
            .I(N__10314));
    Span4Mux_h I__1169 (
            .O(N__10322),
            .I(N__10311));
    LocalMux I__1168 (
            .O(N__10319),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__1167 (
            .O(N__10314),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    Odrv4 I__1166 (
            .O(N__10311),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    InMux I__1165 (
            .O(N__10304),
            .I(N__10301));
    LocalMux I__1164 (
            .O(N__10301),
            .I(\transmit_module.video_signal_controller.n55 ));
    CascadeMux I__1163 (
            .O(N__10298),
            .I(\transmit_module.video_signal_controller.n3478_cascade_ ));
    InMux I__1162 (
            .O(N__10295),
            .I(N__10290));
    InMux I__1161 (
            .O(N__10294),
            .I(N__10287));
    InMux I__1160 (
            .O(N__10293),
            .I(N__10284));
    LocalMux I__1159 (
            .O(N__10290),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1158 (
            .O(N__10287),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1157 (
            .O(N__10284),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    CascadeMux I__1156 (
            .O(N__10277),
            .I(N__10272));
    InMux I__1155 (
            .O(N__10276),
            .I(N__10269));
    InMux I__1154 (
            .O(N__10275),
            .I(N__10264));
    InMux I__1153 (
            .O(N__10272),
            .I(N__10264));
    LocalMux I__1152 (
            .O(N__10269),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    LocalMux I__1151 (
            .O(N__10264),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    InMux I__1150 (
            .O(N__10259),
            .I(N__10256));
    LocalMux I__1149 (
            .O(N__10256),
            .I(N__10253));
    Span4Mux_h I__1148 (
            .O(N__10253),
            .I(N__10250));
    Odrv4 I__1147 (
            .O(N__10250),
            .I(\transmit_module.ADDR_Y_COMPONENT_13 ));
    CEMux I__1146 (
            .O(N__10247),
            .I(N__10243));
    CEMux I__1145 (
            .O(N__10246),
            .I(N__10240));
    LocalMux I__1144 (
            .O(N__10243),
            .I(N__10237));
    LocalMux I__1143 (
            .O(N__10240),
            .I(N__10234));
    Span4Mux_v I__1142 (
            .O(N__10237),
            .I(N__10231));
    Span4Mux_h I__1141 (
            .O(N__10234),
            .I(N__10228));
    Span4Mux_h I__1140 (
            .O(N__10231),
            .I(N__10225));
    Odrv4 I__1139 (
            .O(N__10228),
            .I(\transmit_module.n2073 ));
    Odrv4 I__1138 (
            .O(N__10225),
            .I(\transmit_module.n2073 ));
    CascadeMux I__1137 (
            .O(N__10220),
            .I(N__10216));
    CascadeMux I__1136 (
            .O(N__10219),
            .I(N__10213));
    CascadeBuf I__1135 (
            .O(N__10216),
            .I(N__10210));
    CascadeBuf I__1134 (
            .O(N__10213),
            .I(N__10207));
    CascadeMux I__1133 (
            .O(N__10210),
            .I(N__10204));
    CascadeMux I__1132 (
            .O(N__10207),
            .I(N__10201));
    CascadeBuf I__1131 (
            .O(N__10204),
            .I(N__10198));
    CascadeBuf I__1130 (
            .O(N__10201),
            .I(N__10195));
    CascadeMux I__1129 (
            .O(N__10198),
            .I(N__10192));
    CascadeMux I__1128 (
            .O(N__10195),
            .I(N__10189));
    CascadeBuf I__1127 (
            .O(N__10192),
            .I(N__10186));
    CascadeBuf I__1126 (
            .O(N__10189),
            .I(N__10183));
    CascadeMux I__1125 (
            .O(N__10186),
            .I(N__10180));
    CascadeMux I__1124 (
            .O(N__10183),
            .I(N__10177));
    CascadeBuf I__1123 (
            .O(N__10180),
            .I(N__10174));
    CascadeBuf I__1122 (
            .O(N__10177),
            .I(N__10171));
    CascadeMux I__1121 (
            .O(N__10174),
            .I(N__10168));
    CascadeMux I__1120 (
            .O(N__10171),
            .I(N__10165));
    CascadeBuf I__1119 (
            .O(N__10168),
            .I(N__10162));
    CascadeBuf I__1118 (
            .O(N__10165),
            .I(N__10159));
    CascadeMux I__1117 (
            .O(N__10162),
            .I(N__10156));
    CascadeMux I__1116 (
            .O(N__10159),
            .I(N__10153));
    CascadeBuf I__1115 (
            .O(N__10156),
            .I(N__10150));
    CascadeBuf I__1114 (
            .O(N__10153),
            .I(N__10147));
    CascadeMux I__1113 (
            .O(N__10150),
            .I(N__10144));
    CascadeMux I__1112 (
            .O(N__10147),
            .I(N__10141));
    CascadeBuf I__1111 (
            .O(N__10144),
            .I(N__10138));
    CascadeBuf I__1110 (
            .O(N__10141),
            .I(N__10135));
    CascadeMux I__1109 (
            .O(N__10138),
            .I(N__10132));
    CascadeMux I__1108 (
            .O(N__10135),
            .I(N__10129));
    CascadeBuf I__1107 (
            .O(N__10132),
            .I(N__10126));
    CascadeBuf I__1106 (
            .O(N__10129),
            .I(N__10123));
    CascadeMux I__1105 (
            .O(N__10126),
            .I(N__10120));
    CascadeMux I__1104 (
            .O(N__10123),
            .I(N__10117));
    CascadeBuf I__1103 (
            .O(N__10120),
            .I(N__10114));
    CascadeBuf I__1102 (
            .O(N__10117),
            .I(N__10111));
    CascadeMux I__1101 (
            .O(N__10114),
            .I(N__10108));
    CascadeMux I__1100 (
            .O(N__10111),
            .I(N__10105));
    CascadeBuf I__1099 (
            .O(N__10108),
            .I(N__10102));
    CascadeBuf I__1098 (
            .O(N__10105),
            .I(N__10099));
    CascadeMux I__1097 (
            .O(N__10102),
            .I(N__10096));
    CascadeMux I__1096 (
            .O(N__10099),
            .I(N__10093));
    CascadeBuf I__1095 (
            .O(N__10096),
            .I(N__10090));
    CascadeBuf I__1094 (
            .O(N__10093),
            .I(N__10087));
    CascadeMux I__1093 (
            .O(N__10090),
            .I(N__10084));
    CascadeMux I__1092 (
            .O(N__10087),
            .I(N__10081));
    CascadeBuf I__1091 (
            .O(N__10084),
            .I(N__10078));
    CascadeBuf I__1090 (
            .O(N__10081),
            .I(N__10075));
    CascadeMux I__1089 (
            .O(N__10078),
            .I(N__10072));
    CascadeMux I__1088 (
            .O(N__10075),
            .I(N__10069));
    CascadeBuf I__1087 (
            .O(N__10072),
            .I(N__10066));
    CascadeBuf I__1086 (
            .O(N__10069),
            .I(N__10063));
    CascadeMux I__1085 (
            .O(N__10066),
            .I(N__10060));
    CascadeMux I__1084 (
            .O(N__10063),
            .I(N__10057));
    CascadeBuf I__1083 (
            .O(N__10060),
            .I(N__10054));
    CascadeBuf I__1082 (
            .O(N__10057),
            .I(N__10051));
    CascadeMux I__1081 (
            .O(N__10054),
            .I(N__10048));
    CascadeMux I__1080 (
            .O(N__10051),
            .I(N__10045));
    CascadeBuf I__1079 (
            .O(N__10048),
            .I(N__10042));
    CascadeBuf I__1078 (
            .O(N__10045),
            .I(N__10039));
    CascadeMux I__1077 (
            .O(N__10042),
            .I(N__10036));
    CascadeMux I__1076 (
            .O(N__10039),
            .I(N__10033));
    InMux I__1075 (
            .O(N__10036),
            .I(N__10030));
    InMux I__1074 (
            .O(N__10033),
            .I(N__10027));
    LocalMux I__1073 (
            .O(N__10030),
            .I(N__10024));
    LocalMux I__1072 (
            .O(N__10027),
            .I(N__10021));
    Span4Mux_v I__1071 (
            .O(N__10024),
            .I(N__10018));
    Span12Mux_v I__1070 (
            .O(N__10021),
            .I(N__10015));
    Span4Mux_v I__1069 (
            .O(N__10018),
            .I(N__10012));
    Span12Mux_h I__1068 (
            .O(N__10015),
            .I(N__10009));
    Span4Mux_v I__1067 (
            .O(N__10012),
            .I(N__10006));
    Odrv12 I__1066 (
            .O(N__10009),
            .I(n20));
    Odrv4 I__1065 (
            .O(N__10006),
            .I(n20));
    InMux I__1064 (
            .O(N__10001),
            .I(N__9998));
    LocalMux I__1063 (
            .O(N__9998),
            .I(N__9995));
    Span4Mux_h I__1062 (
            .O(N__9995),
            .I(N__9992));
    Odrv4 I__1061 (
            .O(N__9992),
            .I(\tvp_video_buffer.BUFFER_1_2 ));
    InMux I__1060 (
            .O(N__9989),
            .I(N__9985));
    InMux I__1059 (
            .O(N__9988),
            .I(N__9981));
    LocalMux I__1058 (
            .O(N__9985),
            .I(N__9978));
    InMux I__1057 (
            .O(N__9984),
            .I(N__9975));
    LocalMux I__1056 (
            .O(N__9981),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    Odrv4 I__1055 (
            .O(N__9978),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__1054 (
            .O(N__9975),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    CascadeMux I__1053 (
            .O(N__9968),
            .I(\transmit_module.video_signal_controller.n3485_cascade_ ));
    InMux I__1052 (
            .O(N__9965),
            .I(N__9961));
    InMux I__1051 (
            .O(N__9964),
            .I(N__9957));
    LocalMux I__1050 (
            .O(N__9961),
            .I(N__9954));
    InMux I__1049 (
            .O(N__9960),
            .I(N__9951));
    LocalMux I__1048 (
            .O(N__9957),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    Odrv4 I__1047 (
            .O(N__9954),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__1046 (
            .O(N__9951),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    InMux I__1045 (
            .O(N__9944),
            .I(N__9941));
    LocalMux I__1044 (
            .O(N__9941),
            .I(\transmit_module.video_signal_controller.n3676 ));
    InMux I__1043 (
            .O(N__9938),
            .I(N__9933));
    InMux I__1042 (
            .O(N__9937),
            .I(N__9930));
    InMux I__1041 (
            .O(N__9936),
            .I(N__9927));
    LocalMux I__1040 (
            .O(N__9933),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    LocalMux I__1039 (
            .O(N__9930),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    LocalMux I__1038 (
            .O(N__9927),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    CascadeMux I__1037 (
            .O(N__9920),
            .I(\transmit_module.video_signal_controller.n3464_cascade_ ));
    InMux I__1036 (
            .O(N__9917),
            .I(N__9913));
    InMux I__1035 (
            .O(N__9916),
            .I(N__9910));
    LocalMux I__1034 (
            .O(N__9913),
            .I(\transmit_module.video_signal_controller.n3378 ));
    LocalMux I__1033 (
            .O(N__9910),
            .I(\transmit_module.video_signal_controller.n3378 ));
    InMux I__1032 (
            .O(N__9905),
            .I(N__9902));
    LocalMux I__1031 (
            .O(N__9902),
            .I(N__9899));
    Odrv4 I__1030 (
            .O(N__9899),
            .I(\transmit_module.ADDR_Y_COMPONENT_5 ));
    InMux I__1029 (
            .O(N__9896),
            .I(N__9888));
    InMux I__1028 (
            .O(N__9895),
            .I(N__9888));
    InMux I__1027 (
            .O(N__9894),
            .I(N__9885));
    InMux I__1026 (
            .O(N__9893),
            .I(N__9882));
    LocalMux I__1025 (
            .O(N__9888),
            .I(N__9879));
    LocalMux I__1024 (
            .O(N__9885),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    LocalMux I__1023 (
            .O(N__9882),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    Odrv4 I__1022 (
            .O(N__9879),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    InMux I__1021 (
            .O(N__9872),
            .I(N__9869));
    LocalMux I__1020 (
            .O(N__9869),
            .I(\transmit_module.video_signal_controller.n6_adj_622 ));
    CascadeMux I__1019 (
            .O(N__9866),
            .I(N__9862));
    InMux I__1018 (
            .O(N__9865),
            .I(N__9855));
    InMux I__1017 (
            .O(N__9862),
            .I(N__9855));
    InMux I__1016 (
            .O(N__9861),
            .I(N__9852));
    InMux I__1015 (
            .O(N__9860),
            .I(N__9849));
    LocalMux I__1014 (
            .O(N__9855),
            .I(N__9846));
    LocalMux I__1013 (
            .O(N__9852),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__1012 (
            .O(N__9849),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    Odrv4 I__1011 (
            .O(N__9846),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    InMux I__1010 (
            .O(N__9839),
            .I(N__9835));
    InMux I__1009 (
            .O(N__9838),
            .I(N__9832));
    LocalMux I__1008 (
            .O(N__9835),
            .I(N__9829));
    LocalMux I__1007 (
            .O(N__9832),
            .I(\transmit_module.video_signal_controller.n2019 ));
    Odrv4 I__1006 (
            .O(N__9829),
            .I(\transmit_module.video_signal_controller.n2019 ));
    CEMux I__1005 (
            .O(N__9824),
            .I(N__9819));
    SRMux I__1004 (
            .O(N__9823),
            .I(N__9815));
    SRMux I__1003 (
            .O(N__9822),
            .I(N__9812));
    LocalMux I__1002 (
            .O(N__9819),
            .I(N__9809));
    CEMux I__1001 (
            .O(N__9818),
            .I(N__9806));
    LocalMux I__1000 (
            .O(N__9815),
            .I(N__9803));
    LocalMux I__999 (
            .O(N__9812),
            .I(N__9800));
    Span4Mux_v I__998 (
            .O(N__9809),
            .I(N__9793));
    LocalMux I__997 (
            .O(N__9806),
            .I(N__9793));
    Span4Mux_h I__996 (
            .O(N__9803),
            .I(N__9793));
    Sp12to4 I__995 (
            .O(N__9800),
            .I(N__9790));
    Odrv4 I__994 (
            .O(N__9793),
            .I(\transmit_module.video_signal_controller.n2050 ));
    Odrv12 I__993 (
            .O(N__9790),
            .I(\transmit_module.video_signal_controller.n2050 ));
    CascadeMux I__992 (
            .O(N__9785),
            .I(\transmit_module.video_signal_controller.n2050_cascade_ ));
    SRMux I__991 (
            .O(N__9782),
            .I(N__9779));
    LocalMux I__990 (
            .O(N__9779),
            .I(N__9775));
    SRMux I__989 (
            .O(N__9778),
            .I(N__9772));
    Span4Mux_v I__988 (
            .O(N__9775),
            .I(N__9767));
    LocalMux I__987 (
            .O(N__9772),
            .I(N__9767));
    Odrv4 I__986 (
            .O(N__9767),
            .I(\transmit_module.video_signal_controller.n2398 ));
    InMux I__985 (
            .O(N__9764),
            .I(\transmit_module.video_signal_controller.n3197 ));
    InMux I__984 (
            .O(N__9761),
            .I(\transmit_module.video_signal_controller.n3198 ));
    InMux I__983 (
            .O(N__9758),
            .I(\transmit_module.video_signal_controller.n3199 ));
    InMux I__982 (
            .O(N__9755),
            .I(N__9751));
    InMux I__981 (
            .O(N__9754),
            .I(N__9748));
    LocalMux I__980 (
            .O(N__9751),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    LocalMux I__979 (
            .O(N__9748),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    InMux I__978 (
            .O(N__9743),
            .I(\transmit_module.video_signal_controller.n3200 ));
    InMux I__977 (
            .O(N__9740),
            .I(N__9736));
    InMux I__976 (
            .O(N__9739),
            .I(N__9733));
    LocalMux I__975 (
            .O(N__9736),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    LocalMux I__974 (
            .O(N__9733),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    InMux I__973 (
            .O(N__9728),
            .I(bfn_12_15_0_));
    InMux I__972 (
            .O(N__9725),
            .I(\transmit_module.video_signal_controller.n3202 ));
    InMux I__971 (
            .O(N__9722),
            .I(\transmit_module.video_signal_controller.n3203 ));
    InMux I__970 (
            .O(N__9719),
            .I(\transmit_module.video_signal_controller.n3204 ));
    InMux I__969 (
            .O(N__9716),
            .I(N__9711));
    InMux I__968 (
            .O(N__9715),
            .I(N__9708));
    InMux I__967 (
            .O(N__9714),
            .I(N__9705));
    LocalMux I__966 (
            .O(N__9711),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    LocalMux I__965 (
            .O(N__9708),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    LocalMux I__964 (
            .O(N__9705),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    InMux I__963 (
            .O(N__9698),
            .I(N__9693));
    InMux I__962 (
            .O(N__9697),
            .I(N__9690));
    InMux I__961 (
            .O(N__9696),
            .I(N__9687));
    LocalMux I__960 (
            .O(N__9693),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__959 (
            .O(N__9690),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__958 (
            .O(N__9687),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    InMux I__957 (
            .O(N__9680),
            .I(N__9677));
    LocalMux I__956 (
            .O(N__9677),
            .I(\transmit_module.Y_DELTA_PATTERN_94 ));
    InMux I__955 (
            .O(N__9674),
            .I(N__9671));
    LocalMux I__954 (
            .O(N__9671),
            .I(\transmit_module.Y_DELTA_PATTERN_93 ));
    InMux I__953 (
            .O(N__9668),
            .I(N__9665));
    LocalMux I__952 (
            .O(N__9665),
            .I(\transmit_module.Y_DELTA_PATTERN_92 ));
    InMux I__951 (
            .O(N__9662),
            .I(N__9659));
    LocalMux I__950 (
            .O(N__9659),
            .I(\transmit_module.Y_DELTA_PATTERN_87 ));
    InMux I__949 (
            .O(N__9656),
            .I(N__9653));
    LocalMux I__948 (
            .O(N__9653),
            .I(\transmit_module.Y_DELTA_PATTERN_89 ));
    InMux I__947 (
            .O(N__9650),
            .I(N__9647));
    LocalMux I__946 (
            .O(N__9647),
            .I(\transmit_module.Y_DELTA_PATTERN_88 ));
    InMux I__945 (
            .O(N__9644),
            .I(N__9641));
    LocalMux I__944 (
            .O(N__9641),
            .I(\transmit_module.Y_DELTA_PATTERN_91 ));
    InMux I__943 (
            .O(N__9638),
            .I(N__9635));
    LocalMux I__942 (
            .O(N__9635),
            .I(\transmit_module.Y_DELTA_PATTERN_90 ));
    CEMux I__941 (
            .O(N__9632),
            .I(N__9627));
    CEMux I__940 (
            .O(N__9631),
            .I(N__9624));
    CEMux I__939 (
            .O(N__9630),
            .I(N__9621));
    LocalMux I__938 (
            .O(N__9627),
            .I(N__9618));
    LocalMux I__937 (
            .O(N__9624),
            .I(N__9613));
    LocalMux I__936 (
            .O(N__9621),
            .I(N__9613));
    Span12Mux_h I__935 (
            .O(N__9618),
            .I(N__9610));
    Sp12to4 I__934 (
            .O(N__9613),
            .I(N__9607));
    Odrv12 I__933 (
            .O(N__9610),
            .I(\transmit_module.n2209 ));
    Odrv12 I__932 (
            .O(N__9607),
            .I(\transmit_module.n2209 ));
    InMux I__931 (
            .O(N__9602),
            .I(bfn_12_14_0_));
    InMux I__930 (
            .O(N__9599),
            .I(\transmit_module.video_signal_controller.n3194 ));
    InMux I__929 (
            .O(N__9596),
            .I(\transmit_module.video_signal_controller.n3195 ));
    InMux I__928 (
            .O(N__9593),
            .I(\transmit_module.video_signal_controller.n3196 ));
    InMux I__927 (
            .O(N__9590),
            .I(N__9587));
    LocalMux I__926 (
            .O(N__9587),
            .I(N__9584));
    Span4Mux_v I__925 (
            .O(N__9584),
            .I(N__9581));
    Odrv4 I__924 (
            .O(N__9581),
            .I(\tvp_video_buffer.BUFFER_0_2 ));
    InMux I__923 (
            .O(N__9578),
            .I(N__9575));
    LocalMux I__922 (
            .O(N__9575),
            .I(N__9572));
    Span12Mux_h I__921 (
            .O(N__9572),
            .I(N__9569));
    Odrv12 I__920 (
            .O(N__9569),
            .I(TVP_VIDEO_c_3));
    InMux I__919 (
            .O(N__9566),
            .I(N__9563));
    LocalMux I__918 (
            .O(N__9563),
            .I(\tvp_video_buffer.BUFFER_0_3 ));
    InMux I__917 (
            .O(N__9560),
            .I(N__9557));
    LocalMux I__916 (
            .O(N__9557),
            .I(\transmit_module.X_DELTA_PATTERN_15 ));
    InMux I__915 (
            .O(N__9554),
            .I(N__9551));
    LocalMux I__914 (
            .O(N__9551),
            .I(\transmit_module.X_DELTA_PATTERN_14 ));
    InMux I__913 (
            .O(N__9548),
            .I(\transmit_module.video_signal_controller.n3186 ));
    InMux I__912 (
            .O(N__9545),
            .I(\transmit_module.video_signal_controller.n3187 ));
    InMux I__911 (
            .O(N__9542),
            .I(\transmit_module.video_signal_controller.n3188 ));
    InMux I__910 (
            .O(N__9539),
            .I(\transmit_module.video_signal_controller.n3189 ));
    InMux I__909 (
            .O(N__9536),
            .I(bfn_11_18_0_));
    InMux I__908 (
            .O(N__9533),
            .I(\transmit_module.video_signal_controller.n3191 ));
    InMux I__907 (
            .O(N__9530),
            .I(\transmit_module.video_signal_controller.n3192 ));
    InMux I__906 (
            .O(N__9527),
            .I(\transmit_module.video_signal_controller.n3193 ));
    CEMux I__905 (
            .O(N__9524),
            .I(N__9520));
    CEMux I__904 (
            .O(N__9523),
            .I(N__9517));
    LocalMux I__903 (
            .O(N__9520),
            .I(N__9509));
    LocalMux I__902 (
            .O(N__9517),
            .I(N__9506));
    CEMux I__901 (
            .O(N__9516),
            .I(N__9503));
    CEMux I__900 (
            .O(N__9515),
            .I(N__9499));
    CEMux I__899 (
            .O(N__9514),
            .I(N__9492));
    CEMux I__898 (
            .O(N__9513),
            .I(N__9489));
    CEMux I__897 (
            .O(N__9512),
            .I(N__9486));
    Span4Mux_v I__896 (
            .O(N__9509),
            .I(N__9477));
    Span4Mux_h I__895 (
            .O(N__9506),
            .I(N__9477));
    LocalMux I__894 (
            .O(N__9503),
            .I(N__9477));
    CEMux I__893 (
            .O(N__9502),
            .I(N__9474));
    LocalMux I__892 (
            .O(N__9499),
            .I(N__9471));
    CEMux I__891 (
            .O(N__9498),
            .I(N__9468));
    CEMux I__890 (
            .O(N__9497),
            .I(N__9465));
    CEMux I__889 (
            .O(N__9496),
            .I(N__9462));
    CEMux I__888 (
            .O(N__9495),
            .I(N__9459));
    LocalMux I__887 (
            .O(N__9492),
            .I(N__9456));
    LocalMux I__886 (
            .O(N__9489),
            .I(N__9451));
    LocalMux I__885 (
            .O(N__9486),
            .I(N__9451));
    CEMux I__884 (
            .O(N__9485),
            .I(N__9448));
    CEMux I__883 (
            .O(N__9484),
            .I(N__9445));
    Span4Mux_v I__882 (
            .O(N__9477),
            .I(N__9442));
    LocalMux I__881 (
            .O(N__9474),
            .I(N__9435));
    Span4Mux_h I__880 (
            .O(N__9471),
            .I(N__9435));
    LocalMux I__879 (
            .O(N__9468),
            .I(N__9435));
    LocalMux I__878 (
            .O(N__9465),
            .I(N__9428));
    LocalMux I__877 (
            .O(N__9462),
            .I(N__9428));
    LocalMux I__876 (
            .O(N__9459),
            .I(N__9428));
    Span4Mux_h I__875 (
            .O(N__9456),
            .I(N__9421));
    Span4Mux_h I__874 (
            .O(N__9451),
            .I(N__9421));
    LocalMux I__873 (
            .O(N__9448),
            .I(N__9421));
    LocalMux I__872 (
            .O(N__9445),
            .I(N__9418));
    Span4Mux_h I__871 (
            .O(N__9442),
            .I(N__9415));
    Span4Mux_v I__870 (
            .O(N__9435),
            .I(N__9412));
    Sp12to4 I__869 (
            .O(N__9428),
            .I(N__9409));
    Sp12to4 I__868 (
            .O(N__9421),
            .I(N__9406));
    Span4Mux_h I__867 (
            .O(N__9418),
            .I(N__9403));
    Odrv4 I__866 (
            .O(N__9415),
            .I(\transmit_module.n3683 ));
    Odrv4 I__865 (
            .O(N__9412),
            .I(\transmit_module.n3683 ));
    Odrv12 I__864 (
            .O(N__9409),
            .I(\transmit_module.n3683 ));
    Odrv12 I__863 (
            .O(N__9406),
            .I(\transmit_module.n3683 ));
    Odrv4 I__862 (
            .O(N__9403),
            .I(\transmit_module.n3683 ));
    CascadeMux I__861 (
            .O(N__9392),
            .I(\transmit_module.video_signal_controller.n6_cascade_ ));
    InMux I__860 (
            .O(N__9389),
            .I(N__9386));
    LocalMux I__859 (
            .O(N__9386),
            .I(\transmit_module.ADDR_Y_COMPONENT_11 ));
    InMux I__858 (
            .O(N__9383),
            .I(N__9380));
    LocalMux I__857 (
            .O(N__9380),
            .I(N__9377));
    Odrv4 I__856 (
            .O(N__9377),
            .I(\transmit_module.ADDR_Y_COMPONENT_12 ));
    InMux I__855 (
            .O(N__9374),
            .I(bfn_11_17_0_));
    InMux I__854 (
            .O(N__9371),
            .I(\transmit_module.video_signal_controller.n3183 ));
    InMux I__853 (
            .O(N__9368),
            .I(\transmit_module.video_signal_controller.n3184 ));
    InMux I__852 (
            .O(N__9365),
            .I(\transmit_module.video_signal_controller.n3185 ));
    InMux I__851 (
            .O(N__9362),
            .I(N__9359));
    LocalMux I__850 (
            .O(N__9359),
            .I(N__9356));
    Span4Mux_h I__849 (
            .O(N__9356),
            .I(N__9353));
    Odrv4 I__848 (
            .O(N__9353),
            .I(\transmit_module.Y_DELTA_PATTERN_99 ));
    InMux I__847 (
            .O(N__9350),
            .I(N__9347));
    LocalMux I__846 (
            .O(N__9347),
            .I(\transmit_module.Y_DELTA_PATTERN_98 ));
    InMux I__845 (
            .O(N__9344),
            .I(N__9341));
    LocalMux I__844 (
            .O(N__9341),
            .I(\transmit_module.Y_DELTA_PATTERN_97 ));
    InMux I__843 (
            .O(N__9338),
            .I(N__9335));
    LocalMux I__842 (
            .O(N__9335),
            .I(\transmit_module.Y_DELTA_PATTERN_95 ));
    InMux I__841 (
            .O(N__9332),
            .I(N__9329));
    LocalMux I__840 (
            .O(N__9329),
            .I(\transmit_module.Y_DELTA_PATTERN_60 ));
    InMux I__839 (
            .O(N__9326),
            .I(N__9323));
    LocalMux I__838 (
            .O(N__9323),
            .I(\transmit_module.Y_DELTA_PATTERN_59 ));
    InMux I__837 (
            .O(N__9320),
            .I(N__9317));
    LocalMux I__836 (
            .O(N__9317),
            .I(\transmit_module.Y_DELTA_PATTERN_58 ));
    InMux I__835 (
            .O(N__9314),
            .I(N__9311));
    LocalMux I__834 (
            .O(N__9311),
            .I(\transmit_module.Y_DELTA_PATTERN_54 ));
    InMux I__833 (
            .O(N__9308),
            .I(N__9305));
    LocalMux I__832 (
            .O(N__9305),
            .I(\transmit_module.Y_DELTA_PATTERN_55 ));
    InMux I__831 (
            .O(N__9302),
            .I(N__9299));
    LocalMux I__830 (
            .O(N__9299),
            .I(\transmit_module.Y_DELTA_PATTERN_57 ));
    InMux I__829 (
            .O(N__9296),
            .I(N__9293));
    LocalMux I__828 (
            .O(N__9293),
            .I(\transmit_module.Y_DELTA_PATTERN_56 ));
    InMux I__827 (
            .O(N__9290),
            .I(N__9287));
    LocalMux I__826 (
            .O(N__9287),
            .I(\transmit_module.Y_DELTA_PATTERN_86 ));
    InMux I__825 (
            .O(N__9284),
            .I(N__9281));
    LocalMux I__824 (
            .O(N__9281),
            .I(\transmit_module.Y_DELTA_PATTERN_96 ));
    InMux I__823 (
            .O(N__9278),
            .I(N__9275));
    LocalMux I__822 (
            .O(N__9275),
            .I(\transmit_module.Y_DELTA_PATTERN_47 ));
    InMux I__821 (
            .O(N__9272),
            .I(N__9269));
    LocalMux I__820 (
            .O(N__9269),
            .I(\transmit_module.Y_DELTA_PATTERN_46 ));
    InMux I__819 (
            .O(N__9266),
            .I(N__9263));
    LocalMux I__818 (
            .O(N__9263),
            .I(\transmit_module.Y_DELTA_PATTERN_49 ));
    InMux I__817 (
            .O(N__9260),
            .I(N__9257));
    LocalMux I__816 (
            .O(N__9257),
            .I(\transmit_module.Y_DELTA_PATTERN_48 ));
    InMux I__815 (
            .O(N__9254),
            .I(N__9251));
    LocalMux I__814 (
            .O(N__9251),
            .I(N__9248));
    Odrv12 I__813 (
            .O(N__9248),
            .I(\transmit_module.Y_DELTA_PATTERN_53 ));
    InMux I__812 (
            .O(N__9245),
            .I(N__9242));
    LocalMux I__811 (
            .O(N__9242),
            .I(\transmit_module.Y_DELTA_PATTERN_52 ));
    InMux I__810 (
            .O(N__9239),
            .I(N__9236));
    LocalMux I__809 (
            .O(N__9236),
            .I(\transmit_module.Y_DELTA_PATTERN_51 ));
    InMux I__808 (
            .O(N__9233),
            .I(N__9230));
    LocalMux I__807 (
            .O(N__9230),
            .I(\transmit_module.Y_DELTA_PATTERN_50 ));
    InMux I__806 (
            .O(N__9227),
            .I(N__9224));
    LocalMux I__805 (
            .O(N__9224),
            .I(\transmit_module.Y_DELTA_PATTERN_82 ));
    InMux I__804 (
            .O(N__9221),
            .I(N__9218));
    LocalMux I__803 (
            .O(N__9218),
            .I(\transmit_module.Y_DELTA_PATTERN_81 ));
    InMux I__802 (
            .O(N__9215),
            .I(N__9212));
    LocalMux I__801 (
            .O(N__9212),
            .I(\transmit_module.Y_DELTA_PATTERN_83 ));
    InMux I__800 (
            .O(N__9209),
            .I(N__9206));
    LocalMux I__799 (
            .O(N__9206),
            .I(\transmit_module.Y_DELTA_PATTERN_85 ));
    InMux I__798 (
            .O(N__9203),
            .I(N__9200));
    LocalMux I__797 (
            .O(N__9200),
            .I(\transmit_module.Y_DELTA_PATTERN_84 ));
    InMux I__796 (
            .O(N__9197),
            .I(N__9194));
    LocalMux I__795 (
            .O(N__9194),
            .I(\transmit_module.Y_DELTA_PATTERN_26 ));
    InMux I__794 (
            .O(N__9191),
            .I(N__9188));
    LocalMux I__793 (
            .O(N__9188),
            .I(\transmit_module.Y_DELTA_PATTERN_27 ));
    InMux I__792 (
            .O(N__9185),
            .I(N__9182));
    LocalMux I__791 (
            .O(N__9182),
            .I(\transmit_module.Y_DELTA_PATTERN_28 ));
    InMux I__790 (
            .O(N__9179),
            .I(N__9176));
    LocalMux I__789 (
            .O(N__9176),
            .I(N__9173));
    Odrv12 I__788 (
            .O(N__9173),
            .I(\transmit_module.Y_DELTA_PATTERN_30 ));
    InMux I__787 (
            .O(N__9170),
            .I(N__9167));
    LocalMux I__786 (
            .O(N__9167),
            .I(\transmit_module.Y_DELTA_PATTERN_29 ));
    InMux I__785 (
            .O(N__9164),
            .I(N__9161));
    LocalMux I__784 (
            .O(N__9161),
            .I(\transmit_module.Y_DELTA_PATTERN_75 ));
    InMux I__783 (
            .O(N__9158),
            .I(N__9155));
    LocalMux I__782 (
            .O(N__9155),
            .I(\transmit_module.Y_DELTA_PATTERN_78 ));
    InMux I__781 (
            .O(N__9152),
            .I(N__9149));
    LocalMux I__780 (
            .O(N__9149),
            .I(\transmit_module.Y_DELTA_PATTERN_79 ));
    InMux I__779 (
            .O(N__9146),
            .I(N__9143));
    LocalMux I__778 (
            .O(N__9143),
            .I(\transmit_module.Y_DELTA_PATTERN_77 ));
    InMux I__777 (
            .O(N__9140),
            .I(N__9137));
    LocalMux I__776 (
            .O(N__9137),
            .I(\transmit_module.Y_DELTA_PATTERN_76 ));
    InMux I__775 (
            .O(N__9134),
            .I(N__9131));
    LocalMux I__774 (
            .O(N__9131),
            .I(\transmit_module.Y_DELTA_PATTERN_62 ));
    InMux I__773 (
            .O(N__9128),
            .I(N__9125));
    LocalMux I__772 (
            .O(N__9125),
            .I(\transmit_module.Y_DELTA_PATTERN_61 ));
    InMux I__771 (
            .O(N__9122),
            .I(N__9119));
    LocalMux I__770 (
            .O(N__9119),
            .I(N__9116));
    Odrv12 I__769 (
            .O(N__9116),
            .I(\transmit_module.Y_DELTA_PATTERN_80 ));
    InMux I__768 (
            .O(N__9113),
            .I(N__9110));
    LocalMux I__767 (
            .O(N__9110),
            .I(\transmit_module.Y_DELTA_PATTERN_45 ));
    IoInMux I__766 (
            .O(N__9107),
            .I(N__9104));
    LocalMux I__765 (
            .O(N__9104),
            .I(N__9101));
    IoSpan4Mux I__764 (
            .O(N__9101),
            .I(N__9098));
    Span4Mux_s3_h I__763 (
            .O(N__9098),
            .I(N__9094));
    InMux I__762 (
            .O(N__9097),
            .I(N__9091));
    Span4Mux_h I__761 (
            .O(N__9094),
            .I(N__9086));
    LocalMux I__760 (
            .O(N__9091),
            .I(N__9086));
    Span4Mux_h I__759 (
            .O(N__9086),
            .I(N__9083));
    Sp12to4 I__758 (
            .O(N__9083),
            .I(N__9080));
    Span12Mux_v I__757 (
            .O(N__9080),
            .I(N__9077));
    Odrv12 I__756 (
            .O(N__9077),
            .I(DEBUG_c_5_c));
    InMux I__755 (
            .O(N__9074),
            .I(N__9071));
    LocalMux I__754 (
            .O(N__9071),
            .I(N__9065));
    InMux I__753 (
            .O(N__9070),
            .I(N__9062));
    InMux I__752 (
            .O(N__9069),
            .I(N__9059));
    InMux I__751 (
            .O(N__9068),
            .I(N__9054));
    Span4Mux_h I__750 (
            .O(N__9065),
            .I(N__9051));
    LocalMux I__749 (
            .O(N__9062),
            .I(N__9048));
    LocalMux I__748 (
            .O(N__9059),
            .I(N__9045));
    InMux I__747 (
            .O(N__9058),
            .I(N__9042));
    InMux I__746 (
            .O(N__9057),
            .I(N__9039));
    LocalMux I__745 (
            .O(N__9054),
            .I(N__9035));
    Span4Mux_v I__744 (
            .O(N__9051),
            .I(N__9032));
    Span4Mux_v I__743 (
            .O(N__9048),
            .I(N__9027));
    Span4Mux_v I__742 (
            .O(N__9045),
            .I(N__9027));
    LocalMux I__741 (
            .O(N__9042),
            .I(N__9024));
    LocalMux I__740 (
            .O(N__9039),
            .I(N__9021));
    InMux I__739 (
            .O(N__9038),
            .I(N__9018));
    Span12Mux_h I__738 (
            .O(N__9035),
            .I(N__9015));
    Span4Mux_v I__737 (
            .O(N__9032),
            .I(N__9010));
    Span4Mux_h I__736 (
            .O(N__9027),
            .I(N__9010));
    Span12Mux_s3_v I__735 (
            .O(N__9024),
            .I(N__9007));
    Span12Mux_s4_v I__734 (
            .O(N__9021),
            .I(N__9002));
    LocalMux I__733 (
            .O(N__9018),
            .I(N__9002));
    Span12Mux_v I__732 (
            .O(N__9015),
            .I(N__8992));
    Sp12to4 I__731 (
            .O(N__9010),
            .I(N__8992));
    Span12Mux_v I__730 (
            .O(N__9007),
            .I(N__8992));
    Span12Mux_v I__729 (
            .O(N__9002),
            .I(N__8992));
    InMux I__728 (
            .O(N__9001),
            .I(N__8989));
    Odrv12 I__727 (
            .O(N__8992),
            .I(RX_DATA_3));
    LocalMux I__726 (
            .O(N__8989),
            .I(RX_DATA_3));
    InMux I__725 (
            .O(N__8984),
            .I(N__8981));
    LocalMux I__724 (
            .O(N__8981),
            .I(\tvp_video_buffer.BUFFER_0_5 ));
    InMux I__723 (
            .O(N__8978),
            .I(N__8975));
    LocalMux I__722 (
            .O(N__8975),
            .I(\tvp_video_buffer.BUFFER_1_5 ));
    CascadeMux I__721 (
            .O(N__8972),
            .I(N__8969));
    CascadeBuf I__720 (
            .O(N__8969),
            .I(N__8965));
    CascadeMux I__719 (
            .O(N__8968),
            .I(N__8962));
    CascadeMux I__718 (
            .O(N__8965),
            .I(N__8959));
    CascadeBuf I__717 (
            .O(N__8962),
            .I(N__8956));
    CascadeBuf I__716 (
            .O(N__8959),
            .I(N__8953));
    CascadeMux I__715 (
            .O(N__8956),
            .I(N__8950));
    CascadeMux I__714 (
            .O(N__8953),
            .I(N__8947));
    CascadeBuf I__713 (
            .O(N__8950),
            .I(N__8944));
    CascadeBuf I__712 (
            .O(N__8947),
            .I(N__8941));
    CascadeMux I__711 (
            .O(N__8944),
            .I(N__8938));
    CascadeMux I__710 (
            .O(N__8941),
            .I(N__8935));
    CascadeBuf I__709 (
            .O(N__8938),
            .I(N__8932));
    CascadeBuf I__708 (
            .O(N__8935),
            .I(N__8929));
    CascadeMux I__707 (
            .O(N__8932),
            .I(N__8926));
    CascadeMux I__706 (
            .O(N__8929),
            .I(N__8923));
    CascadeBuf I__705 (
            .O(N__8926),
            .I(N__8920));
    CascadeBuf I__704 (
            .O(N__8923),
            .I(N__8917));
    CascadeMux I__703 (
            .O(N__8920),
            .I(N__8914));
    CascadeMux I__702 (
            .O(N__8917),
            .I(N__8911));
    CascadeBuf I__701 (
            .O(N__8914),
            .I(N__8908));
    CascadeBuf I__700 (
            .O(N__8911),
            .I(N__8905));
    CascadeMux I__699 (
            .O(N__8908),
            .I(N__8902));
    CascadeMux I__698 (
            .O(N__8905),
            .I(N__8899));
    CascadeBuf I__697 (
            .O(N__8902),
            .I(N__8896));
    CascadeBuf I__696 (
            .O(N__8899),
            .I(N__8893));
    CascadeMux I__695 (
            .O(N__8896),
            .I(N__8890));
    CascadeMux I__694 (
            .O(N__8893),
            .I(N__8887));
    CascadeBuf I__693 (
            .O(N__8890),
            .I(N__8884));
    CascadeBuf I__692 (
            .O(N__8887),
            .I(N__8881));
    CascadeMux I__691 (
            .O(N__8884),
            .I(N__8878));
    CascadeMux I__690 (
            .O(N__8881),
            .I(N__8875));
    CascadeBuf I__689 (
            .O(N__8878),
            .I(N__8872));
    CascadeBuf I__688 (
            .O(N__8875),
            .I(N__8869));
    CascadeMux I__687 (
            .O(N__8872),
            .I(N__8866));
    CascadeMux I__686 (
            .O(N__8869),
            .I(N__8863));
    CascadeBuf I__685 (
            .O(N__8866),
            .I(N__8860));
    CascadeBuf I__684 (
            .O(N__8863),
            .I(N__8857));
    CascadeMux I__683 (
            .O(N__8860),
            .I(N__8854));
    CascadeMux I__682 (
            .O(N__8857),
            .I(N__8851));
    CascadeBuf I__681 (
            .O(N__8854),
            .I(N__8848));
    CascadeBuf I__680 (
            .O(N__8851),
            .I(N__8845));
    CascadeMux I__679 (
            .O(N__8848),
            .I(N__8842));
    CascadeMux I__678 (
            .O(N__8845),
            .I(N__8839));
    CascadeBuf I__677 (
            .O(N__8842),
            .I(N__8836));
    CascadeBuf I__676 (
            .O(N__8839),
            .I(N__8833));
    CascadeMux I__675 (
            .O(N__8836),
            .I(N__8830));
    CascadeMux I__674 (
            .O(N__8833),
            .I(N__8827));
    CascadeBuf I__673 (
            .O(N__8830),
            .I(N__8824));
    CascadeBuf I__672 (
            .O(N__8827),
            .I(N__8821));
    CascadeMux I__671 (
            .O(N__8824),
            .I(N__8818));
    CascadeMux I__670 (
            .O(N__8821),
            .I(N__8815));
    CascadeBuf I__669 (
            .O(N__8818),
            .I(N__8812));
    CascadeBuf I__668 (
            .O(N__8815),
            .I(N__8809));
    CascadeMux I__667 (
            .O(N__8812),
            .I(N__8806));
    CascadeMux I__666 (
            .O(N__8809),
            .I(N__8803));
    CascadeBuf I__665 (
            .O(N__8806),
            .I(N__8800));
    CascadeBuf I__664 (
            .O(N__8803),
            .I(N__8797));
    CascadeMux I__663 (
            .O(N__8800),
            .I(N__8794));
    CascadeMux I__662 (
            .O(N__8797),
            .I(N__8791));
    CascadeBuf I__661 (
            .O(N__8794),
            .I(N__8788));
    InMux I__660 (
            .O(N__8791),
            .I(N__8785));
    CascadeMux I__659 (
            .O(N__8788),
            .I(N__8782));
    LocalMux I__658 (
            .O(N__8785),
            .I(N__8779));
    InMux I__657 (
            .O(N__8782),
            .I(N__8776));
    Span4Mux_h I__656 (
            .O(N__8779),
            .I(N__8773));
    LocalMux I__655 (
            .O(N__8776),
            .I(N__8770));
    Span4Mux_v I__654 (
            .O(N__8773),
            .I(N__8767));
    Sp12to4 I__653 (
            .O(N__8770),
            .I(N__8764));
    Sp12to4 I__652 (
            .O(N__8767),
            .I(N__8761));
    Span12Mux_s5_v I__651 (
            .O(N__8764),
            .I(N__8756));
    Span12Mux_h I__650 (
            .O(N__8761),
            .I(N__8756));
    Odrv12 I__649 (
            .O(N__8756),
            .I(n27));
    InMux I__648 (
            .O(N__8753),
            .I(N__8750));
    LocalMux I__647 (
            .O(N__8750),
            .I(N__8747));
    Span4Mux_v I__646 (
            .O(N__8747),
            .I(N__8744));
    Odrv4 I__645 (
            .O(N__8744),
            .I(\line_buffer.n603 ));
    InMux I__644 (
            .O(N__8741),
            .I(N__8738));
    LocalMux I__643 (
            .O(N__8738),
            .I(N__8735));
    Span4Mux_v I__642 (
            .O(N__8735),
            .I(N__8732));
    Odrv4 I__641 (
            .O(N__8732),
            .I(\line_buffer.n595 ));
    InMux I__640 (
            .O(N__8729),
            .I(N__8726));
    LocalMux I__639 (
            .O(N__8726),
            .I(N__8723));
    Span4Mux_v I__638 (
            .O(N__8723),
            .I(N__8720));
    Odrv4 I__637 (
            .O(N__8720),
            .I(\line_buffer.n602 ));
    InMux I__636 (
            .O(N__8717),
            .I(N__8714));
    LocalMux I__635 (
            .O(N__8714),
            .I(N__8711));
    Span4Mux_v I__634 (
            .O(N__8711),
            .I(N__8708));
    Odrv4 I__633 (
            .O(N__8708),
            .I(\line_buffer.n594 ));
    InMux I__632 (
            .O(N__8705),
            .I(N__8702));
    LocalMux I__631 (
            .O(N__8702),
            .I(N__8699));
    IoSpan4Mux I__630 (
            .O(N__8699),
            .I(N__8696));
    Odrv4 I__629 (
            .O(N__8696),
            .I(TVP_VIDEO_c_2));
    InMux I__628 (
            .O(N__8693),
            .I(N__8690));
    LocalMux I__627 (
            .O(N__8690),
            .I(\transmit_module.Y_DELTA_PATTERN_74 ));
    InMux I__626 (
            .O(N__8687),
            .I(N__8684));
    LocalMux I__625 (
            .O(N__8684),
            .I(\transmit_module.Y_DELTA_PATTERN_67 ));
    InMux I__624 (
            .O(N__8681),
            .I(N__8678));
    LocalMux I__623 (
            .O(N__8678),
            .I(\transmit_module.Y_DELTA_PATTERN_65 ));
    InMux I__622 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__621 (
            .O(N__8672),
            .I(\transmit_module.Y_DELTA_PATTERN_64 ));
    InMux I__620 (
            .O(N__8669),
            .I(N__8666));
    LocalMux I__619 (
            .O(N__8666),
            .I(\transmit_module.Y_DELTA_PATTERN_69 ));
    InMux I__618 (
            .O(N__8663),
            .I(N__8660));
    LocalMux I__617 (
            .O(N__8660),
            .I(\transmit_module.Y_DELTA_PATTERN_68 ));
    InMux I__616 (
            .O(N__8657),
            .I(N__8654));
    LocalMux I__615 (
            .O(N__8654),
            .I(N__8651));
    Odrv4 I__614 (
            .O(N__8651),
            .I(\transmit_module.Y_DELTA_PATTERN_24 ));
    InMux I__613 (
            .O(N__8648),
            .I(N__8645));
    LocalMux I__612 (
            .O(N__8645),
            .I(\transmit_module.Y_DELTA_PATTERN_25 ));
    InMux I__611 (
            .O(N__8642),
            .I(N__8639));
    LocalMux I__610 (
            .O(N__8639),
            .I(\transmit_module.Y_DELTA_PATTERN_43 ));
    InMux I__609 (
            .O(N__8636),
            .I(N__8633));
    LocalMux I__608 (
            .O(N__8633),
            .I(N__8630));
    Odrv4 I__607 (
            .O(N__8630),
            .I(\transmit_module.Y_DELTA_PATTERN_42 ));
    InMux I__606 (
            .O(N__8627),
            .I(N__8624));
    LocalMux I__605 (
            .O(N__8624),
            .I(\transmit_module.Y_DELTA_PATTERN_44 ));
    InMux I__604 (
            .O(N__8621),
            .I(N__8618));
    LocalMux I__603 (
            .O(N__8618),
            .I(\transmit_module.Y_DELTA_PATTERN_73 ));
    InMux I__602 (
            .O(N__8615),
            .I(N__8612));
    LocalMux I__601 (
            .O(N__8612),
            .I(\transmit_module.Y_DELTA_PATTERN_72 ));
    InMux I__600 (
            .O(N__8609),
            .I(N__8606));
    LocalMux I__599 (
            .O(N__8606),
            .I(\transmit_module.Y_DELTA_PATTERN_63 ));
    InMux I__598 (
            .O(N__8603),
            .I(N__8600));
    LocalMux I__597 (
            .O(N__8600),
            .I(N__8597));
    Odrv4 I__596 (
            .O(N__8597),
            .I(\transmit_module.Y_DELTA_PATTERN_71 ));
    InMux I__595 (
            .O(N__8594),
            .I(N__8591));
    LocalMux I__594 (
            .O(N__8591),
            .I(\transmit_module.Y_DELTA_PATTERN_70 ));
    InMux I__593 (
            .O(N__8588),
            .I(N__8585));
    LocalMux I__592 (
            .O(N__8585),
            .I(\transmit_module.Y_DELTA_PATTERN_66 ));
    InMux I__591 (
            .O(N__8582),
            .I(N__8579));
    LocalMux I__590 (
            .O(N__8579),
            .I(\transmit_module.Y_DELTA_PATTERN_14 ));
    InMux I__589 (
            .O(N__8576),
            .I(N__8573));
    LocalMux I__588 (
            .O(N__8573),
            .I(\transmit_module.Y_DELTA_PATTERN_39 ));
    InMux I__587 (
            .O(N__8570),
            .I(N__8567));
    LocalMux I__586 (
            .O(N__8567),
            .I(\transmit_module.Y_DELTA_PATTERN_41 ));
    InMux I__585 (
            .O(N__8564),
            .I(N__8561));
    LocalMux I__584 (
            .O(N__8561),
            .I(\transmit_module.Y_DELTA_PATTERN_40 ));
    InMux I__583 (
            .O(N__8558),
            .I(N__8555));
    LocalMux I__582 (
            .O(N__8555),
            .I(N__8552));
    Odrv4 I__581 (
            .O(N__8552),
            .I(\transmit_module.Y_DELTA_PATTERN_13 ));
    InMux I__580 (
            .O(N__8549),
            .I(N__8546));
    LocalMux I__579 (
            .O(N__8546),
            .I(\transmit_module.Y_DELTA_PATTERN_12 ));
    InMux I__578 (
            .O(N__8543),
            .I(N__8540));
    LocalMux I__577 (
            .O(N__8540),
            .I(\transmit_module.Y_DELTA_PATTERN_7 ));
    InMux I__576 (
            .O(N__8537),
            .I(N__8534));
    LocalMux I__575 (
            .O(N__8534),
            .I(\transmit_module.Y_DELTA_PATTERN_6 ));
    InMux I__574 (
            .O(N__8531),
            .I(N__8528));
    LocalMux I__573 (
            .O(N__8528),
            .I(\transmit_module.Y_DELTA_PATTERN_11 ));
    InMux I__572 (
            .O(N__8525),
            .I(N__8522));
    LocalMux I__571 (
            .O(N__8522),
            .I(\transmit_module.Y_DELTA_PATTERN_10 ));
    InMux I__570 (
            .O(N__8519),
            .I(N__8516));
    LocalMux I__569 (
            .O(N__8516),
            .I(\transmit_module.Y_DELTA_PATTERN_22 ));
    InMux I__568 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__567 (
            .O(N__8510),
            .I(\transmit_module.Y_DELTA_PATTERN_21 ));
    InMux I__566 (
            .O(N__8507),
            .I(N__8504));
    LocalMux I__565 (
            .O(N__8504),
            .I(\transmit_module.Y_DELTA_PATTERN_20 ));
    InMux I__564 (
            .O(N__8501),
            .I(N__8498));
    LocalMux I__563 (
            .O(N__8498),
            .I(\transmit_module.Y_DELTA_PATTERN_19 ));
    InMux I__562 (
            .O(N__8495),
            .I(N__8492));
    LocalMux I__561 (
            .O(N__8492),
            .I(\transmit_module.Y_DELTA_PATTERN_18 ));
    InMux I__560 (
            .O(N__8489),
            .I(N__8486));
    LocalMux I__559 (
            .O(N__8486),
            .I(\transmit_module.Y_DELTA_PATTERN_15 ));
    InMux I__558 (
            .O(N__8483),
            .I(N__8480));
    LocalMux I__557 (
            .O(N__8480),
            .I(N__8477));
    Odrv4 I__556 (
            .O(N__8477),
            .I(\transmit_module.Y_DELTA_PATTERN_23 ));
    InMux I__555 (
            .O(N__8474),
            .I(N__8471));
    LocalMux I__554 (
            .O(N__8471),
            .I(\transmit_module.Y_DELTA_PATTERN_17 ));
    InMux I__553 (
            .O(N__8468),
            .I(N__8465));
    LocalMux I__552 (
            .O(N__8465),
            .I(\transmit_module.Y_DELTA_PATTERN_16 ));
    InMux I__551 (
            .O(N__8462),
            .I(N__8459));
    LocalMux I__550 (
            .O(N__8459),
            .I(\transmit_module.Y_DELTA_PATTERN_31 ));
    InMux I__549 (
            .O(N__8456),
            .I(N__8453));
    LocalMux I__548 (
            .O(N__8453),
            .I(\transmit_module.Y_DELTA_PATTERN_32 ));
    InMux I__547 (
            .O(N__8450),
            .I(N__8447));
    LocalMux I__546 (
            .O(N__8447),
            .I(\transmit_module.Y_DELTA_PATTERN_33 ));
    InMux I__545 (
            .O(N__8444),
            .I(N__8441));
    LocalMux I__544 (
            .O(N__8441),
            .I(\transmit_module.Y_DELTA_PATTERN_38 ));
    InMux I__543 (
            .O(N__8438),
            .I(N__8435));
    LocalMux I__542 (
            .O(N__8435),
            .I(\transmit_module.Y_DELTA_PATTERN_35 ));
    InMux I__541 (
            .O(N__8432),
            .I(N__8429));
    LocalMux I__540 (
            .O(N__8429),
            .I(\transmit_module.Y_DELTA_PATTERN_34 ));
    InMux I__539 (
            .O(N__8426),
            .I(N__8423));
    LocalMux I__538 (
            .O(N__8423),
            .I(\transmit_module.Y_DELTA_PATTERN_9 ));
    InMux I__537 (
            .O(N__8420),
            .I(N__8417));
    LocalMux I__536 (
            .O(N__8417),
            .I(\transmit_module.Y_DELTA_PATTERN_8 ));
    InMux I__535 (
            .O(N__8414),
            .I(N__8411));
    LocalMux I__534 (
            .O(N__8411),
            .I(\transmit_module.Y_DELTA_PATTERN_37 ));
    InMux I__533 (
            .O(N__8408),
            .I(N__8405));
    LocalMux I__532 (
            .O(N__8405),
            .I(\transmit_module.Y_DELTA_PATTERN_36 ));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3201 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3190 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\transmit_module.n3169 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\receive_module.rx_counter.n3182 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3217 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\receive_module.n3156 ),
            .carryinitout(bfn_15_12_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_5_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_5_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_5_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i35_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8408),
            .lcout(\transmit_module.Y_DELTA_PATTERN_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23598),
            .ce(N__9513),
            .sr(N__20061));
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_5_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_5_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i37_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8444),
            .lcout(\transmit_module.Y_DELTA_PATTERN_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23598),
            .ce(N__9513),
            .sr(N__20061));
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_5_15_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_5_15_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_5_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i36_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8414),
            .lcout(\transmit_module.Y_DELTA_PATTERN_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23598),
            .ce(N__9513),
            .sr(N__20061));
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_6_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_6_14_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_6_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i31_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8456),
            .lcout(\transmit_module.Y_DELTA_PATTERN_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23729),
            .ce(N__21426),
            .sr(N__20012));
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_6_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_6_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_6_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i30_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8462),
            .lcout(\transmit_module.Y_DELTA_PATTERN_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23729),
            .ce(N__21426),
            .sr(N__20012));
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_6_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_6_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_6_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i32_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8450),
            .lcout(\transmit_module.Y_DELTA_PATTERN_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23729),
            .ce(N__21426),
            .sr(N__20012));
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_6_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_6_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_6_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i33_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8432),
            .lcout(\transmit_module.Y_DELTA_PATTERN_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23686),
            .ce(N__9514),
            .sr(N__20065));
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_6_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_6_15_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_6_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i38_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8576),
            .lcout(\transmit_module.Y_DELTA_PATTERN_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23686),
            .ce(N__9514),
            .sr(N__20065));
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_6_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_6_15_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i34_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(N__8438),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23686),
            .ce(N__9514),
            .sr(N__20065));
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_6_18_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_6_18_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_6_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i9_LC_6_18_1  (
            .in0(N__8525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23708),
            .ce(N__21429),
            .sr(N__20056));
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_6_18_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_6_18_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_6_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i7_LC_6_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8420),
            .lcout(\transmit_module.Y_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23708),
            .ce(N__21429),
            .sr(N__20056));
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_6_18_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_6_18_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_6_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i8_LC_6_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8426),
            .lcout(\transmit_module.Y_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23708),
            .ce(N__21429),
            .sr(N__20056));
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_7_12_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_7_12_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_7_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i22_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8483),
            .lcout(\transmit_module.Y_DELTA_PATTERN_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23599),
            .ce(N__21382),
            .sr(N__20036));
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_7_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_7_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_7_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i20_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8513),
            .lcout(\transmit_module.Y_DELTA_PATTERN_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23601),
            .ce(N__21430),
            .sr(N__20067));
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_7_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_7_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i21_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8519),
            .lcout(\transmit_module.Y_DELTA_PATTERN_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23601),
            .ce(N__21430),
            .sr(N__20067));
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_7_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_7_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_7_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i19_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8507),
            .lcout(\transmit_module.Y_DELTA_PATTERN_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23601),
            .ce(N__21430),
            .sr(N__20067));
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_7_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_7_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i18_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8501),
            .lcout(\transmit_module.Y_DELTA_PATTERN_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23601),
            .ce(N__21430),
            .sr(N__20067));
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_7_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_7_13_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_7_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i17_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8495),
            .lcout(\transmit_module.Y_DELTA_PATTERN_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23601),
            .ce(N__21430),
            .sr(N__20067));
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_7_14_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_7_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i15_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8468),
            .lcout(\transmit_module.Y_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23703),
            .ce(N__21407),
            .sr(N__20007));
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_7_14_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_7_14_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_7_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i14_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8489),
            .lcout(\transmit_module.Y_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23703),
            .ce(N__21407),
            .sr(N__20007));
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_7_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_7_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i23_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8657),
            .lcout(\transmit_module.Y_DELTA_PATTERN_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23703),
            .ce(N__21407),
            .sr(N__20007));
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_7_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_7_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_7_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i16_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8474),
            .lcout(\transmit_module.Y_DELTA_PATTERN_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23703),
            .ce(N__21407),
            .sr(N__20007));
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_7_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_7_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i13_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8582),
            .lcout(\transmit_module.Y_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23703),
            .ce(N__21407),
            .sr(N__20007));
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_7_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_7_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i39_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8564),
            .lcout(\transmit_module.Y_DELTA_PATTERN_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23634),
            .ce(N__9512),
            .sr(N__20060));
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_7_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_7_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_7_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i41_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8636),
            .lcout(\transmit_module.Y_DELTA_PATTERN_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23634),
            .ce(N__9512),
            .sr(N__20060));
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_7_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_7_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i40_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8570),
            .lcout(\transmit_module.Y_DELTA_PATTERN_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23634),
            .ce(N__9512),
            .sr(N__20060));
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_7_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_7_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_7_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i12_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8558),
            .lcout(\transmit_module.Y_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23709),
            .ce(N__21427),
            .sr(N__20045));
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_7_17_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_7_17_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_7_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i11_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8549),
            .lcout(\transmit_module.Y_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23486),
            .ce(N__21431),
            .sr(N__20069));
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_7_17_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_7_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i5_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8537),
            .lcout(\transmit_module.Y_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23486),
            .ce(N__21431),
            .sr(N__20069));
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_7_17_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_7_17_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_7_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i6_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8543),
            .lcout(\transmit_module.Y_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23486),
            .ce(N__21431),
            .sr(N__20069));
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_7_18_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_7_18_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i10_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__8531),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23648),
            .ce(N__21428),
            .sr(N__20049));
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_9_10_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_9_10_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_9_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i71_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8615),
            .lcout(\transmit_module.Y_DELTA_PATTERN_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23715),
            .ce(N__9524),
            .sr(N__20057));
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_9_10_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_9_10_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_9_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i73_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8693),
            .lcout(\transmit_module.Y_DELTA_PATTERN_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23715),
            .ce(N__9524),
            .sr(N__20057));
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_9_10_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_9_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i72_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8621),
            .lcout(\transmit_module.Y_DELTA_PATTERN_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23715),
            .ce(N__9524),
            .sr(N__20057));
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_9_10_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_9_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i78_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9152),
            .lcout(\transmit_module.Y_DELTA_PATTERN_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23715),
            .ce(N__9524),
            .sr(N__20057));
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_9_11_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_9_11_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_9_11_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i62_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__8609),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23600),
            .ce(N__9523),
            .sr(N__20044));
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_9_12_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_9_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_9_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i63_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8675),
            .lcout(\transmit_module.Y_DELTA_PATTERN_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23687),
            .ce(N__9516),
            .sr(N__20011));
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_9_12_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_9_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i69_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8594),
            .lcout(\transmit_module.Y_DELTA_PATTERN_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23687),
            .ce(N__9516),
            .sr(N__20011));
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_9_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_9_12_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_9_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i70_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8603),
            .lcout(\transmit_module.Y_DELTA_PATTERN_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23687),
            .ce(N__9516),
            .sr(N__20011));
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_9_13_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_9_13_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_9_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i66_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8687),
            .lcout(\transmit_module.Y_DELTA_PATTERN_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23646),
            .ce(N__9515),
            .sr(N__19994));
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_9_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_9_13_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_9_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i65_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8588),
            .lcout(\transmit_module.Y_DELTA_PATTERN_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23646),
            .ce(N__9515),
            .sr(N__19994));
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_9_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_9_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i67_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8663),
            .lcout(\transmit_module.Y_DELTA_PATTERN_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23646),
            .ce(N__9515),
            .sr(N__19994));
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_9_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_9_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i64_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8681),
            .lcout(\transmit_module.Y_DELTA_PATTERN_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23646),
            .ce(N__9515),
            .sr(N__19994));
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_13_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i68_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8669),
            .lcout(\transmit_module.Y_DELTA_PATTERN_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23646),
            .ce(N__9515),
            .sr(N__19994));
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_9_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i99_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20684),
            .lcout(\transmit_module.Y_DELTA_PATTERN_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23714),
            .ce(N__21381),
            .sr(N__20006));
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_9_14_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_9_14_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_9_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i24_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8648),
            .lcout(\transmit_module.Y_DELTA_PATTERN_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23714),
            .ce(N__21381),
            .sr(N__20006));
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_9_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_9_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_9_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i25_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9197),
            .lcout(\transmit_module.Y_DELTA_PATTERN_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23714),
            .ce(N__21381),
            .sr(N__20006));
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_9_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_9_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_9_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i43_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8627),
            .lcout(\transmit_module.Y_DELTA_PATTERN_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23467),
            .ce(N__9485),
            .sr(N__20019));
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8642),
            .lcout(\transmit_module.Y_DELTA_PATTERN_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23467),
            .ce(N__9485),
            .sr(N__20019));
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9113),
            .lcout(\transmit_module.Y_DELTA_PATTERN_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23467),
            .ce(N__9485),
            .sr(N__20019));
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_9_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_9_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i45_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9272),
            .lcout(\transmit_module.Y_DELTA_PATTERN_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23467),
            .ce(N__9485),
            .sr(N__20019));
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_9_17_1 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_9_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i4_LC_9_17_1  (
            .in0(N__9097),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24148),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_9_17_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_9_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i3_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8978),
            .lcout(RX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24148),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_9_17_7 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_9_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i12_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8984),
            .lcout(\tvp_video_buffer.BUFFER_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24148),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1646_4_lut_LC_9_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1646_4_lut_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1646_4_lut_LC_9_19_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1646_4_lut_LC_9_19_0  (
            .in0(N__20259),
            .in1(N__14165),
            .in2(N__20059),
            .in3(N__13604),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2194_3_lut_LC_9_20_0 .C_ON=1'b0;
    defparam \line_buffer.i2194_3_lut_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2194_3_lut_LC_9_20_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2194_3_lut_LC_9_20_0  (
            .in0(N__24733),
            .in1(N__8753),
            .in2(_gnd_net_),
            .in3(N__8741),
            .lcout(\line_buffer.n3531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2206_3_lut_LC_9_21_5 .C_ON=1'b0;
    defparam \line_buffer.i2206_3_lut_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2206_3_lut_LC_9_21_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2206_3_lut_LC_9_21_5  (
            .in0(N__24779),
            .in1(N__8729),
            .in2(_gnd_net_),
            .in3(N__8717),
            .lcout(\line_buffer.n3543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_10_1_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_10_1_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_10_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i1_LC_10_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8705),
            .lcout(\tvp_video_buffer.BUFFER_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24098),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_10_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_10_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i74_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9164),
            .lcout(\transmit_module.Y_DELTA_PATTERN_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23728),
            .ce(N__9497),
            .sr(N__20068));
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_10_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i75_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9140),
            .lcout(\transmit_module.Y_DELTA_PATTERN_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23728),
            .ce(N__9497),
            .sr(N__20068));
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_10_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_10_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i77_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9158),
            .lcout(\transmit_module.Y_DELTA_PATTERN_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23728),
            .ce(N__9497),
            .sr(N__20068));
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_10_10_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_10_10_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_10_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i79_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9122),
            .lcout(\transmit_module.Y_DELTA_PATTERN_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23728),
            .ce(N__9497),
            .sr(N__20068));
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_10_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_10_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i76_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9146),
            .lcout(\transmit_module.Y_DELTA_PATTERN_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23728),
            .ce(N__9497),
            .sr(N__20068));
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_10_11_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_10_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i61_LC_10_11_1  (
            .in0(N__9134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23677),
            .ce(N__9502),
            .sr(N__20002));
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_10_11_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_10_11_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_10_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i60_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9128),
            .lcout(\transmit_module.Y_DELTA_PATTERN_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23677),
            .ce(N__9502),
            .sr(N__20002));
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_10_11_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_10_11_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_10_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i53_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9314),
            .lcout(\transmit_module.Y_DELTA_PATTERN_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23677),
            .ce(N__9502),
            .sr(N__20002));
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_10_11_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_10_11_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_10_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i80_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9221),
            .lcout(\transmit_module.Y_DELTA_PATTERN_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23677),
            .ce(N__9502),
            .sr(N__20002));
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9215),
            .lcout(\transmit_module.Y_DELTA_PATTERN_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23704),
            .ce(N__9496),
            .sr(N__20050));
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_10_12_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_10_12_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_10_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i81_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9227),
            .lcout(\transmit_module.Y_DELTA_PATTERN_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23704),
            .ce(N__9496),
            .sr(N__20050));
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9203),
            .lcout(\transmit_module.Y_DELTA_PATTERN_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23635),
            .ce(N__9631),
            .sr(N__20001));
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9290),
            .lcout(\transmit_module.Y_DELTA_PATTERN_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23635),
            .ce(N__9631),
            .sr(N__20001));
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9209),
            .lcout(\transmit_module.Y_DELTA_PATTERN_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23635),
            .ce(N__9631),
            .sr(N__20001));
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_10_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_10_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i26_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9191),
            .lcout(\transmit_module.Y_DELTA_PATTERN_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23710),
            .ce(N__21331),
            .sr(N__19876));
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_10_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_10_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_10_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i27_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9185),
            .lcout(\transmit_module.Y_DELTA_PATTERN_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23710),
            .ce(N__21331),
            .sr(N__19876));
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i28_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9170),
            .lcout(\transmit_module.Y_DELTA_PATTERN_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23710),
            .ce(N__21331),
            .sr(N__19876));
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_10_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_10_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i29_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9179),
            .lcout(\transmit_module.Y_DELTA_PATTERN_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23710),
            .ce(N__21331),
            .sr(N__19876));
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i49_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9233),
            .lcout(\transmit_module.Y_DELTA_PATTERN_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23613),
            .ce(N__9484),
            .sr(N__19971));
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9260),
            .lcout(\transmit_module.Y_DELTA_PATTERN_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23613),
            .ce(N__9484),
            .sr(N__19971));
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_10_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_10_15_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_10_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i51_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9245),
            .lcout(\transmit_module.Y_DELTA_PATTERN_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23613),
            .ce(N__9484),
            .sr(N__19971));
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i46_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9278),
            .lcout(\transmit_module.Y_DELTA_PATTERN_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23613),
            .ce(N__9484),
            .sr(N__19971));
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i48_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9266),
            .lcout(\transmit_module.Y_DELTA_PATTERN_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23613),
            .ce(N__9484),
            .sr(N__19971));
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_10_15_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_10_15_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_10_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i52_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9254),
            .lcout(\transmit_module.Y_DELTA_PATTERN_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23613),
            .ce(N__9484),
            .sr(N__19971));
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i50_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9239),
            .lcout(\transmit_module.Y_DELTA_PATTERN_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23613),
            .ce(N__9484),
            .sr(N__19971));
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_10_16_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_10_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i11_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24641),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23649),
            .ce(N__20764),
            .sr(N__19997));
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_10_16_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_10_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_10_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i5_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13538),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23649),
            .ce(N__20764),
            .sr(N__19997));
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_10_19_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_10_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i9_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14216),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23324),
            .ce(N__20772),
            .sr(N__20054));
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_10_20_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_10_20_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_10_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i13_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23918),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23553),
            .ce(N__20774),
            .sr(N__20055));
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_11_11_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_11_11_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_11_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i58_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9326),
            .lcout(\transmit_module.Y_DELTA_PATTERN_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23637),
            .ce(N__9498),
            .sr(N__20043));
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_11_11_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_11_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i59_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9332),
            .lcout(\transmit_module.Y_DELTA_PATTERN_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23637),
            .ce(N__9498),
            .sr(N__20043));
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9320),
            .lcout(\transmit_module.Y_DELTA_PATTERN_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23474),
            .ce(N__9495),
            .sr(N__19964));
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_11_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_11_12_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i54_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9308),
            .lcout(\transmit_module.Y_DELTA_PATTERN_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23474),
            .ce(N__9495),
            .sr(N__19964));
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_11_12_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_11_12_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i55_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9296),
            .lcout(\transmit_module.Y_DELTA_PATTERN_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23474),
            .ce(N__9495),
            .sr(N__19964));
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_12_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i56_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9302),
            .lcout(\transmit_module.Y_DELTA_PATTERN_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23474),
            .ce(N__9495),
            .sr(N__19964));
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9284),
            .lcout(\transmit_module.Y_DELTA_PATTERN_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23602),
            .ce(N__9630),
            .sr(N__20018));
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_11_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_11_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i86_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9662),
            .lcout(\transmit_module.Y_DELTA_PATTERN_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23602),
            .ce(N__9630),
            .sr(N__20018));
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_11_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i96_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9344),
            .lcout(\transmit_module.Y_DELTA_PATTERN_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23602),
            .ce(N__9630),
            .sr(N__20018));
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_11_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_11_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_11_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i98_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9362),
            .lcout(\transmit_module.Y_DELTA_PATTERN_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23602),
            .ce(N__9630),
            .sr(N__20018));
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_11_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_11_13_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i97_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9350),
            .lcout(\transmit_module.Y_DELTA_PATTERN_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23602),
            .ce(N__9630),
            .sr(N__20018));
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9338),
            .lcout(\transmit_module.Y_DELTA_PATTERN_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23602),
            .ce(N__9630),
            .sr(N__20018));
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_11_14_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_11_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i6_LC_11_14_0  (
            .in0(N__15179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23550),
            .ce(N__20738),
            .sr(N__19963));
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_11_14_1 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_11_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i7_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13490),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23550),
            .ce(N__20738),
            .sr(N__19963));
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_11_14_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_11_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i12_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22269),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23550),
            .ce(N__20738),
            .sr(N__19963));
    defparam \transmit_module.video_signal_controller.i2183_3_lut_LC_11_15_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2183_3_lut_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2183_3_lut_LC_11_15_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2183_3_lut_LC_11_15_0  (
            .in0(N__9861),
            .in1(N__9894),
            .in2(_gnd_net_),
            .in3(N__9838),
            .lcout(\transmit_module.video_signal_controller.n3520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i127_2_lut_4_lut_LC_11_15_2 .C_ON=1'b0;
    defparam \transmit_module.i127_2_lut_4_lut_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i127_2_lut_4_lut_LC_11_15_2 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.i127_2_lut_4_lut_LC_11_15_2  (
            .in0(N__11284),
            .in1(N__10870),
            .in2(N__20034),
            .in3(N__10818),
            .lcout(\transmit_module.n2209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i483_2_lut_LC_11_15_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i483_2_lut_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i483_2_lut_LC_11_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i483_2_lut_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__10958),
            .in2(_gnd_net_),
            .in3(N__11009),
            .lcout(\transmit_module.video_signal_controller.n6_adj_622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i127_2_lut_4_lut_rep_24_LC_11_15_4 .C_ON=1'b0;
    defparam \transmit_module.i127_2_lut_4_lut_rep_24_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i127_2_lut_4_lut_rep_24_LC_11_15_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.i127_2_lut_4_lut_rep_24_LC_11_15_4  (
            .in0(N__11285),
            .in1(N__10871),
            .in2(N__20035),
            .in3(N__10819),
            .lcout(\transmit_module.n3683 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_11_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_11_15_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__9754),
            .in2(_gnd_net_),
            .in3(N__9739),
            .lcout(\transmit_module.video_signal_controller.n3378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_15_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_15_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_15_6  (
            .in0(N__9714),
            .in1(N__9696),
            .in2(_gnd_net_),
            .in3(N__9960),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_11_15_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_11_15_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i4_4_lut_LC_11_15_7  (
            .in0(N__9984),
            .in1(N__9936),
            .in2(N__9392),
            .in3(N__9916),
            .lcout(\transmit_module.video_signal_controller.n2019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_11_16_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_11_16_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i0_LC_11_16_1  (
            .in0(N__9389),
            .in1(N__20252),
            .in2(_gnd_net_),
            .in3(N__13655),
            .lcout(TX_ADDR_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23335),
            .ce(N__10246),
            .sr(N__19981));
    defparam \transmit_module.BRAM_ADDR__i12_LC_11_16_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i12_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i12_LC_11_16_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i12_LC_11_16_5  (
            .in0(N__9383),
            .in1(N__20251),
            .in2(_gnd_net_),
            .in3(N__13643),
            .lcout(TX_ADDR_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23335),
            .ce(N__10246),
            .sr(N__19981));
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_11_17_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_11_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i0_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__10276),
            .in2(_gnd_net_),
            .in3(N__9374),
            .lcout(\transmit_module.video_signal_controller.VGA_X_0 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\transmit_module.video_signal_controller.n3183 ),
            .clk(N__23482),
            .ce(),
            .sr(N__9822));
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_11_17_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_11_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i1_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__12458),
            .in2(_gnd_net_),
            .in3(N__9371),
            .lcout(\transmit_module.video_signal_controller.VGA_X_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3183 ),
            .carryout(\transmit_module.video_signal_controller.n3184 ),
            .clk(N__23482),
            .ce(),
            .sr(N__9822));
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_11_17_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_11_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i2_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__12485),
            .in2(_gnd_net_),
            .in3(N__9368),
            .lcout(\transmit_module.video_signal_controller.VGA_X_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3184 ),
            .carryout(\transmit_module.video_signal_controller.n3185 ),
            .clk(N__23482),
            .ce(),
            .sr(N__9822));
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_11_17_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_11_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i3_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__10399),
            .in2(_gnd_net_),
            .in3(N__9365),
            .lcout(\transmit_module.video_signal_controller.VGA_X_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3185 ),
            .carryout(\transmit_module.video_signal_controller.n3186 ),
            .clk(N__23482),
            .ce(),
            .sr(N__9822));
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_11_17_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_11_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i4_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__10379),
            .in2(_gnd_net_),
            .in3(N__9548),
            .lcout(\transmit_module.video_signal_controller.VGA_X_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3186 ),
            .carryout(\transmit_module.video_signal_controller.n3187 ),
            .clk(N__23482),
            .ce(),
            .sr(N__9822));
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_11_17_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_11_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i5_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__10327),
            .in2(_gnd_net_),
            .in3(N__9545),
            .lcout(\transmit_module.video_signal_controller.VGA_X_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3187 ),
            .carryout(\transmit_module.video_signal_controller.n3188 ),
            .clk(N__23482),
            .ce(),
            .sr(N__9822));
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_11_17_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_11_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i6_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__10357),
            .in2(_gnd_net_),
            .in3(N__9542),
            .lcout(\transmit_module.video_signal_controller.VGA_X_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3188 ),
            .carryout(\transmit_module.video_signal_controller.n3189 ),
            .clk(N__23482),
            .ce(),
            .sr(N__9822));
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_11_17_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_11_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i7_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__10294),
            .in2(_gnd_net_),
            .in3(N__9539),
            .lcout(\transmit_module.video_signal_controller.VGA_X_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3189 ),
            .carryout(\transmit_module.video_signal_controller.n3190 ),
            .clk(N__23482),
            .ce(),
            .sr(N__9822));
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_11_18_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_11_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i8_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__11846),
            .in2(_gnd_net_),
            .in3(N__9536),
            .lcout(\transmit_module.video_signal_controller.VGA_X_8 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\transmit_module.video_signal_controller.n3191 ),
            .clk(N__23647),
            .ce(),
            .sr(N__9823));
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_11_18_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_11_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i9_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__12407),
            .in2(_gnd_net_),
            .in3(N__9533),
            .lcout(\transmit_module.video_signal_controller.VGA_X_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3191 ),
            .carryout(\transmit_module.video_signal_controller.n3192 ),
            .clk(N__23647),
            .ce(),
            .sr(N__9823));
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_11_18_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_11_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i10_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__11548),
            .in2(_gnd_net_),
            .in3(N__9530),
            .lcout(\transmit_module.video_signal_controller.VGA_X_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3192 ),
            .carryout(\transmit_module.video_signal_controller.n3193 ),
            .clk(N__23647),
            .ce(),
            .sr(N__9823));
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_11_18_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_11_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i11_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__14277),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(\transmit_module.video_signal_controller.VGA_X_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23647),
            .ce(),
            .sr(N__9823));
    defparam \transmit_module.i1699_4_lut_LC_11_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1699_4_lut_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1699_4_lut_LC_11_19_0 .LUT_INIT=16'b1111011111110100;
    LogicCell40 \transmit_module.i1699_4_lut_LC_11_19_0  (
            .in0(N__20682),
            .in1(N__20264),
            .in2(N__20033),
            .in3(N__15146),
            .lcout(\transmit_module.n2073 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_12_3_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_12_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i9_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9590),
            .lcout(\tvp_video_buffer.BUFFER_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24099),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_12_7_1 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_12_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i10_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9566),
            .lcout(\tvp_video_buffer.BUFFER_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24114),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_12_7_7 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_12_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i2_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9578),
            .lcout(\tvp_video_buffer.BUFFER_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24114),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_12_9_6 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_12_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i6_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10412),
            .lcout(RX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24121),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_12_12_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_12_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_12_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i15_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14675),
            .lcout(\transmit_module.X_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23604),
            .ce(N__21475),
            .sr(N__21355));
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_12_12_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_12_12_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_12_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i13_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9554),
            .lcout(\transmit_module.X_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23604),
            .ce(N__21475),
            .sr(N__21355));
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_12_12_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_12_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i14_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9560),
            .lcout(\transmit_module.X_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23604),
            .ce(N__21475),
            .sr(N__21355));
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9638),
            .lcout(\transmit_module.Y_DELTA_PATTERN_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23532),
            .ce(N__9632),
            .sr(N__20017));
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_12_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_12_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_12_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i92_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9674),
            .lcout(\transmit_module.Y_DELTA_PATTERN_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23532),
            .ce(N__9632),
            .sr(N__20017));
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_12_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_12_13_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_12_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i93_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9680),
            .lcout(\transmit_module.Y_DELTA_PATTERN_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23532),
            .ce(N__9632),
            .sr(N__20017));
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_12_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_12_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i91_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9668),
            .lcout(\transmit_module.Y_DELTA_PATTERN_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23532),
            .ce(N__9632),
            .sr(N__20017));
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9650),
            .lcout(\transmit_module.Y_DELTA_PATTERN_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23532),
            .ce(N__9632),
            .sr(N__20017));
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9656),
            .lcout(\transmit_module.Y_DELTA_PATTERN_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23532),
            .ce(N__9632),
            .sr(N__20017));
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_12_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_12_13_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_12_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i90_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9644),
            .lcout(\transmit_module.Y_DELTA_PATTERN_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23532),
            .ce(N__9632),
            .sr(N__20017));
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_14_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__10975),
            .in2(_gnd_net_),
            .in3(N__9602),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_0 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\transmit_module.video_signal_controller.n3194 ),
            .clk(N__23667),
            .ce(N__9824),
            .sr(N__9782));
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_14_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__11013),
            .in2(_gnd_net_),
            .in3(N__9599),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3194 ),
            .carryout(\transmit_module.video_signal_controller.n3195 ),
            .clk(N__23667),
            .ce(N__9824),
            .sr(N__9782));
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_14_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__10962),
            .in2(_gnd_net_),
            .in3(N__9596),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3195 ),
            .carryout(\transmit_module.video_signal_controller.n3196 ),
            .clk(N__23667),
            .ce(N__9824),
            .sr(N__9782));
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_14_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__9893),
            .in2(_gnd_net_),
            .in3(N__9593),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3196 ),
            .carryout(\transmit_module.video_signal_controller.n3197 ),
            .clk(N__23667),
            .ce(N__9824),
            .sr(N__9782));
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_14_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__9860),
            .in2(_gnd_net_),
            .in3(N__9764),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3197 ),
            .carryout(\transmit_module.video_signal_controller.n3198 ),
            .clk(N__23667),
            .ce(N__9824),
            .sr(N__9782));
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_14_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__9988),
            .in2(_gnd_net_),
            .in3(N__9761),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3198 ),
            .carryout(\transmit_module.video_signal_controller.n3199 ),
            .clk(N__23667),
            .ce(N__9824),
            .sr(N__9782));
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_14_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__9964),
            .in2(_gnd_net_),
            .in3(N__9758),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3199 ),
            .carryout(\transmit_module.video_signal_controller.n3200 ),
            .clk(N__23667),
            .ce(N__9824),
            .sr(N__9782));
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_14_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__9755),
            .in2(_gnd_net_),
            .in3(N__9743),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3200 ),
            .carryout(\transmit_module.video_signal_controller.n3201 ),
            .clk(N__23667),
            .ce(N__9824),
            .sr(N__9782));
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_15_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__9740),
            .in2(_gnd_net_),
            .in3(N__9728),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_8 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\transmit_module.video_signal_controller.n3202 ),
            .clk(N__23656),
            .ce(N__9818),
            .sr(N__9778));
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_15_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__9938),
            .in2(_gnd_net_),
            .in3(N__9725),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3202 ),
            .carryout(\transmit_module.video_signal_controller.n3203 ),
            .clk(N__23656),
            .ce(N__9818),
            .sr(N__9778));
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_15_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__9698),
            .in2(_gnd_net_),
            .in3(N__9722),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3203 ),
            .carryout(\transmit_module.video_signal_controller.n3204 ),
            .clk(N__23656),
            .ce(N__9818),
            .sr(N__9778));
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_15_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__9716),
            .in2(_gnd_net_),
            .in3(N__9719),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23656),
            .ce(N__9818),
            .sr(N__9778));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_12_16_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_12_16_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__9715),
            .in2(_gnd_net_),
            .in3(N__9697),
            .lcout(\transmit_module.video_signal_controller.n3676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_16_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_16_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_LC_12_16_1  (
            .in0(N__9895),
            .in1(N__10964),
            .in2(_gnd_net_),
            .in3(N__11015),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3485_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_12_16_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_12_16_2 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_LC_12_16_2  (
            .in0(N__9989),
            .in1(N__9865),
            .in2(N__9968),
            .in3(N__9965),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3464_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_12_16_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_12_16_3 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_LC_12_16_3  (
            .in0(N__9944),
            .in1(N__9937),
            .in2(N__9920),
            .in3(N__9917),
            .lcout(\transmit_module.video_signal_controller.n3382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i6_3_lut_LC_12_16_4 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i6_3_lut_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i6_3_lut_LC_12_16_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i6_3_lut_LC_12_16_4  (
            .in0(N__20678),
            .in1(N__9905),
            .in2(_gnd_net_),
            .in3(N__13533),
            .lcout(\transmit_module.n111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_12_16_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_12_16_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_12_16_5  (
            .in0(N__10361),
            .in1(N__10331),
            .in2(_gnd_net_),
            .in3(N__10293),
            .lcout(\transmit_module.video_signal_controller.n2017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_12_16_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_12_16_7 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_12_16_7  (
            .in0(N__9896),
            .in1(N__9872),
            .in2(N__9866),
            .in3(N__9839),
            .lcout(\transmit_module.video_signal_controller.VGA_VISIBLE_N_588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_12_17_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_12_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__10376),
            .in2(_gnd_net_),
            .in3(N__10394),
            .lcout(\transmit_module.video_signal_controller.n3366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1738_4_lut_LC_12_17_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1738_4_lut_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1738_4_lut_LC_12_17_1 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \transmit_module.video_signal_controller.i1738_4_lut_LC_12_17_1  (
            .in0(N__11543),
            .in1(N__14269),
            .in2(N__10925),
            .in3(N__12406),
            .lcout(\transmit_module.video_signal_controller.n2050 ),
            .ltout(\transmit_module.video_signal_controller.n2050_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1163_2_lut_LC_12_17_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1163_2_lut_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1163_2_lut_LC_12_17_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1163_2_lut_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9785),
            .in3(N__13577),
            .lcout(\transmit_module.video_signal_controller.n2398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_17_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_17_3 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_17_3  (
            .in0(N__10377),
            .in1(N__10355),
            .in2(N__10400),
            .in3(N__10325),
            .lcout(\transmit_module.video_signal_controller.n55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_17_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_17_4 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_17_4  (
            .in0(N__12456),
            .in1(N__10395),
            .in2(N__12483),
            .in3(N__10275),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_12_17_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_12_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i3_4_lut_LC_12_17_5  (
            .in0(N__10378),
            .in1(N__10356),
            .in2(N__10334),
            .in3(N__10326),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3478_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_17_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_17_6 .LUT_INIT=16'b0000010101000100;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_17_6  (
            .in0(N__11544),
            .in1(N__10304),
            .in2(N__10298),
            .in3(N__10295),
            .lcout(\transmit_module.video_signal_controller.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1715_2_lut_3_lut_LC_12_17_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1715_2_lut_3_lut_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1715_2_lut_3_lut_LC_12_17_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \transmit_module.video_signal_controller.i1715_2_lut_3_lut_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__12455),
            .in2(N__10277),
            .in3(N__12473),
            .lcout(\transmit_module.video_signal_controller.n2958 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i13_LC_12_18_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i13_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i13_LC_12_18_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i13_LC_12_18_4  (
            .in0(N__10259),
            .in1(N__20253),
            .in2(_gnd_net_),
            .in3(N__13628),
            .lcout(TX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23571),
            .ce(N__10247),
            .sr(N__19935));
    defparam \transmit_module.i1653_4_lut_LC_12_19_7 .C_ON=1'b0;
    defparam \transmit_module.i1653_4_lut_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1653_4_lut_LC_12_19_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1653_4_lut_LC_12_19_7  (
            .in0(N__20226),
            .in1(N__12427),
            .in2(N__19995),
            .in3(N__12370),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_12_20_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_12_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i3_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16409),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23418),
            .ce(N__20773),
            .sr(N__20032));
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_13_5_6 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_13_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i0_LC_13_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10001),
            .lcout(RX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24102),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_13_6_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_13_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i3_LC_13_6_0  (
            .in0(N__10649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24105),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_13_6_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_13_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i11_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10634),
            .lcout(\tvp_video_buffer.BUFFER_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24105),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_13_7_1 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_13_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i7_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10628),
            .lcout(\tvp_video_buffer.BUFFER_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24110),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_13_7_3 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_13_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i1_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10616),
            .lcout(RX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24110),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_13_7_4 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_13_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i2_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10523),
            .lcout(RX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24110),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_13_8_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_13_8_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i15_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24115),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.X_246__i0_LC_13_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i0_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i0_LC_13_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i0_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__12566),
            .in2(_gnd_net_),
            .in3(N__10406),
            .lcout(\receive_module.rx_counter.X_0 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\receive_module.rx_counter.n3210 ),
            .clk(N__24118),
            .ce(),
            .sr(N__12502));
    defparam \receive_module.rx_counter.X_246__i1_LC_13_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i1_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i1_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i1_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__12578),
            .in2(_gnd_net_),
            .in3(N__10403),
            .lcout(\receive_module.rx_counter.X_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3210 ),
            .carryout(\receive_module.rx_counter.n3211 ),
            .clk(N__24118),
            .ce(),
            .sr(N__12502));
    defparam \receive_module.rx_counter.X_246__i2_LC_13_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i2_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i2_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i2_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__12554),
            .in2(_gnd_net_),
            .in3(N__10763),
            .lcout(\receive_module.rx_counter.X_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3211 ),
            .carryout(\receive_module.rx_counter.n3212 ),
            .clk(N__24118),
            .ce(),
            .sr(N__12502));
    defparam \receive_module.rx_counter.X_246__i3_LC_13_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i3_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i3_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i3_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__12989),
            .in2(_gnd_net_),
            .in3(N__10760),
            .lcout(\receive_module.rx_counter.X_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3212 ),
            .carryout(\receive_module.rx_counter.n3213 ),
            .clk(N__24118),
            .ce(),
            .sr(N__12502));
    defparam \receive_module.rx_counter.X_246__i4_LC_13_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i4_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i4_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i4_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__12536),
            .in2(_gnd_net_),
            .in3(N__10757),
            .lcout(\receive_module.rx_counter.X_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3213 ),
            .carryout(\receive_module.rx_counter.n3214 ),
            .clk(N__24118),
            .ce(),
            .sr(N__12502));
    defparam \receive_module.rx_counter.X_246__i5_LC_13_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i5_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i5_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i5_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__12971),
            .in2(_gnd_net_),
            .in3(N__10754),
            .lcout(\receive_module.rx_counter.X_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3214 ),
            .carryout(\receive_module.rx_counter.n3215 ),
            .clk(N__24118),
            .ce(),
            .sr(N__12502));
    defparam \receive_module.rx_counter.X_246__i6_LC_13_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i6_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i6_LC_13_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i6_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__12521),
            .in2(_gnd_net_),
            .in3(N__10751),
            .lcout(\receive_module.rx_counter.X_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3215 ),
            .carryout(\receive_module.rx_counter.n3216 ),
            .clk(N__24118),
            .ce(),
            .sr(N__12502));
    defparam \receive_module.rx_counter.X_246__i7_LC_13_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i7_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i7_LC_13_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i7_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__12953),
            .in2(_gnd_net_),
            .in3(N__10748),
            .lcout(\receive_module.rx_counter.X_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3216 ),
            .carryout(\receive_module.rx_counter.n3217 ),
            .clk(N__24118),
            .ce(),
            .sr(N__12502));
    defparam \receive_module.rx_counter.X_246__i8_LC_13_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_246__i8_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i8_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i8_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__12854),
            .in2(_gnd_net_),
            .in3(N__10745),
            .lcout(\receive_module.rx_counter.X_8 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\receive_module.rx_counter.n3218 ),
            .clk(N__24122),
            .ce(),
            .sr(N__12506));
    defparam \receive_module.rx_counter.X_246__i9_LC_13_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.X_246__i9_LC_13_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_246__i9_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_246__i9_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__12835),
            .in2(_gnd_net_),
            .in3(N__10742),
            .lcout(\receive_module.rx_counter.X_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24122),
            .ce(),
            .sr(N__12506));
    defparam \receive_module.rx_counter.Y__i0_LC_13_11_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i0_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i0_LC_13_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i0_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__13194),
            .in2(_gnd_net_),
            .in3(N__10739),
            .lcout(\receive_module.rx_counter.Y_0 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\receive_module.rx_counter.n3175 ),
            .clk(N__24127),
            .ce(N__12913),
            .sr(N__17554));
    defparam \receive_module.rx_counter.Y__i1_LC_13_11_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i1_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i1_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i1_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__13219),
            .in2(_gnd_net_),
            .in3(N__10787),
            .lcout(\receive_module.rx_counter.Y_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3175 ),
            .carryout(\receive_module.rx_counter.n3176 ),
            .clk(N__24127),
            .ce(N__12913),
            .sr(N__17554));
    defparam \receive_module.rx_counter.Y__i2_LC_13_11_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i2_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i2_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i2_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__13165),
            .in2(_gnd_net_),
            .in3(N__10784),
            .lcout(\receive_module.rx_counter.Y_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3176 ),
            .carryout(\receive_module.rx_counter.n3177 ),
            .clk(N__24127),
            .ce(N__12913),
            .sr(N__17554));
    defparam \receive_module.rx_counter.Y__i3_LC_13_11_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i3_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i3_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i3_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__13135),
            .in2(_gnd_net_),
            .in3(N__10781),
            .lcout(\receive_module.rx_counter.Y_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3177 ),
            .carryout(\receive_module.rx_counter.n3178 ),
            .clk(N__24127),
            .ce(N__12913),
            .sr(N__17554));
    defparam \receive_module.rx_counter.Y__i4_LC_13_11_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i4_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i4_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i4_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__13110),
            .in2(_gnd_net_),
            .in3(N__10778),
            .lcout(\receive_module.rx_counter.Y_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3178 ),
            .carryout(\receive_module.rx_counter.n3179 ),
            .clk(N__24127),
            .ce(N__12913),
            .sr(N__17554));
    defparam \receive_module.rx_counter.Y__i5_LC_13_11_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i5_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i5_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i5_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__12794),
            .in2(_gnd_net_),
            .in3(N__10775),
            .lcout(\receive_module.rx_counter.Y_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3179 ),
            .carryout(\receive_module.rx_counter.n3180 ),
            .clk(N__24127),
            .ce(N__12913),
            .sr(N__17554));
    defparam \receive_module.rx_counter.Y__i6_LC_13_11_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i6_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i6_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i6_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__12812),
            .in2(_gnd_net_),
            .in3(N__10772),
            .lcout(\receive_module.rx_counter.Y_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3180 ),
            .carryout(\receive_module.rx_counter.n3181 ),
            .clk(N__24127),
            .ce(N__12913),
            .sr(N__17554));
    defparam \receive_module.rx_counter.Y__i7_LC_13_11_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i7_LC_13_11_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i7_LC_13_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i7_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__13309),
            .in2(_gnd_net_),
            .in3(N__10769),
            .lcout(\receive_module.rx_counter.Y_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3181 ),
            .carryout(\receive_module.rx_counter.n3182 ),
            .clk(N__24127),
            .ce(N__12913),
            .sr(N__17554));
    defparam \receive_module.rx_counter.Y__i8_LC_13_12_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.Y__i8_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i8_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i8_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__13264),
            .in2(_gnd_net_),
            .in3(N__10766),
            .lcout(\receive_module.rx_counter.Y_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24131),
            .ce(N__12914),
            .sr(N__17541));
    defparam \receive_module.rx_counter.i2_2_lut_LC_13_13_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_LC_13_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__13115),
            .in2(_gnd_net_),
            .in3(N__13310),
            .lcout(\receive_module.rx_counter.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i6_4_lut_LC_13_13_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i6_4_lut_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i6_4_lut_LC_13_13_5 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \receive_module.rx_counter.i6_4_lut_LC_13_13_5  (
            .in0(N__13223),
            .in1(N__13139),
            .in2(N__13268),
            .in3(N__13169),
            .lcout(),
            .ltout(\receive_module.rx_counter.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.SYNC_46_LC_13_13_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.SYNC_46_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.SYNC_46_LC_13_13_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \receive_module.rx_counter.SYNC_46_LC_13_13_6  (
            .in0(N__10910),
            .in1(N__13199),
            .in2(N__10904),
            .in3(N__13283),
            .lcout(RX_TX_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24135),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i127_2_lut_4_lut_rep_23_LC_13_14_0 .C_ON=1'b0;
    defparam \transmit_module.i127_2_lut_4_lut_rep_23_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i127_2_lut_4_lut_rep_23_LC_13_14_0 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \transmit_module.i127_2_lut_4_lut_rep_23_LC_13_14_0  (
            .in0(N__10808),
            .in1(N__19692),
            .in2(N__11283),
            .in3(N__10861),
            .lcout(\transmit_module.n3682 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2193_3_lut_LC_13_14_1 .C_ON=1'b0;
    defparam \line_buffer.i2193_3_lut_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2193_3_lut_LC_13_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2193_3_lut_LC_13_14_1  (
            .in0(N__24714),
            .in1(N__10901),
            .in2(_gnd_net_),
            .in3(N__10886),
            .lcout(\line_buffer.n3530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.old_VGA_HS_40_LC_13_14_2 .C_ON=1'b0;
    defparam \transmit_module.old_VGA_HS_40_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.old_VGA_HS_40_LC_13_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.old_VGA_HS_40_LC_13_14_2  (
            .in0(N__10809),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.old_VGA_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23603),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i2_3_lut_rep_19_LC_13_14_3 .C_ON=1'b0;
    defparam \transmit_module.i2_3_lut_rep_19_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_3_lut_rep_19_LC_13_14_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \transmit_module.i2_3_lut_rep_19_LC_13_14_3  (
            .in0(N__10860),
            .in1(N__10807),
            .in2(_gnd_net_),
            .in3(N__11274),
            .lcout(\transmit_module.n3678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i8_3_lut_LC_13_14_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i8_3_lut_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i8_3_lut_LC_13_14_5 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \transmit_module.mux_12_i8_3_lut_LC_13_14_5  (
            .in0(N__20683),
            .in1(N__10847),
            .in2(N__13486),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_13_15_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_13_15_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \transmit_module.video_signal_controller.VGA_HS_66_LC_13_15_0  (
            .in0(N__11860),
            .in1(N__12416),
            .in2(N__14288),
            .in3(N__10838),
            .lcout(ADV_HSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23302),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i7_LC_13_15_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i7_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i7_LC_13_15_1 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i7_LC_13_15_1  (
            .in0(N__11252),
            .in1(N__20129),
            .in2(N__19721),
            .in3(N__11261),
            .lcout(\transmit_module.TX_ADDR_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23302),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i7_3_lut_LC_13_15_2 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i7_3_lut_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i7_3_lut_LC_13_15_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i7_3_lut_LC_13_15_2  (
            .in0(N__15141),
            .in1(N__15175),
            .in2(_gnd_net_),
            .in3(N__13499),
            .lcout(\transmit_module.n141 ),
            .ltout(\transmit_module.n141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1651_4_lut_LC_13_15_3 .C_ON=1'b0;
    defparam \transmit_module.i1651_4_lut_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1651_4_lut_LC_13_15_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1651_4_lut_LC_13_15_3  (
            .in0(N__19607),
            .in1(N__20127),
            .in2(N__11516),
            .in3(N__15199),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_15_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__14305),
            .in2(_gnd_net_),
            .in3(N__11801),
            .lcout(\transmit_module.VGA_VISIBLE_Y ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23302),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i8_3_lut_LC_13_15_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i8_3_lut_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i8_3_lut_LC_13_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i8_3_lut_LC_13_15_5  (
            .in0(N__15144),
            .in1(N__13482),
            .in2(_gnd_net_),
            .in3(N__13457),
            .lcout(\transmit_module.n140 ),
            .ltout(\transmit_module.n140_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1652_4_lut_LC_13_15_6 .C_ON=1'b0;
    defparam \transmit_module.i1652_4_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1652_4_lut_LC_13_15_6 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.i1652_4_lut_LC_13_15_6  (
            .in0(N__20128),
            .in1(N__19608),
            .in2(N__11255),
            .in3(N__11251),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_13_15_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_13_15_7 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VS_67_LC_13_15_7  (
            .in0(N__11014),
            .in1(N__10988),
            .in2(N__10979),
            .in3(N__10963),
            .lcout(ADV_VSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23302),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1732_4_lut_LC_13_16_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1732_4_lut_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1732_4_lut_LC_13_16_0 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \transmit_module.video_signal_controller.i1732_4_lut_LC_13_16_0  (
            .in0(N__11819),
            .in1(N__11856),
            .in2(N__10937),
            .in3(N__11872),
            .lcout(\transmit_module.video_signal_controller.n2975 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i2_3_lut_LC_13_16_3 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i2_3_lut_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i2_3_lut_LC_13_16_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i2_3_lut_LC_13_16_3  (
            .in0(N__14503),
            .in1(N__15126),
            .in2(_gnd_net_),
            .in3(N__13322),
            .lcout(\transmit_module.n146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i4_LC_13_16_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i4_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i4_LC_13_16_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i4_LC_13_16_4  (
            .in0(N__20180),
            .in1(N__13616),
            .in2(N__19837),
            .in3(N__11789),
            .lcout(\transmit_module.TX_ADDR_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23488),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i5_LC_13_16_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i5_LC_13_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i5_LC_13_16_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i5_LC_13_16_5  (
            .in0(N__20193),
            .in1(N__12104),
            .in2(N__19722),
            .in3(N__12113),
            .lcout(\transmit_module.TX_ADDR_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23488),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i6_3_lut_LC_13_16_6 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i6_3_lut_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i6_3_lut_LC_13_16_6 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \transmit_module.mux_14_i6_3_lut_LC_13_16_6  (
            .in0(N__15127),
            .in1(N__13534),
            .in2(N__13511),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n142 ),
            .ltout(\transmit_module.n142_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1650_4_lut_LC_13_16_7 .C_ON=1'b0;
    defparam \transmit_module.i1650_4_lut_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1650_4_lut_LC_13_16_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1650_4_lut_LC_13_16_7  (
            .in0(N__19612),
            .in1(N__20179),
            .in2(N__12107),
            .in3(N__12103),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1764_4_lut_LC_13_17_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1764_4_lut_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1764_4_lut_LC_13_17_0 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \transmit_module.video_signal_controller.i1764_4_lut_LC_13_17_0  (
            .in0(N__12434),
            .in1(N__11873),
            .in2(N__11861),
            .in3(N__11818),
            .lcout(\transmit_module.video_signal_controller.n3007 ),
            .ltout(\transmit_module.video_signal_controller.n3007_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_13_17_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_13_17_1 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_13_17_1  (
            .in0(N__11555),
            .in1(N__12377),
            .in2(N__11804),
            .in3(N__11800),
            .lcout(\transmit_module.video_signal_controller.n7_adj_624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i8_LC_13_17_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i8_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i8_LC_13_17_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i8_LC_13_17_2  (
            .in0(N__20195),
            .in1(N__12428),
            .in2(N__19866),
            .in3(N__12371),
            .lcout(\transmit_module.TX_ADDR_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23405),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i5_3_lut_LC_13_17_3 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i5_3_lut_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i5_3_lut_LC_13_17_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \transmit_module.mux_14_i5_3_lut_LC_13_17_3  (
            .in0(N__15119),
            .in1(_gnd_net_),
            .in2(N__13553),
            .in3(N__20806),
            .lcout(\transmit_module.n143 ),
            .ltout(\transmit_module.n143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1649_4_lut_LC_13_17_4 .C_ON=1'b0;
    defparam \transmit_module.i1649_4_lut_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1649_4_lut_LC_13_17_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1649_4_lut_LC_13_17_4  (
            .in0(N__19723),
            .in1(N__20181),
            .in2(N__11783),
            .in3(N__13615),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1774_3_lut_LC_13_17_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1774_3_lut_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1774_3_lut_LC_13_17_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \transmit_module.video_signal_controller.i1774_3_lut_LC_13_17_5  (
            .in0(N__11554),
            .in1(N__12415),
            .in2(_gnd_net_),
            .in3(N__11522),
            .lcout(\transmit_module.video_signal_controller.n3017 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i509_2_lut_rep_20_LC_13_17_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i509_2_lut_rep_20_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i509_2_lut_rep_20_LC_13_17_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i509_2_lut_rep_20_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__12484),
            .in2(_gnd_net_),
            .in3(N__12457),
            .lcout(\transmit_module.video_signal_controller.n3679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_18_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_18_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_12_i9_3_lut_LC_13_18_5  (
            .in0(N__14513),
            .in1(N__20661),
            .in2(_gnd_net_),
            .in3(N__14535),
            .lcout(\transmit_module.n108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_2_lut_LC_13_18_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_2_lut_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_2_lut_LC_13_18_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i2_2_lut_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__14273),
            .in2(_gnd_net_),
            .in3(N__12408),
            .lcout(\transmit_module.video_signal_controller.n6_adj_623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i9_3_lut_LC_13_18_7 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i9_3_lut_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i9_3_lut_LC_13_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i9_3_lut_LC_13_18_7  (
            .in0(N__15115),
            .in1(N__14534),
            .in2(_gnd_net_),
            .in3(N__13448),
            .lcout(\transmit_module.n139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i10_3_lut_LC_13_19_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i10_3_lut_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i10_3_lut_LC_13_19_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \transmit_module.mux_14_i10_3_lut_LC_13_19_5  (
            .in0(N__14211),
            .in1(_gnd_net_),
            .in2(N__15143),
            .in3(N__13436),
            .lcout(\transmit_module.n138 ),
            .ltout(\transmit_module.n138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1654_4_lut_LC_13_19_6 .C_ON=1'b0;
    defparam \transmit_module.i1654_4_lut_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1654_4_lut_LC_13_19_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1654_4_lut_LC_13_19_6  (
            .in0(N__19727),
            .in1(N__20194),
            .in2(N__12359),
            .in3(N__14176),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_13_20_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_13_20_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_LC_13_20_2  (
            .in0(N__22306),
            .in1(N__12140),
            .in2(N__23919),
            .in3(N__12131),
            .lcout(\line_buffer.n3620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1144_1_lut_LC_13_20_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1144_1_lut_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1144_1_lut_LC_13_20_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \transmit_module.video_signal_controller.i1144_1_lut_LC_13_20_3  (
            .in0(N__15142),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n2388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i7_LC_13_21_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i7_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i7_LC_13_21_5 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \line_buffer.dout_i7_LC_13_21_5  (
            .in0(N__12743),
            .in1(N__12650),
            .in2(N__23933),
            .in3(N__12119),
            .lcout(TX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23228),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2197_3_lut_LC_13_22_2 .C_ON=1'b0;
    defparam \line_buffer.i2197_3_lut_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2197_3_lut_LC_13_22_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2197_3_lut_LC_13_22_2  (
            .in0(N__12776),
            .in1(N__12761),
            .in2(_gnd_net_),
            .in3(N__24780),
            .lcout(\line_buffer.n3534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i8_LC_13_24_2 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i8_LC_13_24_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i8_LC_13_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i8_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12737),
            .lcout(ADV_B_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23257),
            .ce(),
            .sr(N__22670));
    defparam \line_buffer.i2196_3_lut_LC_13_25_6 .C_ON=1'b0;
    defparam \line_buffer.i2196_3_lut_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2196_3_lut_LC_13_25_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2196_3_lut_LC_13_25_6  (
            .in0(N__12677),
            .in1(N__12665),
            .in2(_gnd_net_),
            .in3(N__24798),
            .lcout(\line_buffer.n3533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_14_9_2 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_14_9_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_LC_14_9_2  (
            .in0(N__14927),
            .in1(N__14828),
            .in2(N__14882),
            .in3(N__18682),
            .lcout(\line_buffer.n542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_adj_23_LC_14_9_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_adj_23_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_adj_23_LC_14_9_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_adj_23_LC_14_9_3  (
            .in0(N__12577),
            .in1(N__12565),
            .in2(_gnd_net_),
            .in3(N__12553),
            .lcout(\receive_module.rx_counter.n3225 ),
            .ltout(\receive_module.rx_counter.n3225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i3_4_lut_LC_14_9_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i3_4_lut_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i3_4_lut_LC_14_9_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \receive_module.rx_counter.i3_4_lut_LC_14_9_4  (
            .in0(N__12534),
            .in1(N__12988),
            .in2(N__12542),
            .in3(N__12969),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3458_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_4_lut_LC_14_9_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_4_lut_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_4_lut_LC_14_9_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \receive_module.rx_counter.i1_4_lut_LC_14_9_5  (
            .in0(N__12520),
            .in1(N__12951),
            .in2(N__12539),
            .in3(N__12852),
            .lcout(\receive_module.rx_counter.n39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_9_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_9_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_9_6  (
            .in0(N__12535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12519),
            .lcout(\receive_module.rx_counter.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_1_lut_LC_14_9_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_1_lut_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_1_lut_LC_14_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \receive_module.rx_counter.i5_1_lut_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14335),
            .lcout(\receive_module.rx_counter.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_2_lut_adj_25_LC_14_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_adj_25_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_adj_25_LC_14_10_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_adj_25_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__12987),
            .in2(_gnd_net_),
            .in3(N__12970),
            .lcout(),
            .ltout(\receive_module.rx_counter.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2092_4_lut_LC_14_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2092_4_lut_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2092_4_lut_LC_14_10_2 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \receive_module.rx_counter.i2092_4_lut_LC_14_10_2  (
            .in0(N__12952),
            .in1(N__12935),
            .in2(N__12929),
            .in3(N__12926),
            .lcout(\receive_module.rx_counter.n3429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_HS_51_LC_14_11_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_HS_51_LC_14_11_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_HS_51_LC_14_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receive_module.rx_counter.old_HS_51_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14344),
            .lcout(\receive_module.rx_counter.old_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24123),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i252_3_lut_LC_14_11_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i252_3_lut_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i252_3_lut_LC_14_11_3 .LUT_INIT=16'b0101111101010101;
    LogicCell40 \receive_module.rx_counter.i252_3_lut_LC_14_11_3  (
            .in0(N__18862),
            .in1(_gnd_net_),
            .in2(N__14345),
            .in3(N__12920),
            .lcout(\receive_module.rx_counter.n2081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_14_11_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_14_11_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_14_11_4  (
            .in0(N__14867),
            .in1(N__18662),
            .in2(N__14827),
            .in3(N__14923),
            .lcout(\line_buffer.n573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i609_2_lut_rep_21_LC_14_11_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i609_2_lut_rep_21_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i609_2_lut_rep_21_LC_14_11_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i609_2_lut_rep_21_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__12811),
            .in2(_gnd_net_),
            .in3(N__12792),
            .lcout(\receive_module.rx_counter.n3680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i58_4_lut_LC_14_11_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i58_4_lut_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i58_4_lut_LC_14_11_6 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \receive_module.rx_counter.i58_4_lut_LC_14_11_6  (
            .in0(N__12860),
            .in1(N__12853),
            .in2(N__12836),
            .in3(N__12821),
            .lcout(\receive_module.rx_counter.n54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_12_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_12_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_12_0  (
            .in0(N__13304),
            .in1(N__12810),
            .in2(_gnd_net_),
            .in3(N__12793),
            .lcout(),
            .ltout(\receive_module.rx_counter.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i3_4_lut_adj_21_LC_14_12_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i3_4_lut_adj_21_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i3_4_lut_adj_21_LC_14_12_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \receive_module.rx_counter.i3_4_lut_adj_21_LC_14_12_1  (
            .in0(N__13262),
            .in1(N__13088),
            .in2(N__13313),
            .in3(N__13145),
            .lcout(\receive_module.rx_counter.n3481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_LC_14_12_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_LC_14_12_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_LC_14_12_2  (
            .in0(N__13218),
            .in1(N__13133),
            .in2(N__13198),
            .in3(N__13163),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_4_lut_adj_22_LC_14_12_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_4_lut_adj_22_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_4_lut_adj_22_LC_14_12_3 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \receive_module.rx_counter.i1_4_lut_adj_22_LC_14_12_3  (
            .in0(N__13114),
            .in1(N__13305),
            .in2(N__13286),
            .in3(N__13279),
            .lcout(),
            .ltout(\receive_module.rx_counter.n4_adj_612_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_14_12_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_14_12_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_14_12_4 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \receive_module.rx_counter.O_VISIBLE_53_LC_14_12_4  (
            .in0(N__13263),
            .in1(N__13238),
            .in2(N__13232),
            .in3(N__13229),
            .lcout(DEBUG_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24128),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_LC_14_12_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_LC_14_12_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_LC_14_12_6  (
            .in0(N__13217),
            .in1(N__13193),
            .in2(_gnd_net_),
            .in3(N__13164),
            .lcout(\receive_module.rx_counter.n3453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_27_LC_14_12_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_27_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_27_LC_14_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_27_LC_14_12_7  (
            .in0(N__13134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13109),
            .lcout(\receive_module.rx_counter.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.BUFFER_0__i1_LC_14_13_2 .C_ON=1'b0;
    defparam \sync_buffer.BUFFER_0__i1_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.BUFFER_0__i1_LC_14_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \sync_buffer.BUFFER_0__i1_LC_14_13_2  (
            .in0(N__13082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sync_buffer.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23531),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_14_13_3 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_14_13_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_14_13_3  (
            .in0(N__14922),
            .in1(N__14879),
            .in2(N__14821),
            .in3(N__18661),
            .lcout(\line_buffer.n477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_14_13_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_14_13_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_14_13_4  (
            .in0(N__14880),
            .in1(N__18659),
            .in2(N__14825),
            .in3(N__14920),
            .lcout(\line_buffer.n541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_14_13_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_14_13_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_14_13_5  (
            .in0(N__14921),
            .in1(N__14881),
            .in2(N__14822),
            .in3(N__18660),
            .lcout(\line_buffer.n605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i2_3_lut_LC_14_14_0 .C_ON=1'b0;
    defparam \transmit_module.i2_3_lut_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_3_lut_LC_14_14_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.i2_3_lut_LC_14_14_0  (
            .in0(N__20162),
            .in1(N__19694),
            .in2(_gnd_net_),
            .in3(N__15145),
            .lcout(\transmit_module.n2087 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2215_3_lut_LC_14_14_1 .C_ON=1'b0;
    defparam \line_buffer.i2215_3_lut_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2215_3_lut_LC_14_14_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2215_3_lut_LC_14_14_1  (
            .in0(N__13370),
            .in1(N__13352),
            .in2(_gnd_net_),
            .in3(N__24715),
            .lcout(\line_buffer.n3552 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.BUFFER_0__i2_LC_14_14_2 .C_ON=1'b0;
    defparam \sync_buffer.BUFFER_0__i2_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.BUFFER_0__i2_LC_14_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.BUFFER_0__i2_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13337),
            .lcout(\sync_buffer.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23666),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_14_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_14_5 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i0_LC_14_14_5  (
            .in0(N__14144),
            .in1(N__20163),
            .in2(N__19836),
            .in3(N__14129),
            .lcout(\transmit_module.TX_ADDR_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23666),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_14_6 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_14_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i7_3_lut_LC_14_14_6  (
            .in0(N__20676),
            .in1(N__13331),
            .in2(_gnd_net_),
            .in3(N__15173),
            .lcout(\transmit_module.n110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1_3_lut_LC_14_14_7 .C_ON=1'b0;
    defparam \transmit_module.i1_3_lut_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1_3_lut_LC_14_14_7 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \transmit_module.i1_3_lut_LC_14_14_7  (
            .in0(N__19693),
            .in1(N__20677),
            .in2(_gnd_net_),
            .in3(N__20161),
            .lcout(\transmit_module.n2313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_2_lut_LC_14_15_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_2_lut_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_2_lut_LC_14_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_2_lut_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__14450),
            .in2(N__14671),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n132 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\transmit_module.n3162 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_3_lut_LC_14_15_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_3_lut_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_3_lut_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_3_lut_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__14492),
            .in2(_gnd_net_),
            .in3(N__13316),
            .lcout(\transmit_module.n131 ),
            .ltout(),
            .carryin(\transmit_module.n3162 ),
            .carryout(\transmit_module.n3163 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_4_lut_LC_14_15_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_4_lut_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_4_lut_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_4_lut_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__20573),
            .in2(_gnd_net_),
            .in3(N__13559),
            .lcout(\transmit_module.n130 ),
            .ltout(),
            .carryin(\transmit_module.n3163 ),
            .carryout(\transmit_module.n3164 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_5_lut_LC_14_15_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_5_lut_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_5_lut_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_5_lut_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16404),
            .in3(N__13556),
            .lcout(\transmit_module.n129 ),
            .ltout(),
            .carryin(\transmit_module.n3164 ),
            .carryout(\transmit_module.n3165 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_6_lut_LC_14_15_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_6_lut_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_6_lut_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_6_lut_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__20804),
            .in2(_gnd_net_),
            .in3(N__13541),
            .lcout(\transmit_module.n128 ),
            .ltout(),
            .carryin(\transmit_module.n3165 ),
            .carryout(\transmit_module.n3166 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_7_lut_LC_14_15_5 .C_ON=1'b1;
    defparam \transmit_module.add_13_7_lut_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_7_lut_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_7_lut_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__13532),
            .in2(_gnd_net_),
            .in3(N__13502),
            .lcout(\transmit_module.n127 ),
            .ltout(),
            .carryin(\transmit_module.n3166 ),
            .carryout(\transmit_module.n3167 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_8_lut_LC_14_15_6 .C_ON=1'b1;
    defparam \transmit_module.add_13_8_lut_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_8_lut_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_8_lut_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15174),
            .in3(N__13493),
            .lcout(\transmit_module.n126 ),
            .ltout(),
            .carryin(\transmit_module.n3167 ),
            .carryout(\transmit_module.n3168 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_9_lut_LC_14_15_7 .C_ON=1'b1;
    defparam \transmit_module.add_13_9_lut_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_9_lut_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_9_lut_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__13478),
            .in2(_gnd_net_),
            .in3(N__13451),
            .lcout(\transmit_module.n125 ),
            .ltout(),
            .carryin(\transmit_module.n3168 ),
            .carryout(\transmit_module.n3169 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_10_lut_LC_14_16_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_10_lut_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_10_lut_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_10_lut_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14539),
            .in3(N__13439),
            .lcout(\transmit_module.n124 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\transmit_module.n3170 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_11_lut_LC_14_16_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_11_lut_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_11_lut_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_11_lut_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14210),
            .in3(N__13424),
            .lcout(\transmit_module.n123 ),
            .ltout(),
            .carryin(\transmit_module.n3170 ),
            .carryout(\transmit_module.n3171 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_12_lut_LC_14_16_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_12_lut_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_12_lut_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_12_lut_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14578),
            .in3(N__13421),
            .lcout(\transmit_module.n122 ),
            .ltout(),
            .carryin(\transmit_module.n3171 ),
            .carryout(\transmit_module.n3172 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_13_lut_LC_14_16_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_13_lut_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_13_lut_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_13_lut_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__24732),
            .in2(_gnd_net_),
            .in3(N__13646),
            .lcout(\transmit_module.n121 ),
            .ltout(),
            .carryin(\transmit_module.n3172 ),
            .carryout(\transmit_module.n3173 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_14_lut_LC_14_16_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_14_lut_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_14_lut_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_14_lut_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__22305),
            .in2(_gnd_net_),
            .in3(N__13634),
            .lcout(\transmit_module.n120 ),
            .ltout(),
            .carryin(\transmit_module.n3173 ),
            .carryout(\transmit_module.n3174 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_15_lut_LC_14_16_5 .C_ON=1'b0;
    defparam \transmit_module.add_13_15_lut_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_15_lut_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_15_lut_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__23917),
            .in2(_gnd_net_),
            .in3(N__13631),
            .lcout(\transmit_module.n119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_16_6 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_16_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i5_3_lut_LC_14_16_6  (
            .in0(N__20672),
            .in1(N__20783),
            .in2(_gnd_net_),
            .in3(N__20805),
            .lcout(\transmit_module.n112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_16_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_16_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i1_LC_14_16_7  (
            .in0(N__20261),
            .in1(N__14164),
            .in2(N__19838),
            .in3(N__13600),
            .lcout(\transmit_module.TX_ADDR_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23560),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.WIRE_OUT_0__9_LC_14_17_1 .C_ON=1'b0;
    defparam \sync_buffer.WIRE_OUT_0__9_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.WIRE_OUT_0__9_LC_14_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.WIRE_OUT_0__9_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13586),
            .lcout(RX_TX_SYNC_BUFF),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23376),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_17_3 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_17_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i11_3_lut_LC_14_17_3  (
            .in0(N__15096),
            .in1(N__14573),
            .in2(_gnd_net_),
            .in3(N__13568),
            .lcout(\transmit_module.n137 ),
            .ltout(\transmit_module.n137_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_17_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_17_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \transmit_module.BRAM_ADDR__i10_LC_14_17_4  (
            .in0(N__13895),
            .in1(N__19739),
            .in2(N__13562),
            .in3(N__20262),
            .lcout(\transmit_module.TX_ADDR_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23376),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_17_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_17_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_17_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i9_LC_14_17_5  (
            .in0(N__20263),
            .in1(N__14180),
            .in2(N__19875),
            .in3(N__14324),
            .lcout(\transmit_module.TX_ADDR_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23376),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_17_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_17_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_17_7  (
            .in0(N__14312),
            .in1(N__14294),
            .in2(N__14287),
            .in3(N__14240),
            .lcout(\transmit_module.VGA_VISIBLE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23376),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_18_0 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \transmit_module.mux_14_i1_3_lut_LC_14_18_0  (
            .in0(N__15097),
            .in1(N__14234),
            .in2(_gnd_net_),
            .in3(N__14460),
            .lcout(\transmit_module.n147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i11_3_lut_LC_14_18_6 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i11_3_lut_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i11_3_lut_LC_14_18_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i11_3_lut_LC_14_18_6  (
            .in0(N__20625),
            .in1(N__14549),
            .in2(_gnd_net_),
            .in3(N__14574),
            .lcout(\transmit_module.n106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_19_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_19_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i10_3_lut_LC_14_19_1  (
            .in0(N__20671),
            .in1(N__14225),
            .in2(_gnd_net_),
            .in3(N__14212),
            .lcout(\transmit_module.n107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_19_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_19_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i2_3_lut_LC_14_19_2  (
            .in0(N__20647),
            .in1(N__14471),
            .in2(_gnd_net_),
            .in3(N__14502),
            .lcout(\transmit_module.n115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_19_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_19_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_12_i1_3_lut_LC_14_19_5  (
            .in0(N__14435),
            .in1(N__20648),
            .in2(_gnd_net_),
            .in3(N__14461),
            .lcout(\transmit_module.n116 ),
            .ltout(\transmit_module.n116_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1640_4_lut_LC_14_19_6 .C_ON=1'b0;
    defparam \transmit_module.i1640_4_lut_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1640_4_lut_LC_14_19_6 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \transmit_module.i1640_4_lut_LC_14_19_6  (
            .in0(N__19873),
            .in1(N__20236),
            .in2(N__14132),
            .in3(N__14125),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1655_4_lut_LC_14_19_7 .C_ON=1'b0;
    defparam \transmit_module.i1655_4_lut_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1655_4_lut_LC_14_19_7 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \transmit_module.i1655_4_lut_LC_14_19_7  (
            .in0(N__13894),
            .in1(N__19874),
            .in2(N__20260),
            .in3(N__13883),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_20_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_20_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14579),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23417),
            .ce(N__20748),
            .sr(N__20058));
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_20_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_20_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14540),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23417),
            .ce(N__20748),
            .sr(N__20058));
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_20_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_20_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14504),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23417),
            .ce(N__20748),
            .sr(N__20058));
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_20_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_20_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14465),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23417),
            .ce(N__20748),
            .sr(N__20058));
    defparam \tvp_vs_buffer.BUFFER_0__i1_LC_15_6_3 .C_ON=1'b0;
    defparam \tvp_vs_buffer.BUFFER_0__i1_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \tvp_vs_buffer.BUFFER_0__i1_LC_15_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_vs_buffer.BUFFER_0__i1_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14413),
            .lcout(\tvp_vs_buffer.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24100),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_15_8_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_15_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i5_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14389),
            .lcout(\tvp_video_buffer.BUFFER_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24106),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_vs_buffer.BUFFER_0__i2_LC_15_8_6 .C_ON=1'b0;
    defparam \tvp_vs_buffer.BUFFER_0__i2_LC_15_8_6 .SEQ_MODE=4'b1000;
    defparam \tvp_vs_buffer.BUFFER_0__i2_LC_15_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_vs_buffer.BUFFER_0__i2_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14360),
            .lcout(\tvp_vs_buffer.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24106),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_15_9_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_15_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i13_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14351),
            .lcout(\tvp_video_buffer.BUFFER_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24111),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_15_9_4 .C_ON=1'b0;
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_15_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_hs_buffer.WIRE_OUT_0__9_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20849),
            .lcout(TVP_HSYNC_buff),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24111),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_15_10_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_15_10_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_15_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i10_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14615),
            .lcout(\transmit_module.X_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23551),
            .ce(N__21476),
            .sr(N__21362));
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_15_10_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_15_10_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_15_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i9_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14627),
            .lcout(\transmit_module.X_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23551),
            .ce(N__21476),
            .sr(N__21362));
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_15_10_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_15_10_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_15_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i8_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14621),
            .lcout(\transmit_module.X_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23551),
            .ce(N__21476),
            .sr(N__21362));
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_15_10_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_15_10_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_15_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i11_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14597),
            .lcout(\transmit_module.X_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23551),
            .ce(N__21476),
            .sr(N__21362));
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_15_10_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_15_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i12_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14609),
            .lcout(\transmit_module.X_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23551),
            .ce(N__21476),
            .sr(N__21362));
    defparam \receive_module.add_12_2_lut_LC_15_11_0 .C_ON=1'b1;
    defparam \receive_module.add_12_2_lut_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_2_lut_LC_15_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_2_lut_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__18099),
            .in2(_gnd_net_),
            .in3(N__14591),
            .lcout(\receive_module.n137 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\receive_module.n3149 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_3_lut_LC_15_11_1 .C_ON=1'b1;
    defparam \receive_module.add_12_3_lut_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_3_lut_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_3_lut_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__15540),
            .in2(_gnd_net_),
            .in3(N__14588),
            .lcout(\receive_module.n136 ),
            .ltout(),
            .carryin(\receive_module.n3149 ),
            .carryout(\receive_module.n3150 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_4_lut_LC_15_11_2 .C_ON=1'b1;
    defparam \receive_module.add_12_4_lut_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_4_lut_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_4_lut_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__15288),
            .in2(_gnd_net_),
            .in3(N__14585),
            .lcout(\receive_module.n135 ),
            .ltout(),
            .carryin(\receive_module.n3150 ),
            .carryout(\receive_module.n3151 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_5_lut_LC_15_11_3 .C_ON=1'b1;
    defparam \receive_module.add_12_5_lut_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_5_lut_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_5_lut_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__17862),
            .in2(_gnd_net_),
            .in3(N__14582),
            .lcout(\receive_module.n134 ),
            .ltout(),
            .carryin(\receive_module.n3151 ),
            .carryout(\receive_module.n3152 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_6_lut_LC_15_11_4 .C_ON=1'b1;
    defparam \receive_module.add_12_6_lut_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_6_lut_LC_15_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_6_lut_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__17244),
            .in2(_gnd_net_),
            .in3(N__14654),
            .lcout(\receive_module.n133 ),
            .ltout(),
            .carryin(\receive_module.n3152 ),
            .carryout(\receive_module.n3153 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_7_lut_LC_15_11_5 .C_ON=1'b1;
    defparam \receive_module.add_12_7_lut_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_7_lut_LC_15_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_7_lut_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__16992),
            .in2(_gnd_net_),
            .in3(N__14651),
            .lcout(\receive_module.n132 ),
            .ltout(),
            .carryin(\receive_module.n3153 ),
            .carryout(\receive_module.n3154 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_8_lut_LC_15_11_6 .C_ON=1'b1;
    defparam \receive_module.add_12_8_lut_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_8_lut_LC_15_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_8_lut_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__16725),
            .in2(_gnd_net_),
            .in3(N__14648),
            .lcout(\receive_module.n131 ),
            .ltout(),
            .carryin(\receive_module.n3154 ),
            .carryout(\receive_module.n3155 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_9_lut_LC_15_11_7 .C_ON=1'b1;
    defparam \receive_module.add_12_9_lut_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_9_lut_LC_15_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_9_lut_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__16464),
            .in2(_gnd_net_),
            .in3(N__14645),
            .lcout(\receive_module.n130 ),
            .ltout(),
            .carryin(\receive_module.n3155 ),
            .carryout(\receive_module.n3156 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_10_lut_LC_15_12_0 .C_ON=1'b1;
    defparam \receive_module.add_12_10_lut_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_10_lut_LC_15_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_10_lut_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__15828),
            .in2(_gnd_net_),
            .in3(N__14642),
            .lcout(\receive_module.n129 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\receive_module.n3157 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_11_lut_LC_15_12_1 .C_ON=1'b1;
    defparam \receive_module.add_12_11_lut_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_11_lut_LC_15_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_11_lut_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__16173),
            .in2(_gnd_net_),
            .in3(N__14639),
            .lcout(\receive_module.n128 ),
            .ltout(),
            .carryin(\receive_module.n3157 ),
            .carryout(\receive_module.n3158 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_12_lut_LC_15_12_2 .C_ON=1'b1;
    defparam \receive_module.add_12_12_lut_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_12_lut_LC_15_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_12_lut_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__17625),
            .in2(_gnd_net_),
            .in3(N__14636),
            .lcout(\receive_module.n127 ),
            .ltout(),
            .carryin(\receive_module.n3158 ),
            .carryout(\receive_module.n3159 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i11_LC_15_12_3 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i11_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i11_LC_15_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i11_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__14916),
            .in2(_gnd_net_),
            .in3(N__14633),
            .lcout(RX_ADDR_11),
            .ltout(),
            .carryin(\receive_module.n3159 ),
            .carryout(\receive_module.n3160 ),
            .clk(N__24124),
            .ce(N__14939),
            .sr(N__17513));
    defparam \receive_module.BRAM_ADDR__i12_LC_15_12_4 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i12_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i12_LC_15_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i12_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__14868),
            .in2(_gnd_net_),
            .in3(N__14630),
            .lcout(RX_ADDR_12),
            .ltout(),
            .carryin(\receive_module.n3160 ),
            .carryout(\receive_module.n3161 ),
            .clk(N__24124),
            .ce(N__14939),
            .sr(N__17513));
    defparam \receive_module.BRAM_ADDR__i13_LC_15_12_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i13_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i13_LC_15_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i13_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__14817),
            .in2(_gnd_net_),
            .in3(N__15038),
            .lcout(RX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24124),
            .ce(N__14939),
            .sr(N__17513));
    defparam \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_13_1 .C_ON=1'b0;
    defparam \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14681),
            .lcout(TVP_VSYNC_buff),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24129),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_15_13_2 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_15_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_15_13_2  (
            .in0(N__14918),
            .in1(N__14865),
            .in2(N__14823),
            .in3(N__18663),
            .lcout(\line_buffer.n606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_15_13_3 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_15_13_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_15_13_3  (
            .in0(N__18665),
            .in1(N__14864),
            .in2(N__14826),
            .in3(N__14917),
            .lcout(\line_buffer.n476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18843),
            .lcout(\receive_module.n3677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i249_2_lut_rep_15_2_lut_LC_15_13_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i249_2_lut_rep_15_2_lut_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i249_2_lut_rep_15_2_lut_LC_15_13_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \receive_module.rx_counter.i249_2_lut_rep_15_2_lut_LC_15_13_5  (
            .in0(N__18844),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18669),
            .lcout(\receive_module.n3674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_15_13_6 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_15_13_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_15_13_6  (
            .in0(N__14919),
            .in1(N__14866),
            .in2(N__14824),
            .in3(N__18664),
            .lcout(\line_buffer.n574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_vs_buffer.BUFFER_0__i3_LC_15_13_7 .C_ON=1'b0;
    defparam \tvp_vs_buffer.BUFFER_0__i3_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \tvp_vs_buffer.BUFFER_0__i3_LC_15_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_vs_buffer.BUFFER_0__i3_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14693),
            .lcout(\tvp_vs_buffer.BUFFER_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24129),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15245),
            .lcout(\transmit_module.X_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23409),
            .ce(N__21464),
            .sr(N__21327));
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15230),
            .lcout(\transmit_module.X_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23409),
            .ce(N__21464),
            .sr(N__21327));
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15239),
            .lcout(\transmit_module.X_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23409),
            .ce(N__21464),
            .sr(N__21327));
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15224),
            .lcout(\transmit_module.X_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23409),
            .ce(N__21464),
            .sr(N__21327));
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_15_14_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_15_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_15_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i3_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15212),
            .lcout(\transmit_module.X_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23409),
            .ce(N__21464),
            .sr(N__21327));
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_15_14_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_15_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_15_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i6_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15218),
            .lcout(\transmit_module.X_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23409),
            .ce(N__21464),
            .sr(N__21327));
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_15_14_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_15_14_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_15_14_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i4_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__21485),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23409),
            .ce(N__21464),
            .sr(N__21327));
    defparam \transmit_module.mux_14_i4_3_lut_LC_15_15_1 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i4_3_lut_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i4_3_lut_LC_15_15_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.mux_14_i4_3_lut_LC_15_15_1  (
            .in0(N__15206),
            .in1(N__15140),
            .in2(_gnd_net_),
            .in3(N__16397),
            .lcout(\transmit_module.n144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_15_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_15_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i6_LC_15_15_2  (
            .in0(N__20254),
            .in1(N__15200),
            .in2(N__19951),
            .in3(N__15188),
            .lcout(\transmit_module.TX_ADDR_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23383),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i3_3_lut_LC_15_16_2 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i3_3_lut_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i3_3_lut_LC_15_16_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i3_3_lut_LC_15_16_2  (
            .in0(N__20577),
            .in1(N__15114),
            .in2(_gnd_net_),
            .in3(N__15044),
            .lcout(\transmit_module.n145 ),
            .ltout(\transmit_module.n145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i2_LC_15_16_3 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i2_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i2_LC_15_16_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i2_LC_15_16_3  (
            .in0(N__20037),
            .in1(N__20255),
            .in2(N__15785),
            .in3(N__20552),
            .lcout(\transmit_module.TX_ADDR_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23133),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i3_LC_15_16_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i3_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i3_LC_15_16_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i3_LC_15_16_7  (
            .in0(N__20256),
            .in1(N__19517),
            .in2(N__20066),
            .in3(N__19495),
            .lcout(\transmit_module.TX_ADDR_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23133),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_15_17_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_15_17_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_15_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i1_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15782),
            .lcout(\transmit_module.Y_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23404),
            .ce(N__21406),
            .sr(N__20041));
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_15_17_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_15_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i2_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15761),
            .lcout(\transmit_module.Y_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23404),
            .ce(N__21406),
            .sr(N__20041));
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_15_17_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_15_17_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_15_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i4_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15776),
            .lcout(\transmit_module.Y_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23404),
            .ce(N__21406),
            .sr(N__20041));
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_15_17_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_15_17_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_15_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i3_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15767),
            .lcout(\transmit_module.Y_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23404),
            .ce(N__21406),
            .sr(N__20041));
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_15_18_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_15_18_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_15_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i0_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15755),
            .lcout(\transmit_module.Y_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23232),
            .ce(N__21405),
            .sr(N__19912));
    defparam \receive_module.BRAM_ADDR__i1_LC_15_19_0 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i1_LC_15_19_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i1_LC_15_19_0 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \receive_module.BRAM_ADDR__i1_LC_15_19_0  (
            .in0(N__18892),
            .in1(N__15749),
            .in2(N__18753),
            .in3(N__15515),
            .lcout(RX_ADDR_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24141),
            .ce(),
            .sr(N__17542));
    defparam \receive_module.BRAM_ADDR__i2_LC_15_19_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i2_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i2_LC_15_19_2 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \receive_module.BRAM_ADDR__i2_LC_15_19_2  (
            .in0(N__15491),
            .in1(N__18895),
            .in2(N__18754),
            .in3(N__15272),
            .lcout(RX_ADDR_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24141),
            .ce(),
            .sr(N__17542));
    defparam \receive_module.BRAM_ADDR__i4_LC_15_19_4 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i4_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i4_LC_15_19_4 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \receive_module.BRAM_ADDR__i4_LC_15_19_4  (
            .in0(N__18893),
            .in1(N__17453),
            .in2(N__18755),
            .in3(N__17219),
            .lcout(RX_ADDR_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24141),
            .ce(),
            .sr(N__17542));
    defparam \receive_module.BRAM_ADDR__i5_LC_15_19_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i5_LC_15_19_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i5_LC_15_19_5 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \receive_module.BRAM_ADDR__i5_LC_15_19_5  (
            .in0(N__18896),
            .in1(N__17189),
            .in2(N__16976),
            .in3(N__18733),
            .lcout(RX_ADDR_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24141),
            .ce(),
            .sr(N__17542));
    defparam \receive_module.BRAM_ADDR__i6_LC_15_19_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i6_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i6_LC_15_19_6 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \receive_module.BRAM_ADDR__i6_LC_15_19_6  (
            .in0(N__18894),
            .in1(N__16700),
            .in2(N__18756),
            .in3(N__16934),
            .lcout(RX_ADDR_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24141),
            .ce(),
            .sr(N__17542));
    defparam \receive_module.BRAM_ADDR__i7_LC_15_19_7 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i7_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i7_LC_15_19_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \receive_module.BRAM_ADDR__i7_LC_15_19_7  (
            .in0(N__18897),
            .in1(N__18737),
            .in2(N__16457),
            .in3(N__16673),
            .lcout(RX_ADDR_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24141),
            .ce(),
            .sr(N__17542));
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_20_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_20_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i4_3_lut_LC_15_20_1  (
            .in0(N__20655),
            .in1(N__16418),
            .in2(_gnd_net_),
            .in3(N__16405),
            .lcout(\transmit_module.n113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i9_LC_15_23_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i9_LC_15_23_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i9_LC_15_23_3 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \receive_module.BRAM_ADDR__i9_LC_15_23_3  (
            .in0(N__18908),
            .in1(N__16145),
            .in2(N__18768),
            .in3(N__16373),
            .lcout(RX_ADDR_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24146),
            .ce(),
            .sr(N__17555));
    defparam GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_15_24_3.C_ON=1'b0;
    defparam GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_15_24_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_15_24_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_15_24_3 (
            .in0(N__24173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_DEBUG_c_3_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i1_LC_15_25_3 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i1_LC_15_25_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i1_LC_15_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i1_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22070),
            .lcout(n1821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22876),
            .ce(),
            .sr(N__22688));
    defparam \receive_module.BRAM_ADDR__i8_LC_15_27_4 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i8_LC_15_27_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i8_LC_15_27_4 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \receive_module.BRAM_ADDR__i8_LC_15_27_4  (
            .in0(N__18918),
            .in1(N__15812),
            .in2(N__18777),
            .in3(N__16034),
            .lcout(RX_ADDR_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24155),
            .ce(),
            .sr(N__17565));
    defparam \receive_module.BRAM_ADDR__i0_LC_15_28_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i0_LC_15_28_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i0_LC_15_28_3 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \receive_module.BRAM_ADDR__i0_LC_15_28_3  (
            .in0(N__18919),
            .in1(N__18302),
            .in2(N__18766),
            .in3(N__18080),
            .lcout(RX_ADDR_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24157),
            .ce(),
            .sr(N__17566));
    defparam \receive_module.BRAM_ADDR__i3_LC_15_31_1 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i3_LC_15_31_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i3_LC_15_31_1 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \receive_module.BRAM_ADDR__i3_LC_15_31_1  (
            .in0(N__18926),
            .in1(N__18056),
            .in2(N__18785),
            .in3(N__17846),
            .lcout(RX_ADDR_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24161),
            .ce(),
            .sr(N__17570));
    defparam \receive_module.BRAM_ADDR__i10_LC_15_31_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i10_LC_15_31_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i10_LC_15_31_3 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \receive_module.BRAM_ADDR__i10_LC_15_31_3  (
            .in0(N__18925),
            .in1(N__17597),
            .in2(N__18784),
            .in3(N__17822),
            .lcout(RX_ADDR_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24161),
            .ce(),
            .sr(N__17570));
    defparam PULSE_1HZ_I_0_2_lut_LC_16_6_1.C_ON=1'b0;
    defparam PULSE_1HZ_I_0_2_lut_LC_16_6_1.SEQ_MODE=4'b0000;
    defparam PULSE_1HZ_I_0_2_lut_LC_16_6_1.LUT_INIT=16'b1111111110101010;
    LogicCell40 PULSE_1HZ_I_0_2_lut_LC_16_6_1 (
            .in0(N__18805),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17477),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_16_8_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_16_8_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \receive_module.rx_counter.PULSE_1HZ_49_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__17473),
            .in2(_gnd_net_),
            .in3(N__18428),
            .lcout(PULSE_1HZ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24103),
            .ce(N__18326),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_26_LC_16_9_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_26_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_26_LC_16_9_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_26_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__18355),
            .in2(_gnd_net_),
            .in3(N__18385),
            .lcout(\receive_module.rx_counter.n7_adj_619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i134_2_lut_rep_16_2_lut_LC_16_9_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i134_2_lut_rep_16_2_lut_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i134_2_lut_rep_16_2_lut_LC_16_9_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \receive_module.rx_counter.i134_2_lut_rep_16_2_lut_LC_16_9_1  (
            .in0(N__18871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17462),
            .lcout(\receive_module.rx_counter.n3675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1307_2_lut_3_lut_3_lut_LC_16_9_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1307_2_lut_3_lut_3_lut_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1307_2_lut_3_lut_3_lut_LC_16_9_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \receive_module.rx_counter.i1307_2_lut_3_lut_3_lut_LC_16_9_4  (
            .in0(N__17461),
            .in1(N__18870),
            .in2(_gnd_net_),
            .in3(N__18427),
            .lcout(\receive_module.rx_counter.n2550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_VS_52_LC_16_9_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_VS_52_LC_16_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_VS_52_LC_16_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receive_module.rx_counter.old_VS_52_LC_16_9_5  (
            .in0(N__18872),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.rx_counter.old_VS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24107),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2185_2_lut_LC_16_9_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2185_2_lut_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2185_2_lut_LC_16_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i2185_2_lut_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__18400),
            .in2(_gnd_net_),
            .in3(N__18337),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3522_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_4_lut_LC_16_9_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_4_lut_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_4_lut_LC_16_9_7 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \receive_module.rx_counter.i5_4_lut_LC_16_9_7  (
            .in0(N__18415),
            .in1(N__18370),
            .in2(N__18437),
            .in3(N__18434),
            .lcout(\receive_module.rx_counter.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i0_LC_16_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i0_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i0_LC_16_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_247__i0_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__18416),
            .in2(_gnd_net_),
            .in3(N__18404),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_0 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\receive_module.rx_counter.n3205 ),
            .clk(N__24112),
            .ce(N__18325),
            .sr(N__19163));
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i1_LC_16_10_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i1_LC_16_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i1_LC_16_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_247__i1_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__18401),
            .in2(_gnd_net_),
            .in3(N__18389),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3205 ),
            .carryout(\receive_module.rx_counter.n3206 ),
            .clk(N__24112),
            .ce(N__18325),
            .sr(N__19163));
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i2_LC_16_10_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i2_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i2_LC_16_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_247__i2_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__18386),
            .in2(_gnd_net_),
            .in3(N__18374),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3206 ),
            .carryout(\receive_module.rx_counter.n3207 ),
            .clk(N__24112),
            .ce(N__18325),
            .sr(N__19163));
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i3_LC_16_10_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i3_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i3_LC_16_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_247__i3_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__18371),
            .in2(_gnd_net_),
            .in3(N__18359),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3207 ),
            .carryout(\receive_module.rx_counter.n3208 ),
            .clk(N__24112),
            .ce(N__18325),
            .sr(N__19163));
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i4_LC_16_10_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i4_LC_16_10_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i4_LC_16_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_247__i4_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__18356),
            .in2(_gnd_net_),
            .in3(N__18344),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3208 ),
            .carryout(\receive_module.rx_counter.n3209 ),
            .clk(N__24112),
            .ce(N__18325),
            .sr(N__19163));
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i5_LC_16_10_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i5_LC_16_10_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_247__i5_LC_16_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_247__i5_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__18338),
            .in2(_gnd_net_),
            .in3(N__18341),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24112),
            .ce(N__18325),
            .sr(N__19163));
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_16_11_3 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_16_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i4_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19157),
            .lcout(RX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24116),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.sync_wd.i2_2_lut_LC_16_12_1 .C_ON=1'b0;
    defparam \receive_module.sync_wd.i2_2_lut_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.sync_wd.i2_2_lut_LC_16_12_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.sync_wd.i2_2_lut_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__19081),
            .in2(_gnd_net_),
            .in3(N__18525),
            .lcout(),
            .ltout(\receive_module.sync_wd.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.sync_wd.i1_4_lut_LC_16_12_2 .C_ON=1'b0;
    defparam \receive_module.sync_wd.i1_4_lut_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.sync_wd.i1_4_lut_LC_16_12_2 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \receive_module.sync_wd.i1_4_lut_LC_16_12_2  (
            .in0(N__18959),
            .in1(N__22456),
            .in2(N__18932),
            .in3(N__18680),
            .lcout(),
            .ltout(\receive_module.sync_wd.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.sync_wd.SYNC_BAD_16_LC_16_12_3 .C_ON=1'b0;
    defparam \receive_module.sync_wd.SYNC_BAD_16_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.sync_wd.SYNC_BAD_16_LC_16_12_3 .LUT_INIT=16'b1100111000000000;
    LogicCell40 \receive_module.sync_wd.SYNC_BAD_16_LC_16_12_3  (
            .in0(N__18602),
            .in1(N__18798),
            .in2(N__18929),
            .in3(N__18854),
            .lcout(DEBUG_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24119),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.sync_wd.old_visible_17_LC_16_12_6 .C_ON=1'b0;
    defparam \receive_module.sync_wd.old_visible_17_LC_16_12_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.sync_wd.old_visible_17_LC_16_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receive_module.sync_wd.old_visible_17_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18681),
            .lcout(\receive_module.sync_wd.old_visible ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24119),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_16_13_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_16_13_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_16_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i7_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22532),
            .lcout(RX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24125),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_14_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_14_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_14_5  (
            .in0(N__24764),
            .in1(N__18500),
            .in2(N__22376),
            .in3(N__18482),
            .lcout(\line_buffer.n3656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2260_LC_16_15_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2260_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2260_LC_16_15_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2260_LC_16_15_2  (
            .in0(N__24772),
            .in1(N__18467),
            .in2(N__22377),
            .in3(N__18449),
            .lcout(\line_buffer.n3590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i1_LC_16_15_7 .C_ON=1'b0;
    defparam \line_buffer.dout_i1_LC_16_15_7 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i1_LC_16_15_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i1_LC_16_15_7  (
            .in0(N__23940),
            .in1(N__21242),
            .in2(_gnd_net_),
            .in3(N__21209),
            .lcout(TX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22908),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_16_16_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_16_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_16_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i4_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20810),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23132),
            .ce(N__20757),
            .sr(N__19911));
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20578),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23375),
            .ce(N__20771),
            .sr(N__20042));
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_18_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_18_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_12_i3_3_lut_LC_16_18_3  (
            .in0(N__20690),
            .in1(N__20626),
            .in2(_gnd_net_),
            .in3(N__20579),
            .lcout(\transmit_module.n114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1647_4_lut_LC_16_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1647_4_lut_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1647_4_lut_LC_16_19_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1647_4_lut_LC_16_19_0  (
            .in0(N__20257),
            .in1(N__20548),
            .in2(N__20013),
            .in3(N__20537),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3626_bdd_4_lut_LC_16_19_2 .C_ON=1'b0;
    defparam \line_buffer.n3626_bdd_4_lut_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3626_bdd_4_lut_LC_16_19_2 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3626_bdd_4_lut_LC_16_19_2  (
            .in0(N__20306),
            .in1(N__22339),
            .in2(N__20285),
            .in3(N__21779),
            .lcout(\line_buffer.n3629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1648_4_lut_LC_16_19_3 .C_ON=1'b0;
    defparam \transmit_module.i1648_4_lut_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1648_4_lut_LC_16_19_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.i1648_4_lut_LC_16_19_3  (
            .in0(N__20258),
            .in1(N__19910),
            .in2(N__19516),
            .in3(N__19499),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i4_LC_16_20_3 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i4_LC_16_20_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i4_LC_16_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i4_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21074),
            .lcout(n1818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22987),
            .ce(),
            .sr(N__22649));
    defparam \line_buffer.n3590_bdd_4_lut_LC_16_21_3 .C_ON=1'b0;
    defparam \line_buffer.n3590_bdd_4_lut_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3590_bdd_4_lut_LC_16_21_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.n3590_bdd_4_lut_LC_16_21_3  (
            .in0(N__22375),
            .in1(N__19205),
            .in2(N__19193),
            .in3(N__19172),
            .lcout(),
            .ltout(\line_buffer.n3593_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i3_LC_16_21_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i3_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i3_LC_16_21_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i3_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__23932),
            .in2(N__21086),
            .in3(N__21083),
            .lcout(TX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23201),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2214_3_lut_LC_16_22_5 .C_ON=1'b0;
    defparam \line_buffer.i2214_3_lut_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2214_3_lut_LC_16_22_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2214_3_lut_LC_16_22_5  (
            .in0(N__21068),
            .in1(N__21053),
            .in2(_gnd_net_),
            .in3(N__24797),
            .lcout(),
            .ltout(\line_buffer.n3551_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i4_LC_16_22_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i4_LC_16_22_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i4_LC_16_22_6 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.dout_i4_LC_16_22_6  (
            .in0(N__23938),
            .in1(N__21035),
            .in2(N__21020),
            .in3(N__21692),
            .lcout(TX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23039),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2200_3_lut_LC_16_23_0 .C_ON=1'b0;
    defparam \line_buffer.i2200_3_lut_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2200_3_lut_LC_16_23_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2200_3_lut_LC_16_23_0  (
            .in0(N__24796),
            .in1(N__21017),
            .in2(_gnd_net_),
            .in3(N__20996),
            .lcout(\line_buffer.n3537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i5_LC_16_24_4 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i5_LC_16_24_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i5_LC_16_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i5_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20978),
            .lcout(n1817),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23125),
            .ce(),
            .sr(N__22680));
    defparam \transmit_module.VGA_R__i2_LC_16_25_2 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i2_LC_16_25_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i2_LC_16_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i2_LC_16_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20906),
            .lcout(n1820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22869),
            .ce(),
            .sr(N__22692));
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_17_9_0 .C_ON=1'b0;
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_17_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_hs_buffer.BUFFER_0__i2_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21608),
            .lcout(\tvp_hs_buffer.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24101),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2199_3_lut_LC_17_9_2 .C_ON=1'b0;
    defparam \line_buffer.i2199_3_lut_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2199_3_lut_LC_17_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2199_3_lut_LC_17_9_2  (
            .in0(N__24794),
            .in1(N__20840),
            .in2(_gnd_net_),
            .in3(N__20822),
            .lcout(\line_buffer.n3536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2235_3_lut_LC_17_10_6 .C_ON=1'b0;
    defparam \line_buffer.i2235_3_lut_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2235_3_lut_LC_17_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2235_3_lut_LC_17_10_6  (
            .in0(N__24795),
            .in1(N__21521),
            .in2(_gnd_net_),
            .in3(N__21503),
            .lcout(\line_buffer.n3572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_17_14_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_17_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i5_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21494),
            .lcout(\transmit_module.X_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23487),
            .ce(N__21474),
            .sr(N__21354));
    defparam \line_buffer.n3650_bdd_4_lut_LC_17_15_3 .C_ON=1'b0;
    defparam \line_buffer.n3650_bdd_4_lut_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3650_bdd_4_lut_LC_17_15_3 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3650_bdd_4_lut_LC_17_15_3  (
            .in0(N__21278),
            .in1(N__22346),
            .in2(N__21260),
            .in3(N__21878),
            .lcout(\line_buffer.n3653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3632_bdd_4_lut_LC_17_16_4 .C_ON=1'b0;
    defparam \line_buffer.n3632_bdd_4_lut_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3632_bdd_4_lut_LC_17_16_4 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n3632_bdd_4_lut_LC_17_16_4  (
            .in0(N__21236),
            .in1(N__21149),
            .in2(N__21224),
            .in3(N__22350),
            .lcout(\line_buffer.n3635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2233_3_lut_LC_17_16_6 .C_ON=1'b0;
    defparam \line_buffer.i2233_3_lut_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2233_3_lut_LC_17_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2233_3_lut_LC_17_16_6  (
            .in0(N__21203),
            .in1(N__21185),
            .in2(_gnd_net_),
            .in3(N__24686),
            .lcout(\line_buffer.n3570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2294_LC_17_17_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2294_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2294_LC_17_17_1 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2294_LC_17_17_1  (
            .in0(N__24745),
            .in1(N__21176),
            .in2(N__22372),
            .in3(N__21167),
            .lcout(\line_buffer.n3632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2269_LC_17_17_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2269_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2269_LC_17_17_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2269_LC_17_17_2  (
            .in0(N__22337),
            .in1(N__21566),
            .in2(N__23950),
            .in3(N__21143),
            .lcout(),
            .ltout(\line_buffer.n3602_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i2_LC_17_17_3 .C_ON=1'b0;
    defparam \line_buffer.dout_i2_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i2_LC_17_17_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.dout_i2_LC_17_17_3  (
            .in0(N__23944),
            .in1(N__21656),
            .in2(N__21131),
            .in3(N__21128),
            .lcout(TX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23336),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3656_bdd_4_lut_LC_17_18_5 .C_ON=1'b0;
    defparam \line_buffer.n3656_bdd_4_lut_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3656_bdd_4_lut_LC_17_18_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3656_bdd_4_lut_LC_17_18_5  (
            .in0(N__21122),
            .in1(N__22338),
            .in2(N__21107),
            .in3(N__21818),
            .lcout(\line_buffer.n3659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2289_LC_17_19_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2289_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2289_LC_17_19_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2289_LC_17_19_3  (
            .in0(N__24765),
            .in1(N__21806),
            .in2(N__22373),
            .in3(N__21791),
            .lcout(\line_buffer.n3626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i3_LC_17_21_2 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i3_LC_17_21_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i3_LC_17_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i3_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21773),
            .lcout(n1819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23227),
            .ce(),
            .sr(N__22687));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2279_LC_17_22_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2279_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2279_LC_17_22_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2279_LC_17_22_4  (
            .in0(N__22374),
            .in1(N__21710),
            .in2(N__23949),
            .in3(N__21704),
            .lcout(\line_buffer.n3614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2232_3_lut_LC_17_25_7 .C_ON=1'b0;
    defparam \line_buffer.i2232_3_lut_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2232_3_lut_LC_17_25_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2232_3_lut_LC_17_25_7  (
            .in0(N__21686),
            .in1(N__21674),
            .in2(_gnd_net_),
            .in3(N__24743),
            .lcout(\line_buffer.n3569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_0 .C_ON=1'b0;
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_0 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21628),
            .lcout(\tvp_hs_buffer.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24108),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2236_3_lut_LC_18_17_5 .C_ON=1'b0;
    defparam \line_buffer.i2236_3_lut_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2236_3_lut_LC_18_17_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2236_3_lut_LC_18_17_5  (
            .in0(N__24763),
            .in1(N__21602),
            .in2(_gnd_net_),
            .in3(N__21587),
            .lcout(\line_buffer.n3573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i5_LC_18_18_1 .C_ON=1'b0;
    defparam \line_buffer.dout_i5_LC_18_18_1 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i5_LC_18_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i5_LC_18_18_1  (
            .in0(N__23939),
            .in1(N__21908),
            .in2(_gnd_net_),
            .in3(N__21560),
            .lcout(TX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23570),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2299_LC_18_19_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2299_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2299_LC_18_19_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2299_LC_18_19_3  (
            .in0(N__24784),
            .in1(N__21554),
            .in2(N__22381),
            .in3(N__21536),
            .lcout(\line_buffer.n3638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3638_bdd_4_lut_LC_18_21_0 .C_ON=1'b0;
    defparam \line_buffer.n3638_bdd_4_lut_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3638_bdd_4_lut_LC_18_21_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3638_bdd_4_lut_LC_18_21_0  (
            .in0(N__22124),
            .in1(N__22389),
            .in2(N__22109),
            .in3(N__22085),
            .lcout(\line_buffer.n3641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i0_LC_18_22_1 .C_ON=1'b0;
    defparam \line_buffer.dout_i0_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i0_LC_18_22_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \line_buffer.dout_i0_LC_18_22_1  (
            .in0(N__23937),
            .in1(N__22076),
            .in2(_gnd_net_),
            .in3(N__22010),
            .lcout(TX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23439),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3644_bdd_4_lut_LC_18_23_3 .C_ON=1'b0;
    defparam \line_buffer.n3644_bdd_4_lut_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3644_bdd_4_lut_LC_18_23_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.n3644_bdd_4_lut_LC_18_23_3  (
            .in0(N__22390),
            .in1(N__22058),
            .in2(N__22034),
            .in3(N__22577),
            .lcout(\line_buffer.n3647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i6_LC_18_25_7 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i6_LC_18_25_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i6_LC_18_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i6_LC_18_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22004),
            .lcout(n1816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23038),
            .ce(),
            .sr(N__22694));
    defparam \line_buffer.n3596_bdd_4_lut_LC_19_17_1 .C_ON=1'b0;
    defparam \line_buffer.n3596_bdd_4_lut_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3596_bdd_4_lut_LC_19_17_1 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3596_bdd_4_lut_LC_19_17_1  (
            .in0(N__21950),
            .in1(N__22391),
            .in2(N__21932),
            .in3(N__22175),
            .lcout(\line_buffer.n3599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2309_LC_19_19_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2309_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2309_LC_19_19_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2309_LC_19_19_5  (
            .in0(N__24785),
            .in1(N__21902),
            .in2(N__22393),
            .in3(N__21893),
            .lcout(\line_buffer.n3650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2239_3_lut_LC_19_19_7 .C_ON=1'b0;
    defparam \line_buffer.i2239_3_lut_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2239_3_lut_LC_19_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2239_3_lut_LC_19_19_7  (
            .in0(N__24786),
            .in1(N__21866),
            .in2(_gnd_net_),
            .in3(N__21848),
            .lcout(\line_buffer.n3576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2274_LC_19_21_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2274_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2274_LC_19_21_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2274_LC_19_21_0  (
            .in0(N__22388),
            .in1(N__21827),
            .in2(N__23951),
            .in3(N__24530),
            .lcout(),
            .ltout(\line_buffer.n3608_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i6_LC_19_21_1 .C_ON=1'b0;
    defparam \line_buffer.dout_i6_LC_19_21_1 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i6_LC_19_21_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.dout_i6_LC_19_21_1  (
            .in0(N__23948),
            .in1(N__22541),
            .in2(N__23813),
            .in3(N__23810),
            .lcout(TX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23248),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i7_LC_19_22_1 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i7_LC_19_22_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i7_LC_19_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i7_LC_19_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23801),
            .lcout(n1815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23440),
            .ce(),
            .sr(N__22693));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2304_LC_19_23_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2304_LC_19_23_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2304_LC_19_23_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2304_LC_19_23_0  (
            .in0(N__24799),
            .in1(N__22613),
            .in2(N__22394),
            .in3(N__22598),
            .lcout(\line_buffer.n3644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2238_3_lut_LC_19_25_7 .C_ON=1'b0;
    defparam \line_buffer.i2238_3_lut_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2238_3_lut_LC_19_25_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2238_3_lut_LC_19_25_7  (
            .in0(N__22571),
            .in1(N__22556),
            .in2(_gnd_net_),
            .in3(N__24744),
            .lcout(\line_buffer.n3575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_20_13_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_20_13_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_20_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i16_LC_20_13_0  (
            .in0(N__24185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24132),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_20_17_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_20_17_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_20_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i5_LC_20_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24806),
            .lcout(RX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24139),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2284_LC_20_17_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2284_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2284_LC_20_17_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2284_LC_20_17_1  (
            .in0(N__24793),
            .in1(N__22406),
            .in2(N__22392),
            .in3(N__22193),
            .lcout(\line_buffer.n3596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_20_17_4 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_20_17_4 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_20_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i6_LC_20_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22165),
            .lcout(\tvp_video_buffer.BUFFER_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24139),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_20_17_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_20_17_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_20_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i14_LC_20_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24812),
            .lcout(\tvp_video_buffer.BUFFER_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24139),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2205_3_lut_LC_20_21_0 .C_ON=1'b0;
    defparam \line_buffer.i2205_3_lut_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2205_3_lut_LC_20_21_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2205_3_lut_LC_20_21_0  (
            .in0(N__24800),
            .in1(N__24566),
            .in2(_gnd_net_),
            .in3(N__24551),
            .lcout(\line_buffer.n3542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_22_19_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_22_19_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_22_19_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_22_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_24_9_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_24_9_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_24_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i8_LC_24_9_5  (
            .in0(N__24194),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24133),
            .ce(),
            .sr(_gnd_net_));
endmodule // main
