-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 15 2018 02:00:50

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    TVP_VIDEO : in std_logic_vector(9 downto 0);
    ADV_B : out std_logic_vector(7 downto 0);
    ADV_G : out std_logic_vector(7 downto 0);
    ADV_R : out std_logic_vector(7 downto 0);
    DEBUG : inout std_logic_vector(7 downto 0);
    TVP_CLK : in std_logic;
    ADV_CLK : out std_logic;
    TVP_HSYNC : in std_logic;
    ADV_HSYNC : out std_logic;
    TVP_VSYNC : in std_logic;
    ADV_VSYNC : out std_logic;
    ADV_BLANK_N : out std_logic;
    LED : out std_logic;
    ADV_SYNC_N : out std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7876\ : std_logic;
signal \TVP_VIDEO_c_3\ : std_logic;
signal \VCCG0\ : std_logic;
signal \TVP_VIDEO_c_5\ : std_logic;
signal \TVP_VIDEO_c_4\ : std_logic;
signal \GNDG0\ : std_logic;
signal \TVP_VIDEO_c_7\ : std_logic;
signal \TVP_VIDEO_c_6\ : std_logic;
signal \TVP_VIDEO_c_8\ : std_logic;
signal \TVP_VIDEO_c_9\ : std_logic;
signal \TVP_VIDEO_c_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_55\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_54\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_53\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_52\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_16\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_17\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_19\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_18\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_71\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_70\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_60\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_59\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_42\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_41\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_69\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_56\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_58\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_57\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_61\ : std_logic;
signal \line_buffer.n639\ : std_logic;
signal \line_buffer.n631\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_24\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_20\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_21\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_23\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_22\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_45\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_77\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_46\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_78\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_68\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_79\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_48\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_47\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_67\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_82\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_44\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_43\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_81\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_80\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_66\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_76\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_75\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_51\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_63\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_62\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_74\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_50\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_49\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_65\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_64\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_13\ : std_logic;
signal \old_HS\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \receive_module.rx_counter.n3349\ : std_logic;
signal \receive_module.rx_counter.n3350\ : std_logic;
signal \receive_module.rx_counter.n3351\ : std_logic;
signal \receive_module.rx_counter.n3352\ : std_logic;
signal \receive_module.rx_counter.n3353\ : std_logic;
signal \receive_module.rx_counter.n3354\ : std_logic;
signal \receive_module.rx_counter.n3355\ : std_logic;
signal \receive_module.rx_counter.n3356\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal n2057 : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_26\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_25\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_27\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_83\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_84\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_95\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_94\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_93\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_85\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_86\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_92\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_91\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3377\ : std_logic;
signal \transmit_module.video_signal_controller.n3378\ : std_logic;
signal \transmit_module.video_signal_controller.n3379\ : std_logic;
signal \transmit_module.video_signal_controller.n3380\ : std_logic;
signal \transmit_module.video_signal_controller.n3381\ : std_logic;
signal \transmit_module.video_signal_controller.n3382\ : std_logic;
signal \transmit_module.video_signal_controller.n3383\ : std_logic;
signal \transmit_module.video_signal_controller.n3384\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3385\ : std_logic;
signal \transmit_module.video_signal_controller.n3386\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_28\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_29\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_30\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_31\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_73\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_72\ : std_logic;
signal n22 : std_logic;
signal \transmit_module.X_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_14\ : std_logic;
signal \line_buffer.n630\ : std_logic;
signal \line_buffer.n638\ : std_logic;
signal \receive_module.rx_counter.Y_6\ : std_logic;
signal \receive_module.rx_counter.Y_5\ : std_logic;
signal \receive_module.rx_counter.n3619_cascade_\ : std_logic;
signal \line_buffer.n642\ : std_logic;
signal \line_buffer.n578\ : std_logic;
signal \receive_module.rx_counter.n14_cascade_\ : std_logic;
signal \receive_module.rx_counter.Y_8\ : std_logic;
signal \receive_module.rx_counter.Y_7\ : std_logic;
signal \receive_module.rx_counter.n15_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3861\ : std_logic;
signal \receive_module.rx_counter.Y_0\ : std_logic;
signal \receive_module.rx_counter.n10_adj_570\ : std_logic;
signal \receive_module.rx_counter.Y_2\ : std_logic;
signal \line_buffer.n610\ : std_logic;
signal \line_buffer.n512\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_99\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_90\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_87\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_89\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_88\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_98\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_97\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_96\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_1\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_2\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_0\ : std_logic;
signal \transmit_module.video_signal_controller.n8_adj_569_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3029_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3857_cascade_\ : std_logic;
signal \transmit_module.n2125\ : std_logic;
signal \transmit_module.n3859_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_7\ : std_logic;
signal \transmit_module.video_signal_controller.n4_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_6\ : std_logic;
signal \transmit_module.video_signal_controller.n23_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_10\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_9\ : std_logic;
signal \transmit_module.n214\ : std_logic;
signal \transmit_module.n182\ : std_logic;
signal \transmit_module.n214_cascade_\ : std_logic;
signal n20 : std_logic;
signal \transmit_module.n215_cascade_\ : std_logic;
signal n23 : std_logic;
signal \transmit_module.n183\ : std_logic;
signal \transmit_module.n215\ : std_logic;
signal \transmit_module.n212\ : std_logic;
signal \transmit_module.n180\ : std_logic;
signal \transmit_module.n212_cascade_\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_6\ : std_logic;
signal \line_buffer.n574\ : std_logic;
signal \line_buffer.n3785\ : std_logic;
signal \line_buffer.n566\ : std_logic;
signal \line_buffer.n577\ : std_logic;
signal \line_buffer.n513\ : std_logic;
signal \receive_module.rx_counter.Y_4\ : std_logic;
signal \receive_module.rx_counter.n4\ : std_logic;
signal \receive_module.rx_counter.Y_3\ : std_logic;
signal \receive_module.rx_counter.Y_1\ : std_logic;
signal \receive_module.rx_counter.n3657\ : std_logic;
signal \receive_module.rx_counter.n3619\ : std_logic;
signal \receive_module.rx_counter.n3648_cascade_\ : std_logic;
signal \DEBUG_c_5_cascade_\ : std_logic;
signal \line_buffer.n641\ : std_logic;
signal \line_buffer.n609\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \receive_module.rx_counter.n3387\ : std_logic;
signal \receive_module.rx_counter.n3388\ : std_logic;
signal \receive_module.rx_counter.n3389\ : std_logic;
signal \receive_module.rx_counter.n3390\ : std_logic;
signal \receive_module.rx_counter.n3391\ : std_logic;
signal \DEBUG_c_5\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_4\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_3\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_5\ : std_logic;
signal \transmit_module.video_signal_controller.n21\ : std_logic;
signal \transmit_module.video_signal_controller.n3023_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3697_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n8\ : std_logic;
signal \transmit_module.video_signal_controller.n3577\ : std_logic;
signal \transmit_module.video_signal_controller.n6_adj_568_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3603\ : std_logic;
signal \transmit_module.video_signal_controller.n6_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3575\ : std_logic;
signal \transmit_module.video_signal_controller.n2015\ : std_logic;
signal \transmit_module.video_signal_controller.n3857\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_8\ : std_logic;
signal \transmit_module.video_signal_controller.n3856\ : std_logic;
signal \transmit_module.n220_cascade_\ : std_logic;
signal n28 : std_logic;
signal \transmit_module.BRAM_ADDR_13_N_256_13\ : std_logic;
signal \transmit_module.n219_cascade_\ : std_logic;
signal n27 : std_logic;
signal n1850 : std_logic;
signal n1849 : std_logic;
signal n1848 : std_logic;
signal n1847 : std_logic;
signal n1846 : std_logic;
signal n1845 : std_logic;
signal n1844 : std_logic;
signal \ADV_B_c\ : std_logic;
signal \INVADV_R__i1C_net\ : std_logic;
signal n2404 : std_logic;
signal \transmit_module.n220\ : std_logic;
signal \transmit_module.n218_cascade_\ : std_logic;
signal n26 : std_logic;
signal \transmit_module.n187\ : std_logic;
signal \transmit_module.n219\ : std_logic;
signal \transmit_module.n187_cascade_\ : std_logic;
signal \transmit_module.n218\ : std_logic;
signal \transmit_module.n186\ : std_logic;
signal \transmit_module.n204\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \transmit_module.n203\ : std_logic;
signal \transmit_module.n3336\ : std_logic;
signal \transmit_module.n202\ : std_logic;
signal \transmit_module.n3337\ : std_logic;
signal \transmit_module.n3338\ : std_logic;
signal \transmit_module.n3339\ : std_logic;
signal \transmit_module.n199\ : std_logic;
signal \transmit_module.n3340\ : std_logic;
signal \transmit_module.n198\ : std_logic;
signal \transmit_module.n3341\ : std_logic;
signal \transmit_module.n3342\ : std_logic;
signal \transmit_module.n3343\ : std_logic;
signal \transmit_module.n196\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \transmit_module.n3344\ : std_logic;
signal \transmit_module.n3345\ : std_logic;
signal \transmit_module.n193\ : std_logic;
signal \transmit_module.n3346\ : std_logic;
signal \transmit_module.n192\ : std_logic;
signal \transmit_module.n3347\ : std_logic;
signal \transmit_module.n3348\ : std_logic;
signal \transmit_module.n191\ : std_logic;
signal \transmit_module.TX_ADDR_8\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_8\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.n2099\ : std_logic;
signal \line_buffer.n3788\ : std_logic;
signal \TX_DATA_6\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_4\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_2\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_5\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_1\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_0\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_3\ : std_logic;
signal \receive_module.rx_counter.n3693_cascade_\ : std_logic;
signal \receive_module.rx_counter.n7\ : std_logic;
signal \receive_module.rx_counter.n11_cascade_\ : std_logic;
signal \receive_module.rx_counter.PULSE_1HZ_N_94\ : std_logic;
signal \receive_module.rx_counter.n2562\ : std_logic;
signal \RX_ADDR_0\ : std_logic;
signal \receive_module.n136\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \RX_ADDR_1\ : std_logic;
signal \receive_module.n135\ : std_logic;
signal \receive_module.n3323\ : std_logic;
signal \RX_ADDR_2\ : std_logic;
signal \receive_module.n134\ : std_logic;
signal \receive_module.n3324\ : std_logic;
signal \RX_ADDR_3\ : std_logic;
signal \receive_module.n133\ : std_logic;
signal \receive_module.n3325\ : std_logic;
signal \RX_ADDR_4\ : std_logic;
signal \receive_module.n132\ : std_logic;
signal \receive_module.n3326\ : std_logic;
signal \RX_ADDR_5\ : std_logic;
signal \receive_module.n131\ : std_logic;
signal \receive_module.n3327\ : std_logic;
signal \RX_ADDR_6\ : std_logic;
signal \receive_module.n130\ : std_logic;
signal \receive_module.n3328\ : std_logic;
signal \RX_ADDR_7\ : std_logic;
signal \receive_module.n129\ : std_logic;
signal \receive_module.n3329\ : std_logic;
signal \receive_module.n3330\ : std_logic;
signal \RX_ADDR_8\ : std_logic;
signal \receive_module.n128\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \RX_ADDR_9\ : std_logic;
signal \receive_module.n127\ : std_logic;
signal \receive_module.n3331\ : std_logic;
signal \RX_ADDR_10\ : std_logic;
signal \receive_module.n126\ : std_logic;
signal \receive_module.n3332\ : std_logic;
signal \RX_ADDR_11\ : std_logic;
signal \receive_module.n3333\ : std_logic;
signal \RX_ADDR_12\ : std_logic;
signal \receive_module.n3334\ : std_logic;
signal \receive_module.n3854\ : std_logic;
signal \DEBUG_c_3\ : std_logic;
signal \receive_module.n3335\ : std_logic;
signal \receive_module.n123\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_0\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_1\ : std_logic;
signal \transmit_module.video_signal_controller.n3366\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_2\ : std_logic;
signal \transmit_module.video_signal_controller.n3367\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_3\ : std_logic;
signal \transmit_module.video_signal_controller.n3368\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_4\ : std_logic;
signal \transmit_module.video_signal_controller.n3369\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_5\ : std_logic;
signal \transmit_module.video_signal_controller.n3370\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_6\ : std_logic;
signal \transmit_module.video_signal_controller.n3371\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_7\ : std_logic;
signal \transmit_module.video_signal_controller.n3372\ : std_logic;
signal \transmit_module.video_signal_controller.n3373\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_8\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_9\ : std_logic;
signal \transmit_module.video_signal_controller.n3374\ : std_logic;
signal \transmit_module.video_signal_controller.n3375\ : std_logic;
signal \transmit_module.video_signal_controller.n3376\ : std_logic;
signal \transmit_module.old_VGA_HS\ : std_logic;
signal \ADV_HSYNC_c\ : std_logic;
signal \transmit_module.n188\ : std_logic;
signal \transmit_module.n3859\ : std_logic;
signal \transmit_module.TX_ADDR_1\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_1\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_11\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_12\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_13\ : std_logic;
signal \transmit_module.TX_ADDR_0\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_0\ : std_logic;
signal \transmit_module.TX_ADDR_5\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_5\ : std_logic;
signal \transmit_module.TX_ADDR_6\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_6\ : std_logic;
signal \transmit_module.TX_ADDR_2\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_2\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_7\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_4\ : std_logic;
signal \transmit_module.n184_cascade_\ : std_logic;
signal \transmit_module.n200\ : std_logic;
signal \transmit_module.TX_ADDR_4\ : std_logic;
signal \transmit_module.n197\ : std_logic;
signal \transmit_module.n213_cascade_\ : std_logic;
signal \transmit_module.TX_ADDR_7\ : std_logic;
signal \transmit_module.n184\ : std_logic;
signal \transmit_module.n216\ : std_logic;
signal n24 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_9\ : std_logic;
signal \transmit_module.n181\ : std_logic;
signal \transmit_module.n213\ : std_logic;
signal n21 : std_logic;
signal \line_buffer.n509\ : std_logic;
signal \line_buffer.n501\ : std_logic;
signal \line_buffer.n3770\ : std_logic;
signal \line_buffer.n571\ : std_logic;
signal \line_buffer.n563\ : std_logic;
signal \receive_module.rx_counter.n11\ : std_logic;
signal \LED_c\ : std_logic;
signal \receive_module.rx_counter.n3862\ : std_logic;
signal \TVP_VSYNC_c\ : std_logic;
signal \receive_module.BRAM_ADDR_13__N_31\ : std_logic;
signal \transmit_module.video_signal_controller.n2030\ : std_logic;
signal \transmit_module.video_signal_controller.n2551\ : std_logic;
signal \DEBUG_c_6\ : std_logic;
signal \transmit_module.video_signal_controller.SYNC_BUFF1\ : std_logic;
signal \transmit_module.video_signal_controller.SYNC_BUFF2\ : std_logic;
signal n3852 : std_logic;
signal \transmit_module.n2039\ : std_logic;
signal \line_buffer.n603\ : std_logic;
signal \line_buffer.n595\ : std_logic;
signal \line_buffer.n569\ : std_logic;
signal \line_buffer.n561\ : std_logic;
signal \line_buffer.n3830_cascade_\ : std_logic;
signal \TX_DATA_1\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_11\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_10\ : std_logic;
signal \transmit_module.video_signal_controller.n3858\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_38\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_35\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_37\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_36\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_40\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_39\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_34\ : std_logic;
signal \transmit_module.n3865\ : std_logic;
signal \line_buffer.n570\ : std_logic;
signal \line_buffer.n562\ : std_logic;
signal \line_buffer.n3705\ : std_logic;
signal \line_buffer.n3715\ : std_logic;
signal \line_buffer.n3773_cascade_\ : std_logic;
signal \TX_DATA_3\ : std_logic;
signal \line_buffer.n594\ : std_logic;
signal \line_buffer.n602\ : std_logic;
signal \line_buffer.n497\ : std_logic;
signal \line_buffer.n3803_cascade_\ : std_logic;
signal \line_buffer.n505\ : std_logic;
signal \line_buffer.n3806_cascade_\ : std_logic;
signal \line_buffer.n3782\ : std_logic;
signal \TX_DATA_2\ : std_logic;
signal \line_buffer.n635\ : std_logic;
signal \line_buffer.n627\ : std_logic;
signal \line_buffer.n3706\ : std_logic;
signal \line_buffer.n626\ : std_logic;
signal \line_buffer.n634\ : std_logic;
signal \line_buffer.n3779\ : std_logic;
signal \line_buffer.n3703\ : std_logic;
signal \line_buffer.n3791_cascade_\ : std_logic;
signal \TX_DATA_7\ : std_logic;
signal \line_buffer.n575\ : std_logic;
signal \line_buffer.n567\ : std_logic;
signal \line_buffer.n3702\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_3\ : std_logic;
signal \transmit_module.n2321\ : std_logic;
signal \line_buffer.n625\ : std_logic;
signal \line_buffer.n633\ : std_logic;
signal \line_buffer.n3827\ : std_logic;
signal \line_buffer.n598\ : std_logic;
signal \line_buffer.n606\ : std_logic;
signal \line_buffer.n3767\ : std_logic;
signal \line_buffer.n506\ : std_logic;
signal \line_buffer.n498\ : std_logic;
signal \line_buffer.n3714\ : std_logic;
signal \line_buffer.n510\ : std_logic;
signal \line_buffer.n502\ : std_logic;
signal \line_buffer.n3717\ : std_logic;
signal \receive_module.rx_counter.n3547_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3547\ : std_logic;
signal \receive_module.rx_counter.n3646_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3613\ : std_logic;
signal \receive_module.rx_counter.n28\ : std_logic;
signal \line_buffer.n629\ : std_logic;
signal \line_buffer.n637\ : std_logic;
signal \line_buffer.n565\ : std_logic;
signal \line_buffer.n3761_cascade_\ : std_logic;
signal \line_buffer.n573\ : std_logic;
signal \line_buffer.n3764\ : std_logic;
signal \TX_DATA_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_33\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_32\ : std_logic;
signal \transmit_module.n3864\ : std_logic;
signal \line_buffer.n607\ : std_logic;
signal \line_buffer.n599\ : std_logic;
signal \line_buffer.n3718\ : std_logic;
signal \transmit_module.n194\ : std_logic;
signal \transmit_module.n210_cascade_\ : std_logic;
signal \transmit_module.n201\ : std_logic;
signal \transmit_module.n217_cascade_\ : std_logic;
signal \transmit_module.TX_ADDR_3\ : std_logic;
signal \transmit_module.n3855\ : std_logic;
signal \transmit_module.n195\ : std_logic;
signal \transmit_module.TX_ADDR_9\ : std_logic;
signal \transmit_module.n3549\ : std_logic;
signal \transmit_module.n217\ : std_logic;
signal \transmit_module.n185\ : std_logic;
signal n25 : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_10\ : std_logic;
signal \transmit_module.TX_ADDR_10\ : std_logic;
signal \transmit_module.n178\ : std_logic;
signal \transmit_module.n210\ : std_logic;
signal \transmit_module.n178_cascade_\ : std_logic;
signal n18 : std_logic;
signal \GB_BUFFER_TVP_CLK_c_THRU_CO\ : std_logic;
signal \TVP_HSYNC_c\ : std_logic;
signal \receive_module.rx_counter.n10\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \receive_module.rx_counter.n9\ : std_logic;
signal \receive_module.rx_counter.n3357\ : std_logic;
signal \receive_module.rx_counter.n8\ : std_logic;
signal \receive_module.rx_counter.n3358\ : std_logic;
signal \receive_module.rx_counter.X_3\ : std_logic;
signal \receive_module.rx_counter.n3359\ : std_logic;
signal \receive_module.rx_counter.X_4\ : std_logic;
signal \receive_module.rx_counter.n3360\ : std_logic;
signal \receive_module.rx_counter.X_5\ : std_logic;
signal \receive_module.rx_counter.n3361\ : std_logic;
signal \receive_module.rx_counter.X_6\ : std_logic;
signal \receive_module.rx_counter.n3362\ : std_logic;
signal \receive_module.rx_counter.X_7\ : std_logic;
signal \receive_module.rx_counter.n3363\ : std_logic;
signal \receive_module.rx_counter.n3364\ : std_logic;
signal \receive_module.rx_counter.X_8\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \receive_module.rx_counter.n3365\ : std_logic;
signal \receive_module.rx_counter.X_9\ : std_logic;
signal \TVP_CLK_c\ : std_logic;
signal n3860 : std_logic;
signal \line_buffer.n597\ : std_logic;
signal \line_buffer.n605\ : std_logic;
signal \line_buffer.n604\ : std_logic;
signal \line_buffer.n596\ : std_logic;
signal \line_buffer.n508\ : std_logic;
signal \line_buffer.n3833\ : std_logic;
signal \line_buffer.n500\ : std_logic;
signal \line_buffer.n3836\ : std_logic;
signal \line_buffer.n3721\ : std_logic;
signal \TX_DATA_4\ : std_logic;
signal \transmit_module.n179\ : std_logic;
signal \transmit_module.n211\ : std_logic;
signal \ADV_VSYNC_c\ : std_logic;
signal \transmit_module.n3853\ : std_logic;
signal n19 : std_logic;
signal \line_buffer.n507\ : std_logic;
signal \line_buffer.n499\ : std_logic;
signal \line_buffer.n3720\ : std_logic;
signal \line_buffer.n592\ : std_logic;
signal \line_buffer.n600\ : std_logic;
signal \line_buffer.n572\ : std_logic;
signal \line_buffer.n564\ : std_logic;
signal \line_buffer.n503\ : std_logic;
signal \line_buffer.n3815\ : std_logic;
signal \line_buffer.n495\ : std_logic;
signal \line_buffer.n568\ : std_logic;
signal \line_buffer.n560\ : std_logic;
signal \line_buffer.n3824_cascade_\ : std_logic;
signal \line_buffer.n3818\ : std_logic;
signal \TX_DATA_0\ : std_logic;
signal \ADV_CLK_c\ : std_logic;
signal \line_buffer.n3699\ : std_logic;
signal \DEBUG_c_2\ : std_logic;
signal \line_buffer.n3797\ : std_logic;
signal \line_buffer.n636\ : std_logic;
signal \line_buffer.n628\ : std_logic;
signal \line_buffer.n3700\ : std_logic;
signal \line_buffer.n624\ : std_logic;
signal \line_buffer.n632\ : std_logic;
signal \line_buffer.n3821\ : std_logic;
signal \line_buffer.n593\ : std_logic;
signal \line_buffer.n601\ : std_logic;
signal \TX_ADDR_11\ : std_logic;
signal \TX_ADDR_12\ : std_logic;
signal \line_buffer.n496\ : std_logic;
signal \line_buffer.n3809_cascade_\ : std_logic;
signal \line_buffer.n504\ : std_logic;
signal \line_buffer.n3812\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \TVP_CLK_wire\ : std_logic;
signal \ADV_CLK_wire\ : std_logic;
signal \TVP_VIDEO_wire\ : std_logic_vector(9 downto 0);
signal \ADV_G_wire\ : std_logic_vector(7 downto 0);
signal \ADV_R_wire\ : std_logic_vector(7 downto 0);
signal \ADV_B_wire\ : std_logic_vector(7 downto 0);
signal \ADV_SYNC_N_wire\ : std_logic;
signal \TVP_HSYNC_wire\ : std_logic;
signal \TVP_VSYNC_wire\ : std_logic;
signal \ADV_BLANK_N_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \ADV_HSYNC_wire\ : std_logic;
signal \ADV_VSYNC_wire\ : std_logic;
signal \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \line_buffer.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \TVP_CLK_wire\ <= TVP_CLK;
    ADV_CLK <= \ADV_CLK_wire\;
    \TVP_VIDEO_wire\ <= TVP_VIDEO;
    ADV_G <= \ADV_G_wire\;
    ADV_R <= \ADV_R_wire\;
    ADV_B <= \ADV_B_wire\;
    ADV_SYNC_N <= \ADV_SYNC_N_wire\;
    \TVP_HSYNC_wire\ <= TVP_HSYNC;
    \TVP_VSYNC_wire\ <= TVP_VSYNC;
    ADV_BLANK_N <= \ADV_BLANK_N_wire\;
    LED <= \LED_wire\;
    ADV_HSYNC <= \ADV_HSYNC_wire\;
    ADV_VSYNC <= \ADV_VSYNC_wire\;
    \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.n510\ <= \line_buffer.mem2_physical_RDATA_wire\(11);
    \line_buffer.n509\ <= \line_buffer.mem2_physical_RDATA_wire\(3);
    \line_buffer.mem2_physical_RADDR_wire\ <= \N__18946\&\N__19984\&\N__10507\&\N__16900\&\N__9670\&\N__10279\&\N__17137\&\N__19336\&\N__12127\&\N__11581\&\N__11806\;
    \line_buffer.mem2_physical_WADDR_wire\ <= \N__16030\&\N__13693\&\N__13948\&\N__14203\&\N__14437\&\N__14698\&\N__14926\&\N__15193\&\N__15454\&\N__13090\&\N__13324\;
    \line_buffer.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8493\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8636\&'0'&'0'&'0';
    \line_buffer.n597\ <= \line_buffer.mem14_physical_RDATA_wire\(11);
    \line_buffer.n596\ <= \line_buffer.mem14_physical_RDATA_wire\(3);
    \line_buffer.mem14_physical_RADDR_wire\ <= \N__19018\&\N__20056\&\N__10579\&\N__16972\&\N__9742\&\N__10351\&\N__17209\&\N__19408\&\N__12199\&\N__11653\&\N__11878\;
    \line_buffer.mem14_physical_WADDR_wire\ <= \N__16102\&\N__13765\&\N__14020\&\N__14275\&\N__14509\&\N__14770\&\N__14998\&\N__15265\&\N__15526\&\N__13162\&\N__13396\;
    \line_buffer.mem14_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem14_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8421\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8291\&'0'&'0'&'0';
    \line_buffer.n607\ <= \line_buffer.mem5_physical_RDATA_wire\(11);
    \line_buffer.n606\ <= \line_buffer.mem5_physical_RDATA_wire\(3);
    \line_buffer.mem5_physical_RADDR_wire\ <= \N__18949\&\N__19999\&\N__10510\&\N__16909\&\N__9679\&\N__10288\&\N__17146\&\N__19345\&\N__12130\&\N__11596\&\N__11827\;
    \line_buffer.mem5_physical_WADDR_wire\ <= \N__16045\&\N__13708\&\N__13969\&\N__14212\&\N__14452\&\N__14695\&\N__14953\&\N__15208\&\N__15463\&\N__13099\&\N__13357\;
    \line_buffer.mem5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8520\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8637\&'0'&'0'&'0';
    \line_buffer.n565\ <= \line_buffer.mem11_physical_RDATA_wire\(11);
    \line_buffer.n564\ <= \line_buffer.mem11_physical_RDATA_wire\(3);
    \line_buffer.mem11_physical_RADDR_wire\ <= \N__19054\&\N__20092\&\N__10615\&\N__17008\&\N__9778\&\N__10387\&\N__17245\&\N__19444\&\N__12235\&\N__11689\&\N__11914\;
    \line_buffer.mem11_physical_WADDR_wire\ <= \N__16138\&\N__13801\&\N__14056\&\N__14311\&\N__14545\&\N__14806\&\N__15034\&\N__15301\&\N__15562\&\N__13198\&\N__13432\;
    \line_buffer.mem11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem11_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8381\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8270\&'0'&'0'&'0';
    \line_buffer.n627\ <= \line_buffer.mem21_physical_RDATA_wire\(11);
    \line_buffer.n626\ <= \line_buffer.mem21_physical_RDATA_wire\(3);
    \line_buffer.mem21_physical_RADDR_wire\ <= \N__18922\&\N__19960\&\N__10483\&\N__16876\&\N__9646\&\N__10255\&\N__17113\&\N__19312\&\N__12103\&\N__11557\&\N__11782\;
    \line_buffer.mem21_physical_WADDR_wire\ <= \N__16006\&\N__13669\&\N__13924\&\N__14179\&\N__14413\&\N__14674\&\N__14902\&\N__15169\&\N__15430\&\N__13066\&\N__13300\;
    \line_buffer.mem21_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem21_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8210\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8108\&'0'&'0'&'0';
    \line_buffer.n563\ <= \line_buffer.mem12_physical_RDATA_wire\(11);
    \line_buffer.n562\ <= \line_buffer.mem12_physical_RDATA_wire\(3);
    \line_buffer.mem12_physical_RADDR_wire\ <= \N__19042\&\N__20080\&\N__10603\&\N__16996\&\N__9766\&\N__10375\&\N__17233\&\N__19432\&\N__12223\&\N__11677\&\N__11902\;
    \line_buffer.mem12_physical_WADDR_wire\ <= \N__16126\&\N__13789\&\N__14044\&\N__14299\&\N__14533\&\N__14794\&\N__15022\&\N__15289\&\N__15550\&\N__13186\&\N__13420\;
    \line_buffer.mem12_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem12_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8167\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8100\&'0'&'0'&'0';
    \line_buffer.n506\ <= \line_buffer.mem18_physical_RDATA_wire\(11);
    \line_buffer.n505\ <= \line_buffer.mem18_physical_RDATA_wire\(3);
    \line_buffer.mem18_physical_RADDR_wire\ <= \N__18970\&\N__20008\&\N__10531\&\N__16924\&\N__9694\&\N__10303\&\N__17161\&\N__19360\&\N__12151\&\N__11605\&\N__11830\;
    \line_buffer.mem18_physical_WADDR_wire\ <= \N__16054\&\N__13717\&\N__13972\&\N__14227\&\N__14461\&\N__14722\&\N__14950\&\N__15217\&\N__15478\&\N__13114\&\N__13348\;
    \line_buffer.mem18_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem18_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8199\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8101\&'0'&'0'&'0';
    \line_buffer.n571\ <= \line_buffer.mem24_physical_RDATA_wire\(11);
    \line_buffer.n570\ <= \line_buffer.mem24_physical_RDATA_wire\(3);
    \line_buffer.mem24_physical_RADDR_wire\ <= \N__19069\&\N__20119\&\N__10630\&\N__17029\&\N__9799\&\N__10408\&\N__17266\&\N__19465\&\N__12250\&\N__11716\&\N__11947\;
    \line_buffer.mem24_physical_WADDR_wire\ <= \N__16165\&\N__13828\&\N__14089\&\N__14332\&\N__14572\&\N__14815\&\N__15071\&\N__15328\&\N__15583\&\N__13219\&\N__13472\;
    \line_buffer.mem24_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem24_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8136\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8025\&'0'&'0'&'0';
    \line_buffer.n599\ <= \line_buffer.mem1_physical_RDATA_wire\(11);
    \line_buffer.n598\ <= \line_buffer.mem1_physical_RDATA_wire\(3);
    \line_buffer.mem1_physical_RADDR_wire\ <= \N__19078\&\N__20116\&\N__10639\&\N__17032\&\N__9802\&\N__10411\&\N__17269\&\N__19468\&\N__12259\&\N__11713\&\N__11938\;
    \line_buffer.mem1_physical_WADDR_wire\ <= \N__16162\&\N__13825\&\N__14080\&\N__14335\&\N__14569\&\N__14828\&\N__15058\&\N__15325\&\N__15586\&\N__13222\&\N__13456\;
    \line_buffer.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8474\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8600\&'0'&'0'&'0';
    \line_buffer.n595\ <= \line_buffer.mem15_physical_RDATA_wire\(11);
    \line_buffer.n594\ <= \line_buffer.mem15_physical_RDATA_wire\(3);
    \line_buffer.mem15_physical_RADDR_wire\ <= \N__19006\&\N__20044\&\N__10567\&\N__16960\&\N__9730\&\N__10339\&\N__17197\&\N__19396\&\N__12187\&\N__11641\&\N__11866\;
    \line_buffer.mem15_physical_WADDR_wire\ <= \N__16090\&\N__13753\&\N__14008\&\N__14263\&\N__14497\&\N__14758\&\N__14986\&\N__15253\&\N__15514\&\N__13150\&\N__13384\;
    \line_buffer.mem15_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem15_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8180\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8092\&'0'&'0'&'0';
    \line_buffer.n603\ <= \line_buffer.mem27_physical_RDATA_wire\(11);
    \line_buffer.n602\ <= \line_buffer.mem27_physical_RDATA_wire\(3);
    \line_buffer.mem27_physical_RADDR_wire\ <= \N__19033\&\N__20083\&\N__10594\&\N__16993\&\N__9763\&\N__10372\&\N__17230\&\N__19429\&\N__12214\&\N__11680\&\N__11911\;
    \line_buffer.mem27_physical_WADDR_wire\ <= \N__16129\&\N__13792\&\N__14053\&\N__14296\&\N__14536\&\N__14779\&\N__15037\&\N__15292\&\N__15547\&\N__13183\&\N__13441\;
    \line_buffer.mem27_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem27_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8161\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8056\&'0'&'0'&'0';
    \line_buffer.n575\ <= \line_buffer.mem4_physical_RDATA_wire\(11);
    \line_buffer.n574\ <= \line_buffer.mem4_physical_RDATA_wire\(3);
    \line_buffer.mem4_physical_RADDR_wire\ <= \N__18961\&\N__20011\&\N__10522\&\N__16921\&\N__9691\&\N__10300\&\N__17158\&\N__19357\&\N__12142\&\N__11608\&\N__11839\;
    \line_buffer.mem4_physical_WADDR_wire\ <= \N__16057\&\N__13720\&\N__13981\&\N__14224\&\N__14464\&\N__14707\&\N__14965\&\N__15220\&\N__15475\&\N__13111\&\N__13369\;
    \line_buffer.mem4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8499\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8626\&'0'&'0'&'0';
    \line_buffer.n593\ <= \line_buffer.mem16_physical_RDATA_wire\(11);
    \line_buffer.n592\ <= \line_buffer.mem16_physical_RDATA_wire\(3);
    \line_buffer.mem16_physical_RADDR_wire\ <= \N__18994\&\N__20032\&\N__10555\&\N__16948\&\N__9718\&\N__10327\&\N__17185\&\N__19384\&\N__12175\&\N__11629\&\N__11854\;
    \line_buffer.mem16_physical_WADDR_wire\ <= \N__16078\&\N__13741\&\N__13996\&\N__14251\&\N__14485\&\N__14746\&\N__14974\&\N__15241\&\N__15502\&\N__13138\&\N__13372\;
    \line_buffer.mem16_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem16_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7962\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8758\&'0'&'0'&'0';
    \line_buffer.n635\ <= \line_buffer.mem30_physical_RDATA_wire\(11);
    \line_buffer.n634\ <= \line_buffer.mem30_physical_RDATA_wire\(3);
    \line_buffer.mem30_physical_RADDR_wire\ <= \N__18985\&\N__20035\&\N__10546\&\N__16945\&\N__9715\&\N__10324\&\N__17182\&\N__19381\&\N__12166\&\N__11632\&\N__11863\;
    \line_buffer.mem30_physical_WADDR_wire\ <= \N__16081\&\N__13744\&\N__14005\&\N__14248\&\N__14488\&\N__14731\&\N__14989\&\N__15244\&\N__15499\&\N__13135\&\N__13393\;
    \line_buffer.mem30_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem30_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8186\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8088\&'0'&'0'&'0';
    \line_buffer.n502\ <= \line_buffer.mem7_physical_RDATA_wire\(11);
    \line_buffer.n501\ <= \line_buffer.mem7_physical_RDATA_wire\(3);
    \line_buffer.mem7_physical_RADDR_wire\ <= \N__18925\&\N__19975\&\N__10486\&\N__16885\&\N__9655\&\N__10264\&\N__17122\&\N__19321\&\N__12106\&\N__11572\&\N__11803\;
    \line_buffer.mem7_physical_WADDR_wire\ <= \N__16021\&\N__13684\&\N__13945\&\N__14188\&\N__14428\&\N__14671\&\N__14929\&\N__15184\&\N__15439\&\N__13075\&\N__13333\;
    \line_buffer.mem7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem7_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8528\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8642\&'0'&'0'&'0';
    \line_buffer.n629\ <= \line_buffer.mem20_physical_RDATA_wire\(11);
    \line_buffer.n628\ <= \line_buffer.mem20_physical_RDATA_wire\(3);
    \line_buffer.mem20_physical_RADDR_wire\ <= \N__18934\&\N__19972\&\N__10495\&\N__16888\&\N__9658\&\N__10267\&\N__17125\&\N__19324\&\N__12115\&\N__11569\&\N__11794\;
    \line_buffer.mem20_physical_WADDR_wire\ <= \N__16018\&\N__13681\&\N__13936\&\N__14191\&\N__14425\&\N__14686\&\N__14914\&\N__15181\&\N__15442\&\N__13078\&\N__13312\;
    \line_buffer.mem20_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem20_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8420\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8312\&'0'&'0'&'0';
    \line_buffer.n561\ <= \line_buffer.mem13_physical_RDATA_wire\(11);
    \line_buffer.n560\ <= \line_buffer.mem13_physical_RDATA_wire\(3);
    \line_buffer.mem13_physical_RADDR_wire\ <= \N__19030\&\N__20068\&\N__10591\&\N__16984\&\N__9754\&\N__10363\&\N__17221\&\N__19420\&\N__12211\&\N__11665\&\N__11890\;
    \line_buffer.mem13_physical_WADDR_wire\ <= \N__16114\&\N__13777\&\N__14032\&\N__14287\&\N__14521\&\N__14782\&\N__15010\&\N__15277\&\N__15538\&\N__13174\&\N__13408\;
    \line_buffer.mem13_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem13_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7947\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8751\&'0'&'0'&'0';
    \line_buffer.n504\ <= \line_buffer.mem19_physical_RDATA_wire\(11);
    \line_buffer.n503\ <= \line_buffer.mem19_physical_RDATA_wire\(3);
    \line_buffer.mem19_physical_RADDR_wire\ <= \N__18958\&\N__19996\&\N__10519\&\N__16912\&\N__9682\&\N__10291\&\N__17149\&\N__19348\&\N__12139\&\N__11593\&\N__11818\;
    \line_buffer.mem19_physical_WADDR_wire\ <= \N__16042\&\N__13705\&\N__13960\&\N__14215\&\N__14449\&\N__14710\&\N__14938\&\N__15205\&\N__15466\&\N__13102\&\N__13336\;
    \line_buffer.mem19_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem19_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7969\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8770\&'0'&'0'&'0';
    \line_buffer.n573\ <= \line_buffer.mem23_physical_RDATA_wire\(11);
    \line_buffer.n572\ <= \line_buffer.mem23_physical_RDATA_wire\(3);
    \line_buffer.mem23_physical_RADDR_wire\ <= \N__19081\&\N__20129\&\N__10642\&\N__17041\&\N__9811\&\N__10420\&\N__17278\&\N__19477\&\N__12262\&\N__11726\&\N__11954\;
    \line_buffer.mem23_physical_WADDR_wire\ <= \N__16175\&\N__13838\&\N__14096\&\N__14344\&\N__14582\&\N__14827\&\N__15077\&\N__15338\&\N__15595\&\N__13231\&\N__13478\;
    \line_buffer.mem23_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem23_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8397\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8238\&'0'&'0'&'0';
    \line_buffer.n567\ <= \line_buffer.mem0_physical_RDATA_wire\(11);
    \line_buffer.n566\ <= \line_buffer.mem0_physical_RDATA_wire\(3);
    \line_buffer.mem0_physical_RADDR_wire\ <= \N__19085\&\N__20128\&\N__10646\&\N__17042\&\N__9812\&\N__10421\&\N__17279\&\N__19478\&\N__12266\&\N__11725\&\N__11950\;
    \line_buffer.mem0_physical_WADDR_wire\ <= \N__16174\&\N__13837\&\N__14092\&\N__14345\&\N__14581\&\N__14834\&\N__15070\&\N__15337\&\N__15596\&\N__13232\&\N__13468\;
    \line_buffer.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8449\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8599\&'0'&'0'&'0';
    \line_buffer.n605\ <= \line_buffer.mem26_physical_RDATA_wire\(11);
    \line_buffer.n604\ <= \line_buffer.mem26_physical_RDATA_wire\(3);
    \line_buffer.mem26_physical_RADDR_wire\ <= \N__19045\&\N__20095\&\N__10606\&\N__17005\&\N__9775\&\N__10384\&\N__17242\&\N__19441\&\N__12226\&\N__11692\&\N__11923\;
    \line_buffer.mem26_physical_WADDR_wire\ <= \N__16141\&\N__13804\&\N__14065\&\N__14308\&\N__14548\&\N__14791\&\N__15049\&\N__15304\&\N__15559\&\N__13195\&\N__13453\;
    \line_buffer.mem26_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem26_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8380\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8263\&'0'&'0'&'0';
    \line_buffer.n631\ <= \line_buffer.mem3_physical_RDATA_wire\(11);
    \line_buffer.n630\ <= \line_buffer.mem3_physical_RDATA_wire\(3);
    \line_buffer.mem3_physical_RADDR_wire\ <= \N__18997\&\N__20047\&\N__10558\&\N__16957\&\N__9727\&\N__10336\&\N__17194\&\N__19393\&\N__12178\&\N__11644\&\N__11875\;
    \line_buffer.mem3_physical_WADDR_wire\ <= \N__16093\&\N__13756\&\N__14017\&\N__14260\&\N__14500\&\N__14743\&\N__15001\&\N__15256\&\N__15511\&\N__13147\&\N__13405\;
    \line_buffer.mem3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8506\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8612\&'0'&'0'&'0';
    \line_buffer.n508\ <= \line_buffer.mem17_physical_RDATA_wire\(11);
    \line_buffer.n507\ <= \line_buffer.mem17_physical_RDATA_wire\(3);
    \line_buffer.mem17_physical_RADDR_wire\ <= \N__18982\&\N__20020\&\N__10543\&\N__16936\&\N__9706\&\N__10315\&\N__17173\&\N__19372\&\N__12163\&\N__11617\&\N__11842\;
    \line_buffer.mem17_physical_WADDR_wire\ <= \N__16066\&\N__13729\&\N__13984\&\N__14239\&\N__14473\&\N__14734\&\N__14962\&\N__15229\&\N__15490\&\N__13126\&\N__13360\;
    \line_buffer.mem17_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem17_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8404\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8301\&'0'&'0'&'0';
    \line_buffer.n633\ <= \line_buffer.mem31_physical_RDATA_wire\(11);
    \line_buffer.n632\ <= \line_buffer.mem31_physical_RDATA_wire\(3);
    \line_buffer.mem31_physical_RADDR_wire\ <= \N__18973\&\N__20023\&\N__10534\&\N__16933\&\N__9703\&\N__10312\&\N__17170\&\N__19369\&\N__12154\&\N__11620\&\N__11851\;
    \line_buffer.mem31_physical_WADDR_wire\ <= \N__16069\&\N__13732\&\N__13993\&\N__14236\&\N__14476\&\N__14719\&\N__14977\&\N__15232\&\N__15487\&\N__13123\&\N__13381\;
    \line_buffer.mem31_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem31_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7929\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8736\&'0'&'0'&'0';
    \line_buffer.n498\ <= \line_buffer.mem9_physical_RDATA_wire\(11);
    \line_buffer.n497\ <= \line_buffer.mem9_physical_RDATA_wire\(3);
    \line_buffer.mem9_physical_RADDR_wire\ <= \N__18901\&\N__19951\&\N__10462\&\N__16861\&\N__9631\&\N__10240\&\N__17098\&\N__19297\&\N__12082\&\N__11548\&\N__11779\;
    \line_buffer.mem9_physical_WADDR_wire\ <= \N__15997\&\N__13660\&\N__13921\&\N__14164\&\N__14404\&\N__14647\&\N__14905\&\N__15160\&\N__15415\&\N__13051\&\N__13309\;
    \line_buffer.mem9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem9_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8209\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8099\&'0'&'0'&'0';
    \line_buffer.n637\ <= \line_buffer.mem29_physical_RDATA_wire\(11);
    \line_buffer.n636\ <= \line_buffer.mem29_physical_RDATA_wire\(3);
    \line_buffer.mem29_physical_RADDR_wire\ <= \N__19009\&\N__20059\&\N__10570\&\N__16969\&\N__9739\&\N__10348\&\N__17206\&\N__19405\&\N__12190\&\N__11656\&\N__11887\;
    \line_buffer.mem29_physical_WADDR_wire\ <= \N__16105\&\N__13768\&\N__14029\&\N__14272\&\N__14512\&\N__14755\&\N__15013\&\N__15268\&\N__15523\&\N__13159\&\N__13417\;
    \line_buffer.mem29_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem29_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8422\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8276\&'0'&'0'&'0';
    \line_buffer.n639\ <= \line_buffer.mem6_physical_RDATA_wire\(11);
    \line_buffer.n638\ <= \line_buffer.mem6_physical_RDATA_wire\(3);
    \line_buffer.mem6_physical_RADDR_wire\ <= \N__18937\&\N__19987\&\N__10498\&\N__16897\&\N__9667\&\N__10276\&\N__17134\&\N__19333\&\N__12118\&\N__11584\&\N__11815\;
    \line_buffer.mem6_physical_WADDR_wire\ <= \N__16033\&\N__13696\&\N__13957\&\N__14200\&\N__14440\&\N__14683\&\N__14941\&\N__15196\&\N__15451\&\N__13087\&\N__13345\;
    \line_buffer.mem6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8527\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8638\&'0'&'0'&'0';
    \line_buffer.n496\ <= \line_buffer.mem10_physical_RDATA_wire\(11);
    \line_buffer.n495\ <= \line_buffer.mem10_physical_RDATA_wire\(3);
    \line_buffer.mem10_physical_RADDR_wire\ <= \N__19066\&\N__20104\&\N__10627\&\N__17020\&\N__9790\&\N__10399\&\N__17257\&\N__19456\&\N__12247\&\N__11701\&\N__11926\;
    \line_buffer.mem10_physical_WADDR_wire\ <= \N__16150\&\N__13813\&\N__14068\&\N__14323\&\N__14557\&\N__14818\&\N__15046\&\N__15313\&\N__15574\&\N__13210\&\N__13444\;
    \line_buffer.mem10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem10_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7938\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8737\&'0'&'0'&'0';
    \line_buffer.n625\ <= \line_buffer.mem22_physical_RDATA_wire\(11);
    \line_buffer.n624\ <= \line_buffer.mem22_physical_RDATA_wire\(3);
    \line_buffer.mem22_physical_RADDR_wire\ <= \N__18910\&\N__19948\&\N__10471\&\N__16864\&\N__9634\&\N__10243\&\N__17101\&\N__19300\&\N__12091\&\N__11545\&\N__11770\;
    \line_buffer.mem22_physical_WADDR_wire\ <= \N__15994\&\N__13657\&\N__13912\&\N__14167\&\N__14401\&\N__14662\&\N__14890\&\N__15157\&\N__15418\&\N__13054\&\N__13288\;
    \line_buffer.mem22_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem22_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7976\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8777\&'0'&'0'&'0';
    \line_buffer.n569\ <= \line_buffer.mem25_physical_RDATA_wire\(11);
    \line_buffer.n568\ <= \line_buffer.mem25_physical_RDATA_wire\(3);
    \line_buffer.mem25_physical_RADDR_wire\ <= \N__19057\&\N__20107\&\N__10618\&\N__17017\&\N__9787\&\N__10396\&\N__17254\&\N__19453\&\N__12238\&\N__11704\&\N__11935\;
    \line_buffer.mem25_physical_WADDR_wire\ <= \N__16153\&\N__13816\&\N__14077\&\N__14320\&\N__14560\&\N__14803\&\N__15061\&\N__15316\&\N__15571\&\N__13207\&\N__13465\;
    \line_buffer.mem25_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem25_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7920\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8705\&'0'&'0'&'0';
    \line_buffer.n500\ <= \line_buffer.mem8_physical_RDATA_wire\(11);
    \line_buffer.n499\ <= \line_buffer.mem8_physical_RDATA_wire\(3);
    \line_buffer.mem8_physical_RADDR_wire\ <= \N__18913\&\N__19963\&\N__10474\&\N__16873\&\N__9643\&\N__10252\&\N__17110\&\N__19309\&\N__12094\&\N__11560\&\N__11791\;
    \line_buffer.mem8_physical_WADDR_wire\ <= \N__16009\&\N__13672\&\N__13933\&\N__14176\&\N__14416\&\N__14659\&\N__14917\&\N__15172\&\N__15427\&\N__13063\&\N__13321\;
    \line_buffer.mem8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem8_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8426\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8311\&'0'&'0'&'0';
    \line_buffer.n601\ <= \line_buffer.mem28_physical_RDATA_wire\(11);
    \line_buffer.n600\ <= \line_buffer.mem28_physical_RDATA_wire\(3);
    \line_buffer.mem28_physical_RADDR_wire\ <= \N__19021\&\N__20071\&\N__10582\&\N__16981\&\N__9751\&\N__10360\&\N__17218\&\N__19417\&\N__12202\&\N__11668\&\N__11899\;
    \line_buffer.mem28_physical_WADDR_wire\ <= \N__16117\&\N__13780\&\N__14041\&\N__14284\&\N__14524\&\N__14767\&\N__15025\&\N__15280\&\N__15535\&\N__13171\&\N__13429\;
    \line_buffer.mem28_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem28_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7919\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8718\&'0'&'0'&'0';

    \tx_pll.TX_PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0100110",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \ADV_CLK_c\,
            REFERENCECLK => \N__18875\,
            RESETB => \N__22507\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \line_buffer.mem2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem2_physical_RDATA_wire\,
            RADDR => \line_buffer.mem2_physical_RADDR_wire\,
            WADDR => \line_buffer.mem2_physical_WADDR_wire\,
            MASK => \line_buffer.mem2_physical_MASK_wire\,
            WDATA => \line_buffer.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21957\,
            RE => \N__22516\,
            WCLKE => 'H',
            WCLK => \N__21039\,
            WE => \N__10778\
        );

    \line_buffer.mem14_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem14_physical_RDATA_wire\,
            RADDR => \line_buffer.mem14_physical_RADDR_wire\,
            WADDR => \line_buffer.mem14_physical_WADDR_wire\,
            MASK => \line_buffer.mem14_physical_MASK_wire\,
            WDATA => \line_buffer.mem14_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22053\,
            RE => \N__22621\,
            WCLKE => 'H',
            WCLK => \N__21024\,
            WE => \N__10970\
        );

    \line_buffer.mem5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem5_physical_RDATA_wire\,
            RADDR => \line_buffer.mem5_physical_RADDR_wire\,
            WADDR => \line_buffer.mem5_physical_WADDR_wire\,
            MASK => \line_buffer.mem5_physical_MASK_wire\,
            WDATA => \line_buffer.mem5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21490\,
            RE => \N__22607\,
            WCLKE => 'H',
            WCLK => \N__21035\,
            WE => \N__9917\
        );

    \line_buffer.mem11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem11_physical_RDATA_wire\,
            RADDR => \line_buffer.mem11_physical_RADDR_wire\,
            WADDR => \line_buffer.mem11_physical_WADDR_wire\,
            MASK => \line_buffer.mem11_physical_MASK_wire\,
            WDATA => \line_buffer.mem11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22150\,
            RE => \N__22667\,
            WCLKE => 'H',
            WCLK => \N__21016\,
            WE => \N__10831\
        );

    \line_buffer.mem21_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem21_physical_RDATA_wire\,
            RADDR => \line_buffer.mem21_physical_RADDR_wire\,
            WADDR => \line_buffer.mem21_physical_WADDR_wire\,
            MASK => \line_buffer.mem21_physical_MASK_wire\,
            WDATA => \line_buffer.mem21_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21808\,
            RE => \N__22471\,
            WCLKE => 'H',
            WCLK => \N__21043\,
            WE => \N__11033\
        );

    \line_buffer.mem12_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem12_physical_RDATA_wire\,
            RADDR => \line_buffer.mem12_physical_RADDR_wire\,
            WADDR => \line_buffer.mem12_physical_WADDR_wire\,
            MASK => \line_buffer.mem12_physical_MASK_wire\,
            WDATA => \line_buffer.mem12_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22124\,
            RE => \N__22508\,
            WCLKE => 'H',
            WCLK => \N__21020\,
            WE => \N__10814\
        );

    \line_buffer.mem18_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem18_physical_RDATA_wire\,
            RADDR => \line_buffer.mem18_physical_RADDR_wire\,
            WADDR => \line_buffer.mem18_physical_WADDR_wire\,
            MASK => \line_buffer.mem18_physical_MASK_wire\,
            WDATA => \line_buffer.mem18_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21765\,
            RE => \N__22557\,
            WCLKE => 'H',
            WCLK => \N__21032\,
            WE => \N__10774\
        );

    \line_buffer.mem24_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem24_physical_RDATA_wire\,
            RADDR => \line_buffer.mem24_physical_RADDR_wire\,
            WADDR => \line_buffer.mem24_physical_WADDR_wire\,
            MASK => \line_buffer.mem24_physical_MASK_wire\,
            WDATA => \line_buffer.mem24_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21682\,
            RE => \N__22693\,
            WCLKE => 'H',
            WCLK => \N__21007\,
            WE => \N__9468\
        );

    \line_buffer.mem1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem1_physical_RDATA_wire\,
            RADDR => \line_buffer.mem1_physical_RADDR_wire\,
            WADDR => \line_buffer.mem1_physical_WADDR_wire\,
            MASK => \line_buffer.mem1_physical_MASK_wire\,
            WDATA => \line_buffer.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22159\,
            RE => \N__22684\,
            WCLKE => 'H',
            WCLK => \N__21004\,
            WE => \N__10977\
        );

    \line_buffer.mem15_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem15_physical_RDATA_wire\,
            RADDR => \line_buffer.mem15_physical_RADDR_wire\,
            WADDR => \line_buffer.mem15_physical_WADDR_wire\,
            MASK => \line_buffer.mem15_physical_MASK_wire\,
            WDATA => \line_buffer.mem15_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22052\,
            RE => \N__22620\,
            WCLKE => 'H',
            WCLK => \N__21026\,
            WE => \N__10978\
        );

    \line_buffer.mem27_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem27_physical_RDATA_wire\,
            RADDR => \line_buffer.mem27_physical_RADDR_wire\,
            WADDR => \line_buffer.mem27_physical_WADDR_wire\,
            MASK => \line_buffer.mem27_physical_MASK_wire\,
            WDATA => \line_buffer.mem27_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21959\,
            RE => \N__22672\,
            WCLKE => 'H',
            WCLK => \N__21021\,
            WE => \N__9896\
        );

    \line_buffer.mem4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem4_physical_RDATA_wire\,
            RADDR => \line_buffer.mem4_physical_RADDR_wire\,
            WADDR => \line_buffer.mem4_physical_WADDR_wire\,
            MASK => \line_buffer.mem4_physical_MASK_wire\,
            WDATA => \line_buffer.mem4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21723\,
            RE => \N__22608\,
            WCLKE => 'H',
            WCLK => \N__21033\,
            WE => \N__9476\
        );

    \line_buffer.mem16_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem16_physical_RDATA_wire\,
            RADDR => \line_buffer.mem16_physical_RADDR_wire\,
            WADDR => \line_buffer.mem16_physical_WADDR_wire\,
            MASK => \line_buffer.mem16_physical_MASK_wire\,
            WDATA => \line_buffer.mem16_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21926\,
            RE => \N__22592\,
            WCLKE => 'H',
            WCLK => \N__21028\,
            WE => \N__10979\
        );

    \line_buffer.mem30_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem30_physical_RDATA_wire\,
            RADDR => \line_buffer.mem30_physical_RADDR_wire\,
            WADDR => \line_buffer.mem30_physical_WADDR_wire\,
            MASK => \line_buffer.mem30_physical_MASK_wire\,
            WDATA => \line_buffer.mem30_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22089\,
            RE => \N__22590\,
            WCLKE => 'H',
            WCLK => \N__21029\,
            WE => \N__9507\
        );

    \line_buffer.mem7_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem7_physical_RDATA_wire\,
            RADDR => \line_buffer.mem7_physical_RADDR_wire\,
            WADDR => \line_buffer.mem7_physical_WADDR_wire\,
            MASK => \line_buffer.mem7_physical_MASK_wire\,
            WDATA => \line_buffer.mem7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21446\,
            RE => \N__22574\,
            WCLKE => 'H',
            WCLK => \N__21042\,
            WE => \N__9861\
        );

    \line_buffer.mem20_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem20_physical_RDATA_wire\,
            RADDR => \line_buffer.mem20_physical_RADDR_wire\,
            WADDR => \line_buffer.mem20_physical_WADDR_wire\,
            MASK => \line_buffer.mem20_physical_MASK_wire\,
            WDATA => \line_buffer.mem20_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21809\,
            RE => \N__22515\,
            WCLKE => 'H',
            WCLK => \N__21041\,
            WE => \N__11028\
        );

    \line_buffer.mem13_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem13_physical_RDATA_wire\,
            RADDR => \line_buffer.mem13_physical_RADDR_wire\,
            WADDR => \line_buffer.mem13_physical_WADDR_wire\,
            MASK => \line_buffer.mem13_physical_MASK_wire\,
            WDATA => \line_buffer.mem13_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22123\,
            RE => \N__22645\,
            WCLKE => 'H',
            WCLK => \N__21022\,
            WE => \N__10824\
        );

    \line_buffer.mem19_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem19_physical_RDATA_wire\,
            RADDR => \line_buffer.mem19_physical_RADDR_wire\,
            WADDR => \line_buffer.mem19_physical_WADDR_wire\,
            MASK => \line_buffer.mem19_physical_MASK_wire\,
            WDATA => \line_buffer.mem19_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21958\,
            RE => \N__22556\,
            WCLKE => 'H',
            WCLK => \N__21034\,
            WE => \N__10773\
        );

    \line_buffer.mem23_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem23_physical_RDATA_wire\,
            RADDR => \line_buffer.mem23_physical_RADDR_wire\,
            WADDR => \line_buffer.mem23_physical_WADDR_wire\,
            MASK => \line_buffer.mem23_physical_MASK_wire\,
            WDATA => \line_buffer.mem23_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22137\,
            RE => \N__22694\,
            WCLKE => 'H',
            WCLK => \N__21003\,
            WE => \N__9475\
        );

    \line_buffer.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem0_physical_RDATA_wire\,
            RADDR => \line_buffer.mem0_physical_RADDR_wire\,
            WADDR => \line_buffer.mem0_physical_WADDR_wire\,
            MASK => \line_buffer.mem0_physical_MASK_wire\,
            WDATA => \line_buffer.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22160\,
            RE => \N__22555\,
            WCLKE => 'H',
            WCLK => \N__21001\,
            WE => \N__10832\
        );

    \line_buffer.mem26_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem26_physical_RDATA_wire\,
            RADDR => \line_buffer.mem26_physical_RADDR_wire\,
            WADDR => \line_buffer.mem26_physical_WADDR_wire\,
            MASK => \line_buffer.mem26_physical_MASK_wire\,
            WDATA => \line_buffer.mem26_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22158\,
            RE => \N__22685\,
            WCLKE => 'H',
            WCLK => \N__21019\,
            WE => \N__9907\
        );

    \line_buffer.mem3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem3_physical_RDATA_wire\,
            RADDR => \line_buffer.mem3_physical_RADDR_wire\,
            WADDR => \line_buffer.mem3_physical_WADDR_wire\,
            MASK => \line_buffer.mem3_physical_MASK_wire\,
            WDATA => \line_buffer.mem3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21553\,
            RE => \N__22652\,
            WCLKE => 'H',
            WCLK => \N__21027\,
            WE => \N__11027\
        );

    \line_buffer.mem17_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem17_physical_RDATA_wire\,
            RADDR => \line_buffer.mem17_physical_RADDR_wire\,
            WADDR => \line_buffer.mem17_physical_WADDR_wire\,
            MASK => \line_buffer.mem17_physical_MASK_wire\,
            WDATA => \line_buffer.mem17_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21925\,
            RE => \N__22591\,
            WCLKE => 'H',
            WCLK => \N__21030\,
            WE => \N__10766\
        );

    \line_buffer.mem31_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem31_physical_RDATA_wire\,
            RADDR => \line_buffer.mem31_physical_RADDR_wire\,
            WADDR => \line_buffer.mem31_physical_WADDR_wire\,
            MASK => \line_buffer.mem31_physical_MASK_wire\,
            WDATA => \line_buffer.mem31_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22119\,
            RE => \N__22631\,
            WCLKE => 'H',
            WCLK => \N__21031\,
            WE => \N__9514\
        );

    \line_buffer.mem9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem9_physical_RDATA_wire\,
            RADDR => \line_buffer.mem9_physical_RADDR_wire\,
            WADDR => \line_buffer.mem9_physical_WADDR_wire\,
            MASK => \line_buffer.mem9_physical_MASK_wire\,
            WDATA => \line_buffer.mem9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21509\,
            RE => \N__22533\,
            WCLKE => 'H',
            WCLK => \N__21046\,
            WE => \N__9869\
        );

    \line_buffer.mem29_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem29_physical_RDATA_wire\,
            RADDR => \line_buffer.mem29_physical_RADDR_wire\,
            WADDR => \line_buffer.mem29_physical_WADDR_wire\,
            MASK => \line_buffer.mem29_physical_MASK_wire\,
            WDATA => \line_buffer.mem29_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21817\,
            RE => \N__22653\,
            WCLKE => 'H',
            WCLK => \N__21025\,
            WE => \N__9498\
        );

    \line_buffer.mem6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem6_physical_RDATA_wire\,
            RADDR => \line_buffer.mem6_physical_RADDR_wire\,
            WADDR => \line_buffer.mem6_physical_WADDR_wire\,
            MASK => \line_buffer.mem6_physical_MASK_wire\,
            WDATA => \line_buffer.mem6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21782\,
            RE => \N__22575\,
            WCLKE => 'H',
            WCLK => \N__21040\,
            WE => \N__9518\
        );

    \line_buffer.mem10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem10_physical_RDATA_wire\,
            RADDR => \line_buffer.mem10_physical_RADDR_wire\,
            WADDR => \line_buffer.mem10_physical_WADDR_wire\,
            MASK => \line_buffer.mem10_physical_MASK_wire\,
            WDATA => \line_buffer.mem10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22151\,
            RE => \N__22554\,
            WCLKE => 'H',
            WCLK => \N__21008\,
            WE => \N__9852\
        );

    \line_buffer.mem22_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem22_physical_RDATA_wire\,
            RADDR => \line_buffer.mem22_physical_RADDR_wire\,
            WADDR => \line_buffer.mem22_physical_WADDR_wire\,
            MASK => \line_buffer.mem22_physical_MASK_wire\,
            WDATA => \line_buffer.mem22_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21804\,
            RE => \N__22432\,
            WCLKE => 'H',
            WCLK => \N__21045\,
            WE => \N__11029\
        );

    \line_buffer.mem25_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem25_physical_RDATA_wire\,
            RADDR => \line_buffer.mem25_physical_RADDR_wire\,
            WADDR => \line_buffer.mem25_physical_WADDR_wire\,
            MASK => \line_buffer.mem25_physical_MASK_wire\,
            WDATA => \line_buffer.mem25_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22073\,
            RE => \N__22686\,
            WCLKE => 'H',
            WCLK => \N__21011\,
            WE => \N__9458\
        );

    \line_buffer.mem8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem8_physical_RDATA_wire\,
            RADDR => \line_buffer.mem8_physical_RADDR_wire\,
            WADDR => \line_buffer.mem8_physical_WADDR_wire\,
            MASK => \line_buffer.mem8_physical_MASK_wire\,
            WDATA => \line_buffer.mem8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21628\,
            RE => \N__22534\,
            WCLKE => 'H',
            WCLK => \N__21044\,
            WE => \N__9868\
        );

    \line_buffer.mem28_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem28_physical_RDATA_wire\,
            RADDR => \line_buffer.mem28_physical_RADDR_wire\,
            WADDR => \line_buffer.mem28_physical_WADDR_wire\,
            MASK => \line_buffer.mem28_physical_MASK_wire\,
            WDATA => \line_buffer.mem28_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22144\,
            RE => \N__22671\,
            WCLKE => 'H',
            WCLK => \N__21023\,
            WE => \N__9906\
        );

    \TVP_CLK_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__23673\,
            GLOBALBUFFEROUTPUT => \TVP_CLK_c\
        );

    \TVP_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23675\,
            DIN => \N__23674\,
            DOUT => \N__23673\,
            PACKAGEPIN => \TVP_CLK_wire\
        );

    \TVP_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23675\,
            PADOUT => \N__23674\,
            PADIN => \N__23673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23664\,
            DIN => \N__23663\,
            DOUT => \N__23662\,
            PACKAGEPIN => \ADV_CLK_wire\
        );

    \ADV_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23664\,
            PADOUT => \N__23663\,
            PADIN => \N__23662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21956\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23655\,
            DIN => \N__23654\,
            DOUT => \N__23653\,
            PACKAGEPIN => DEBUG(3)
        );

    \DEBUG_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23655\,
            PADOUT => \N__23654\,
            PADIN => \N__23653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15773\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23646\,
            DIN => \N__23645\,
            DOUT => \N__23644\,
            PACKAGEPIN => \TVP_VIDEO_wire\(2)
        );

    \TVP_VIDEO_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23646\,
            PADOUT => \N__23645\,
            PADIN => \N__23644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23637\,
            DIN => \N__23636\,
            DOUT => \N__23635\,
            PACKAGEPIN => \ADV_G_wire\(5)
        );

    \ADV_G_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23637\,
            PADOUT => \N__23636\,
            PADIN => \N__23635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12470\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23628\,
            DIN => \N__23627\,
            DOUT => \N__23626\,
            PACKAGEPIN => \ADV_R_wire\(3)
        );

    \ADV_R_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23628\,
            PADOUT => \N__23627\,
            PADIN => \N__23626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12579\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23619\,
            DIN => \N__23618\,
            DOUT => \N__23617\,
            PACKAGEPIN => \ADV_B_wire\(5)
        );

    \ADV_B_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23619\,
            PADOUT => \N__23618\,
            PADIN => \N__23617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12469\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23610\,
            DIN => \N__23609\,
            DOUT => \N__23608\,
            PACKAGEPIN => DEBUG(7)
        );

    \DEBUG_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23610\,
            PADOUT => \N__23609\,
            PADIN => \N__23608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23601\,
            DIN => \N__23600\,
            DOUT => \N__23599\,
            PACKAGEPIN => \TVP_VIDEO_wire\(6)
        );

    \TVP_VIDEO_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23601\,
            PADOUT => \N__23600\,
            PADIN => \N__23599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23592\,
            DIN => \N__23591\,
            DOUT => \N__23590\,
            PACKAGEPIN => \ADV_G_wire\(1)
        );

    \ADV_G_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23592\,
            PADOUT => \N__23591\,
            PADIN => \N__23590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11453\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23583\,
            DIN => \N__23582\,
            DOUT => \N__23581\,
            PACKAGEPIN => \ADV_R_wire\(0)
        );

    \ADV_R_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23583\,
            PADOUT => \N__23582\,
            PADIN => \N__23581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11506\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23574\,
            DIN => \N__23573\,
            DOUT => \N__23572\,
            PACKAGEPIN => DEBUG(2)
        );

    \DEBUG_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23574\,
            PADOUT => \N__23573\,
            PADIN => \N__23572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21296\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23565\,
            DIN => \N__23564\,
            DOUT => \N__23563\,
            PACKAGEPIN => \TVP_VIDEO_wire\(3)
        );

    \TVP_VIDEO_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23565\,
            PADOUT => \N__23564\,
            PADIN => \N__23563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23556\,
            DIN => \N__23555\,
            DOUT => \N__23554\,
            PACKAGEPIN => \ADV_G_wire\(4)
        );

    \ADV_G_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23556\,
            PADOUT => \N__23555\,
            PADIN => \N__23554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12516\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23547\,
            DIN => \N__23546\,
            DOUT => \N__23545\,
            PACKAGEPIN => \ADV_R_wire\(5)
        );

    \ADV_R_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23547\,
            PADOUT => \N__23546\,
            PADIN => \N__23545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12468\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23538\,
            DIN => \N__23537\,
            DOUT => \N__23536\,
            PACKAGEPIN => \TVP_VIDEO_wire\(9)
        );

    \TVP_VIDEO_pad_9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23538\,
            PADOUT => \N__23537\,
            PADIN => \N__23536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23529\,
            DIN => \N__23528\,
            DOUT => \N__23527\,
            PACKAGEPIN => DEBUG(1)
        );

    \DEBUG_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23529\,
            PADOUT => \N__23528\,
            PADIN => \N__23527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23520\,
            DIN => \N__23519\,
            DOUT => \N__23518\,
            PACKAGEPIN => \ADV_B_wire\(1)
        );

    \ADV_B_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23520\,
            PADOUT => \N__23519\,
            PADIN => \N__23518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11448\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_SYNC_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23511\,
            DIN => \N__23510\,
            DOUT => \N__23509\,
            PACKAGEPIN => \ADV_SYNC_N_wire\
        );

    \ADV_SYNC_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23511\,
            PADOUT => \N__23510\,
            PADIN => \N__23509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23502\,
            DIN => \N__23501\,
            DOUT => \N__23500\,
            PACKAGEPIN => \ADV_B_wire\(6)
        );

    \ADV_B_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23502\,
            PADOUT => \N__23501\,
            PADIN => \N__23500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12416\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23493\,
            DIN => \N__23492\,
            DOUT => \N__23491\,
            PACKAGEPIN => DEBUG(6)
        );

    \DEBUG_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23493\,
            PADOUT => \N__23492\,
            PADIN => \N__23491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17573\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23484\,
            DIN => \N__23483\,
            DOUT => \N__23482\,
            PACKAGEPIN => \TVP_VIDEO_wire\(7)
        );

    \TVP_VIDEO_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23484\,
            PADOUT => \N__23483\,
            PADIN => \N__23482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23475\,
            DIN => \N__23474\,
            DOUT => \N__23473\,
            PACKAGEPIN => \ADV_G_wire\(0)
        );

    \ADV_G_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23475\,
            PADOUT => \N__23474\,
            PADIN => \N__23473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11507\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23466\,
            DIN => \N__23465\,
            DOUT => \N__23464\,
            PACKAGEPIN => \ADV_R_wire\(1)
        );

    \ADV_R_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23466\,
            PADOUT => \N__23465\,
            PADIN => \N__23464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11449\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23457\,
            DIN => \N__23456\,
            DOUT => \N__23455\,
            PACKAGEPIN => DEBUG(5)
        );

    \DEBUG_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23457\,
            PADOUT => \N__23456\,
            PADIN => \N__23455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11333\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23448\,
            DIN => \N__23447\,
            DOUT => \N__23446\,
            PACKAGEPIN => \TVP_HSYNC_wire\
        );

    \TVP_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23448\,
            PADOUT => \N__23447\,
            PADIN => \N__23446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_HSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23439\,
            DIN => \N__23438\,
            DOUT => \N__23437\,
            PACKAGEPIN => \ADV_G_wire\(7)
        );

    \ADV_G_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23439\,
            PADOUT => \N__23438\,
            PADIN => \N__23437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12345\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23430\,
            DIN => \N__23429\,
            DOUT => \N__23428\,
            PACKAGEPIN => \ADV_R_wire\(6)
        );

    \ADV_R_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23430\,
            PADOUT => \N__23429\,
            PADIN => \N__23428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12412\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23421\,
            DIN => \N__23420\,
            DOUT => \N__23419\,
            PACKAGEPIN => \TVP_VSYNC_wire\
        );

    \TVP_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23421\,
            PADOUT => \N__23420\,
            PADIN => \N__23419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_BLANK_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23412\,
            DIN => \N__23411\,
            DOUT => \N__23410\,
            PACKAGEPIN => \ADV_BLANK_N_wire\
        );

    \ADV_BLANK_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23412\,
            PADOUT => \N__23411\,
            PADIN => \N__23410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22506\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23403\,
            DIN => \N__23402\,
            DOUT => \N__23401\,
            PACKAGEPIN => DEBUG(0)
        );

    \DEBUG_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23403\,
            PADOUT => \N__23402\,
            PADIN => \N__23401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23394\,
            DIN => \N__23393\,
            DOUT => \N__23392\,
            PACKAGEPIN => \ADV_B_wire\(2)
        );

    \ADV_B_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23394\,
            PADOUT => \N__23393\,
            PADIN => \N__23392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12637\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23385\,
            DIN => \N__23384\,
            DOUT => \N__23383\,
            PACKAGEPIN => \ADV_B_wire\(7)
        );

    \ADV_B_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23385\,
            PADOUT => \N__23384\,
            PADIN => \N__23383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12353\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23376\,
            DIN => \N__23375\,
            DOUT => \N__23374\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23376\,
            PADOUT => \N__23375\,
            PADIN => \N__23374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16748\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23367\,
            DIN => \N__23366\,
            DOUT => \N__23365\,
            PACKAGEPIN => \TVP_VIDEO_wire\(4)
        );

    \TVP_VIDEO_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23367\,
            PADOUT => \N__23366\,
            PADIN => \N__23365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23358\,
            DIN => \N__23357\,
            DOUT => \N__23356\,
            PACKAGEPIN => \ADV_G_wire\(3)
        );

    \ADV_G_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23358\,
            PADOUT => \N__23357\,
            PADIN => \N__23356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12580\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23349\,
            DIN => \N__23348\,
            DOUT => \N__23347\,
            PACKAGEPIN => \ADV_HSYNC_wire\
        );

    \ADV_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23349\,
            PADOUT => \N__23348\,
            PADIN => \N__23347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16235\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23340\,
            DIN => \N__23339\,
            DOUT => \N__23338\,
            PACKAGEPIN => \ADV_R_wire\(2)
        );

    \ADV_R_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23340\,
            PADOUT => \N__23339\,
            PADIN => \N__23338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12636\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23331\,
            DIN => \N__23330\,
            DOUT => \N__23329\,
            PACKAGEPIN => \ADV_B_wire\(4)
        );

    \ADV_B_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23331\,
            PADOUT => \N__23330\,
            PADIN => \N__23329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12524\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23322\,
            DIN => \N__23321\,
            DOUT => \N__23320\,
            PACKAGEPIN => DEBUG(4)
        );

    \DEBUG_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23322\,
            PADOUT => \N__23321\,
            PADIN => \N__23320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17528\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23313\,
            DIN => \N__23312\,
            DOUT => \N__23311\,
            PACKAGEPIN => \ADV_G_wire\(6)
        );

    \ADV_G_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23313\,
            PADOUT => \N__23312\,
            PADIN => \N__23311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12411\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23304\,
            DIN => \N__23303\,
            DOUT => \N__23302\,
            PACKAGEPIN => \ADV_R_wire\(7)
        );

    \ADV_R_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23304\,
            PADOUT => \N__23303\,
            PADIN => \N__23302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12349\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23295\,
            DIN => \N__23294\,
            DOUT => \N__23293\,
            PACKAGEPIN => \ADV_B_wire\(3)
        );

    \ADV_B_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23295\,
            PADOUT => \N__23294\,
            PADIN => \N__23293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12581\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23286\,
            DIN => \N__23285\,
            DOUT => \N__23284\,
            PACKAGEPIN => \ADV_R_wire\(4)
        );

    \ADV_R_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23286\,
            PADOUT => \N__23285\,
            PADIN => \N__23284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12523\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23277\,
            DIN => \N__23276\,
            DOUT => \N__23275\,
            PACKAGEPIN => \TVP_VIDEO_wire\(8)
        );

    \TVP_VIDEO_pad_8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23277\,
            PADOUT => \N__23276\,
            PADIN => \N__23275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23268\,
            DIN => \N__23267\,
            DOUT => \N__23266\,
            PACKAGEPIN => \ADV_B_wire\(0)
        );

    \ADV_B_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23268\,
            PADOUT => \N__23267\,
            PADIN => \N__23266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11496\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23259\,
            DIN => \N__23258\,
            DOUT => \N__23257\,
            PACKAGEPIN => \TVP_VIDEO_wire\(5)
        );

    \TVP_VIDEO_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23259\,
            PADOUT => \N__23258\,
            PADIN => \N__23257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23250\,
            DIN => \N__23249\,
            DOUT => \N__23248\,
            PACKAGEPIN => \ADV_G_wire\(2)
        );

    \ADV_G_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23250\,
            PADOUT => \N__23249\,
            PADIN => \N__23248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12638\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23241\,
            DIN => \N__23240\,
            DOUT => \N__23239\,
            PACKAGEPIN => \ADV_VSYNC_wire\
        );

    \ADV_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23241\,
            PADOUT => \N__23240\,
            PADIN => \N__23239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20699\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5604\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23219\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__5601\ : Span4Mux_v
    port map (
            O => \N__23213\,
            I => \N__23210\
        );

    \I__5600\ : Sp12to4
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__5599\ : Span12Mux_h
    port map (
            O => \N__23207\,
            I => \N__23204\
        );

    \I__5598\ : Odrv12
    port map (
            O => \N__23204\,
            I => \line_buffer.n624\
        );

    \I__5597\ : CascadeMux
    port map (
            O => \N__23201\,
            I => \N__23198\
        );

    \I__5596\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__23195\,
            I => \N__23192\
        );

    \I__5594\ : Span4Mux_v
    port map (
            O => \N__23192\,
            I => \N__23189\
        );

    \I__5593\ : Sp12to4
    port map (
            O => \N__23189\,
            I => \N__23186\
        );

    \I__5592\ : Odrv12
    port map (
            O => \N__23186\,
            I => \line_buffer.n632\
        );

    \I__5591\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23180\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__23180\,
            I => \N__23177\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__23177\,
            I => \line_buffer.n3821\
        );

    \I__5588\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23171\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__23171\,
            I => \N__23168\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__23168\,
            I => \N__23165\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__23165\,
            I => \N__23162\
        );

    \I__5584\ : Odrv4
    port map (
            O => \N__23162\,
            I => \line_buffer.n593\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__23159\,
            I => \N__23156\
        );

    \I__5582\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__23153\,
            I => \N__23150\
        );

    \I__5580\ : Span12Mux_v
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__5579\ : Odrv12
    port map (
            O => \N__23147\,
            I => \line_buffer.n601\
        );

    \I__5578\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23138\
        );

    \I__5577\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23126\
        );

    \I__5576\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23122\
        );

    \I__5575\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23119\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__23138\,
            I => \N__23114\
        );

    \I__5573\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23109\
        );

    \I__5572\ : InMux
    port map (
            O => \N__23136\,
            I => \N__23109\
        );

    \I__5571\ : InMux
    port map (
            O => \N__23135\,
            I => \N__23101\
        );

    \I__5570\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23101\
        );

    \I__5569\ : InMux
    port map (
            O => \N__23133\,
            I => \N__23098\
        );

    \I__5568\ : InMux
    port map (
            O => \N__23132\,
            I => \N__23095\
        );

    \I__5567\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23087\
        );

    \I__5566\ : InMux
    port map (
            O => \N__23130\,
            I => \N__23084\
        );

    \I__5565\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23081\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__23126\,
            I => \N__23078\
        );

    \I__5563\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23075\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__23122\,
            I => \N__23072\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__23119\,
            I => \N__23069\
        );

    \I__5560\ : InMux
    port map (
            O => \N__23118\,
            I => \N__23066\
        );

    \I__5559\ : InMux
    port map (
            O => \N__23117\,
            I => \N__23063\
        );

    \I__5558\ : Span4Mux_v
    port map (
            O => \N__23114\,
            I => \N__23060\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__23109\,
            I => \N__23057\
        );

    \I__5556\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23054\
        );

    \I__5555\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23051\
        );

    \I__5554\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23048\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__23045\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__23098\,
            I => \N__23042\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__23095\,
            I => \N__23039\
        );

    \I__5550\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23036\
        );

    \I__5549\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23033\
        );

    \I__5548\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23030\
        );

    \I__5547\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23025\
        );

    \I__5546\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23025\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__23087\,
            I => \N__23016\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__23016\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__23081\,
            I => \N__23016\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__23078\,
            I => \N__23016\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__23075\,
            I => \N__23013\
        );

    \I__5540\ : Span4Mux_v
    port map (
            O => \N__23072\,
            I => \N__23008\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__23069\,
            I => \N__23008\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23005\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__23063\,
            I => \N__23002\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__23060\,
            I => \N__22997\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__23057\,
            I => \N__22997\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__23054\,
            I => \N__22994\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__23051\,
            I => \N__22991\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__23048\,
            I => \N__22986\
        );

    \I__5531\ : Span4Mux_v
    port map (
            O => \N__23045\,
            I => \N__22986\
        );

    \I__5530\ : Span4Mux_h
    port map (
            O => \N__23042\,
            I => \N__22981\
        );

    \I__5529\ : Span4Mux_v
    port map (
            O => \N__23039\,
            I => \N__22981\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__23036\,
            I => \N__22970\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__23033\,
            I => \N__22970\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__23030\,
            I => \N__22970\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__22970\
        );

    \I__5524\ : Span4Mux_v
    port map (
            O => \N__23016\,
            I => \N__22970\
        );

    \I__5523\ : Span4Mux_v
    port map (
            O => \N__23013\,
            I => \N__22965\
        );

    \I__5522\ : Span4Mux_h
    port map (
            O => \N__23008\,
            I => \N__22965\
        );

    \I__5521\ : Span4Mux_v
    port map (
            O => \N__23005\,
            I => \N__22960\
        );

    \I__5520\ : Span4Mux_v
    port map (
            O => \N__23002\,
            I => \N__22960\
        );

    \I__5519\ : Span4Mux_h
    port map (
            O => \N__22997\,
            I => \N__22955\
        );

    \I__5518\ : Span4Mux_v
    port map (
            O => \N__22994\,
            I => \N__22955\
        );

    \I__5517\ : Span4Mux_v
    port map (
            O => \N__22991\,
            I => \N__22946\
        );

    \I__5516\ : Span4Mux_h
    port map (
            O => \N__22986\,
            I => \N__22946\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__22981\,
            I => \N__22946\
        );

    \I__5514\ : Span4Mux_v
    port map (
            O => \N__22970\,
            I => \N__22946\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__22965\,
            I => \N__22943\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__22960\,
            I => \TX_ADDR_11\
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__22955\,
            I => \TX_ADDR_11\
        );

    \I__5510\ : Odrv4
    port map (
            O => \N__22946\,
            I => \TX_ADDR_11\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__22943\,
            I => \TX_ADDR_11\
        );

    \I__5508\ : InMux
    port map (
            O => \N__22934\,
            I => \N__22922\
        );

    \I__5507\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22915\
        );

    \I__5506\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22912\
        );

    \I__5505\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22909\
        );

    \I__5504\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22904\
        );

    \I__5503\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22901\
        );

    \I__5502\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22898\
        );

    \I__5501\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22893\
        );

    \I__5500\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22888\
        );

    \I__5499\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22885\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__22922\,
            I => \N__22882\
        );

    \I__5497\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22873\
        );

    \I__5496\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22873\
        );

    \I__5495\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22873\
        );

    \I__5494\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22873\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__22915\,
            I => \N__22867\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__22912\,
            I => \N__22867\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__22909\,
            I => \N__22861\
        );

    \I__5490\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22858\
        );

    \I__5489\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22855\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__22904\,
            I => \N__22850\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__22901\,
            I => \N__22850\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__22898\,
            I => \N__22847\
        );

    \I__5485\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22842\
        );

    \I__5484\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22842\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__22893\,
            I => \N__22839\
        );

    \I__5482\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22836\
        );

    \I__5481\ : InMux
    port map (
            O => \N__22891\,
            I => \N__22833\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__22888\,
            I => \N__22827\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__22885\,
            I => \N__22827\
        );

    \I__5478\ : Span4Mux_h
    port map (
            O => \N__22882\,
            I => \N__22824\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__22873\,
            I => \N__22821\
        );

    \I__5476\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22818\
        );

    \I__5475\ : Span4Mux_v
    port map (
            O => \N__22867\,
            I => \N__22815\
        );

    \I__5474\ : InMux
    port map (
            O => \N__22866\,
            I => \N__22812\
        );

    \I__5473\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22807\
        );

    \I__5472\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22807\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__22861\,
            I => \N__22802\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__22858\,
            I => \N__22802\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__22855\,
            I => \N__22795\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__22850\,
            I => \N__22795\
        );

    \I__5467\ : Span4Mux_h
    port map (
            O => \N__22847\,
            I => \N__22795\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__22842\,
            I => \N__22788\
        );

    \I__5465\ : Span4Mux_v
    port map (
            O => \N__22839\,
            I => \N__22788\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__22836\,
            I => \N__22788\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__22833\,
            I => \N__22785\
        );

    \I__5462\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22782\
        );

    \I__5461\ : Span4Mux_v
    port map (
            O => \N__22827\,
            I => \N__22779\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__22824\,
            I => \N__22774\
        );

    \I__5459\ : Span4Mux_h
    port map (
            O => \N__22821\,
            I => \N__22774\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__22818\,
            I => \N__22765\
        );

    \I__5457\ : Sp12to4
    port map (
            O => \N__22815\,
            I => \N__22765\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__22812\,
            I => \N__22765\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__22807\,
            I => \N__22765\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__22802\,
            I => \N__22758\
        );

    \I__5453\ : Span4Mux_v
    port map (
            O => \N__22795\,
            I => \N__22758\
        );

    \I__5452\ : Span4Mux_h
    port map (
            O => \N__22788\,
            I => \N__22758\
        );

    \I__5451\ : Span12Mux_h
    port map (
            O => \N__22785\,
            I => \N__22753\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__22782\,
            I => \N__22753\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__22779\,
            I => \TX_ADDR_12\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__22774\,
            I => \TX_ADDR_12\
        );

    \I__5447\ : Odrv12
    port map (
            O => \N__22765\,
            I => \TX_ADDR_12\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__22758\,
            I => \TX_ADDR_12\
        );

    \I__5445\ : Odrv12
    port map (
            O => \N__22753\,
            I => \TX_ADDR_12\
        );

    \I__5444\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__5441\ : Span4Mux_h
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__5440\ : Span4Mux_v
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__22727\,
            I => \line_buffer.n496\
        );

    \I__5438\ : CascadeMux
    port map (
            O => \N__22724\,
            I => \line_buffer.n3809_cascade_\
        );

    \I__5437\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__5435\ : Span4Mux_v
    port map (
            O => \N__22715\,
            I => \N__22712\
        );

    \I__5434\ : Span4Mux_v
    port map (
            O => \N__22712\,
            I => \N__22709\
        );

    \I__5433\ : Span4Mux_h
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__5432\ : Odrv4
    port map (
            O => \N__22706\,
            I => \line_buffer.n504\
        );

    \I__5431\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22700\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__5429\ : Odrv12
    port map (
            O => \N__22697\,
            I => \line_buffer.n3812\
        );

    \I__5428\ : SRMux
    port map (
            O => \N__22694\,
            I => \N__22690\
        );

    \I__5427\ : SRMux
    port map (
            O => \N__22693\,
            I => \N__22687\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__22690\,
            I => \N__22679\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__22687\,
            I => \N__22679\
        );

    \I__5424\ : SRMux
    port map (
            O => \N__22686\,
            I => \N__22676\
        );

    \I__5423\ : SRMux
    port map (
            O => \N__22685\,
            I => \N__22673\
        );

    \I__5422\ : SRMux
    port map (
            O => \N__22684\,
            I => \N__22668\
        );

    \I__5421\ : Span4Mux_s2_v
    port map (
            O => \N__22679\,
            I => \N__22660\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__22676\,
            I => \N__22660\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__22673\,
            I => \N__22660\
        );

    \I__5418\ : SRMux
    port map (
            O => \N__22672\,
            I => \N__22657\
        );

    \I__5417\ : SRMux
    port map (
            O => \N__22671\,
            I => \N__22654\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__22668\,
            I => \N__22649\
        );

    \I__5415\ : SRMux
    port map (
            O => \N__22667\,
            I => \N__22646\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__22660\,
            I => \N__22638\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__22657\,
            I => \N__22638\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22638\
        );

    \I__5411\ : SRMux
    port map (
            O => \N__22653\,
            I => \N__22635\
        );

    \I__5410\ : SRMux
    port map (
            O => \N__22652\,
            I => \N__22632\
        );

    \I__5409\ : Span4Mux_h
    port map (
            O => \N__22649\,
            I => \N__22628\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22625\
        );

    \I__5407\ : SRMux
    port map (
            O => \N__22645\,
            I => \N__22622\
        );

    \I__5406\ : Span4Mux_v
    port map (
            O => \N__22638\,
            I => \N__22615\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__22635\,
            I => \N__22615\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__22632\,
            I => \N__22612\
        );

    \I__5403\ : SRMux
    port map (
            O => \N__22631\,
            I => \N__22609\
        );

    \I__5402\ : Span4Mux_v
    port map (
            O => \N__22628\,
            I => \N__22602\
        );

    \I__5401\ : Span4Mux_h
    port map (
            O => \N__22625\,
            I => \N__22602\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__22622\,
            I => \N__22599\
        );

    \I__5399\ : SRMux
    port map (
            O => \N__22621\,
            I => \N__22596\
        );

    \I__5398\ : SRMux
    port map (
            O => \N__22620\,
            I => \N__22593\
        );

    \I__5397\ : Span4Mux_v
    port map (
            O => \N__22615\,
            I => \N__22585\
        );

    \I__5396\ : Span4Mux_h
    port map (
            O => \N__22612\,
            I => \N__22585\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__22609\,
            I => \N__22582\
        );

    \I__5394\ : SRMux
    port map (
            O => \N__22608\,
            I => \N__22579\
        );

    \I__5393\ : SRMux
    port map (
            O => \N__22607\,
            I => \N__22576\
        );

    \I__5392\ : Span4Mux_v
    port map (
            O => \N__22602\,
            I => \N__22567\
        );

    \I__5391\ : Span4Mux_h
    port map (
            O => \N__22599\,
            I => \N__22567\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__22596\,
            I => \N__22567\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__22593\,
            I => \N__22564\
        );

    \I__5388\ : SRMux
    port map (
            O => \N__22592\,
            I => \N__22561\
        );

    \I__5387\ : SRMux
    port map (
            O => \N__22591\,
            I => \N__22558\
        );

    \I__5386\ : SRMux
    port map (
            O => \N__22590\,
            I => \N__22551\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__22585\,
            I => \N__22546\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__22582\,
            I => \N__22546\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__22579\,
            I => \N__22541\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__22576\,
            I => \N__22541\
        );

    \I__5381\ : SRMux
    port map (
            O => \N__22575\,
            I => \N__22538\
        );

    \I__5380\ : SRMux
    port map (
            O => \N__22574\,
            I => \N__22535\
        );

    \I__5379\ : Span4Mux_v
    port map (
            O => \N__22567\,
            I => \N__22526\
        );

    \I__5378\ : Span4Mux_h
    port map (
            O => \N__22564\,
            I => \N__22526\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__22561\,
            I => \N__22526\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__22558\,
            I => \N__22523\
        );

    \I__5375\ : SRMux
    port map (
            O => \N__22557\,
            I => \N__22520\
        );

    \I__5374\ : SRMux
    port map (
            O => \N__22556\,
            I => \N__22517\
        );

    \I__5373\ : SRMux
    port map (
            O => \N__22555\,
            I => \N__22512\
        );

    \I__5372\ : SRMux
    port map (
            O => \N__22554\,
            I => \N__22509\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__22551\,
            I => \N__22503\
        );

    \I__5370\ : Span4Mux_v
    port map (
            O => \N__22546\,
            I => \N__22494\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__22541\,
            I => \N__22494\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22494\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__22535\,
            I => \N__22494\
        );

    \I__5366\ : SRMux
    port map (
            O => \N__22534\,
            I => \N__22491\
        );

    \I__5365\ : SRMux
    port map (
            O => \N__22533\,
            I => \N__22488\
        );

    \I__5364\ : Span4Mux_v
    port map (
            O => \N__22526\,
            I => \N__22481\
        );

    \I__5363\ : Span4Mux_h
    port map (
            O => \N__22523\,
            I => \N__22481\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22481\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__22517\,
            I => \N__22478\
        );

    \I__5360\ : SRMux
    port map (
            O => \N__22516\,
            I => \N__22475\
        );

    \I__5359\ : SRMux
    port map (
            O => \N__22515\,
            I => \N__22472\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__22512\,
            I => \N__22466\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__22509\,
            I => \N__22466\
        );

    \I__5356\ : SRMux
    port map (
            O => \N__22508\,
            I => \N__22463\
        );

    \I__5355\ : IoInMux
    port map (
            O => \N__22507\,
            I => \N__22460\
        );

    \I__5354\ : IoInMux
    port map (
            O => \N__22506\,
            I => \N__22457\
        );

    \I__5353\ : Sp12to4
    port map (
            O => \N__22503\,
            I => \N__22454\
        );

    \I__5352\ : Span4Mux_v
    port map (
            O => \N__22494\,
            I => \N__22449\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22449\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__22488\,
            I => \N__22446\
        );

    \I__5349\ : Span4Mux_v
    port map (
            O => \N__22481\,
            I => \N__22439\
        );

    \I__5348\ : Span4Mux_h
    port map (
            O => \N__22478\,
            I => \N__22439\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__22475\,
            I => \N__22439\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22436\
        );

    \I__5345\ : SRMux
    port map (
            O => \N__22471\,
            I => \N__22433\
        );

    \I__5344\ : Span12Mux_s6_v
    port map (
            O => \N__22466\,
            I => \N__22427\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__22463\,
            I => \N__22427\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__22460\,
            I => \N__22422\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__22457\,
            I => \N__22422\
        );

    \I__5340\ : Span12Mux_v
    port map (
            O => \N__22454\,
            I => \N__22419\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__22449\,
            I => \N__22414\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__22446\,
            I => \N__22414\
        );

    \I__5337\ : Span4Mux_v
    port map (
            O => \N__22439\,
            I => \N__22407\
        );

    \I__5336\ : Span4Mux_h
    port map (
            O => \N__22436\,
            I => \N__22407\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__22433\,
            I => \N__22407\
        );

    \I__5334\ : SRMux
    port map (
            O => \N__22432\,
            I => \N__22404\
        );

    \I__5333\ : Span12Mux_v
    port map (
            O => \N__22427\,
            I => \N__22401\
        );

    \I__5332\ : Span4Mux_s2_v
    port map (
            O => \N__22422\,
            I => \N__22398\
        );

    \I__5331\ : Span12Mux_h
    port map (
            O => \N__22419\,
            I => \N__22395\
        );

    \I__5330\ : Sp12to4
    port map (
            O => \N__22414\,
            I => \N__22392\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__22407\,
            I => \N__22387\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__22404\,
            I => \N__22387\
        );

    \I__5327\ : Span12Mux_v
    port map (
            O => \N__22401\,
            I => \N__22384\
        );

    \I__5326\ : Span4Mux_h
    port map (
            O => \N__22398\,
            I => \N__22381\
        );

    \I__5325\ : Span12Mux_v
    port map (
            O => \N__22395\,
            I => \N__22374\
        );

    \I__5324\ : Span12Mux_h
    port map (
            O => \N__22392\,
            I => \N__22374\
        );

    \I__5323\ : Sp12to4
    port map (
            O => \N__22387\,
            I => \N__22374\
        );

    \I__5322\ : Odrv12
    port map (
            O => \N__22384\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__22381\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5320\ : Odrv12
    port map (
            O => \N__22374\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5319\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__5317\ : Odrv12
    port map (
            O => \N__22361\,
            I => \line_buffer.n507\
        );

    \I__5316\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__5314\ : Span4Mux_v
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__5313\ : Sp12to4
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__5312\ : Span12Mux_h
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__5311\ : Odrv12
    port map (
            O => \N__22343\,
            I => \line_buffer.n499\
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__5309\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__22331\,
            I => \line_buffer.n3720\
        );

    \I__5306\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__5304\ : Span4Mux_v
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__22316\,
            I => \line_buffer.n592\
        );

    \I__5301\ : CascadeMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__5300\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__5298\ : Span4Mux_v
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__22295\,
            I => \line_buffer.n600\
        );

    \I__5294\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__22289\,
            I => \N__22286\
        );

    \I__5292\ : Sp12to4
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__5291\ : Span12Mux_v
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__5290\ : Odrv12
    port map (
            O => \N__22280\,
            I => \line_buffer.n572\
        );

    \I__5289\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__5287\ : Span4Mux_v
    port map (
            O => \N__22271\,
            I => \N__22268\
        );

    \I__5286\ : Span4Mux_h
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__22265\,
            I => \line_buffer.n564\
        );

    \I__5284\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__5282\ : Span4Mux_h
    port map (
            O => \N__22256\,
            I => \N__22253\
        );

    \I__5281\ : Span4Mux_v
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__5280\ : Span4Mux_v
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__5279\ : Span4Mux_h
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__22244\,
            I => \line_buffer.n503\
        );

    \I__5277\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22238\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__22238\,
            I => \line_buffer.n3815\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__22235\,
            I => \N__22232\
        );

    \I__5274\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22229\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__22229\,
            I => \N__22226\
        );

    \I__5272\ : Span4Mux_v
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__5271\ : Span4Mux_h
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__5270\ : Span4Mux_v
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__5269\ : Span4Mux_v
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__22214\,
            I => \line_buffer.n495\
        );

    \I__5267\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__5265\ : Sp12to4
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__5264\ : Span12Mux_v
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__5263\ : Odrv12
    port map (
            O => \N__22199\,
            I => \line_buffer.n568\
        );

    \I__5262\ : CascadeMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__5261\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__22181\,
            I => \line_buffer.n560\
        );

    \I__5256\ : CascadeMux
    port map (
            O => \N__22178\,
            I => \line_buffer.n3824_cascade_\
        );

    \I__5255\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__22172\,
            I => \line_buffer.n3818\
        );

    \I__5253\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__5251\ : Odrv12
    port map (
            O => \N__22163\,
            I => \TX_DATA_0\
        );

    \I__5250\ : ClkMux
    port map (
            O => \N__22160\,
            I => \N__22155\
        );

    \I__5249\ : ClkMux
    port map (
            O => \N__22159\,
            I => \N__22152\
        );

    \I__5248\ : ClkMux
    port map (
            O => \N__22158\,
            I => \N__22146\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__22155\,
            I => \N__22134\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__22152\,
            I => \N__22131\
        );

    \I__5245\ : ClkMux
    port map (
            O => \N__22151\,
            I => \N__22128\
        );

    \I__5244\ : ClkMux
    port map (
            O => \N__22150\,
            I => \N__22125\
        );

    \I__5243\ : ClkMux
    port map (
            O => \N__22149\,
            I => \N__22120\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__22146\,
            I => \N__22114\
        );

    \I__5241\ : ClkMux
    port map (
            O => \N__22145\,
            I => \N__22111\
        );

    \I__5240\ : ClkMux
    port map (
            O => \N__22144\,
            I => \N__22108\
        );

    \I__5239\ : ClkMux
    port map (
            O => \N__22143\,
            I => \N__22105\
        );

    \I__5238\ : ClkMux
    port map (
            O => \N__22142\,
            I => \N__22100\
        );

    \I__5237\ : ClkMux
    port map (
            O => \N__22141\,
            I => \N__22096\
        );

    \I__5236\ : ClkMux
    port map (
            O => \N__22140\,
            I => \N__22092\
        );

    \I__5235\ : ClkMux
    port map (
            O => \N__22139\,
            I => \N__22081\
        );

    \I__5234\ : ClkMux
    port map (
            O => \N__22138\,
            I => \N__22078\
        );

    \I__5233\ : ClkMux
    port map (
            O => \N__22137\,
            I => \N__22074\
        );

    \I__5232\ : Span4Mux_s2_v
    port map (
            O => \N__22134\,
            I => \N__22063\
        );

    \I__5231\ : Span4Mux_h
    port map (
            O => \N__22131\,
            I => \N__22063\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22063\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__22125\,
            I => \N__22060\
        );

    \I__5228\ : ClkMux
    port map (
            O => \N__22124\,
            I => \N__22057\
        );

    \I__5227\ : ClkMux
    port map (
            O => \N__22123\,
            I => \N__22054\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__22120\,
            I => \N__22049\
        );

    \I__5225\ : ClkMux
    port map (
            O => \N__22119\,
            I => \N__22046\
        );

    \I__5224\ : ClkMux
    port map (
            O => \N__22118\,
            I => \N__22043\
        );

    \I__5223\ : ClkMux
    port map (
            O => \N__22117\,
            I => \N__22038\
        );

    \I__5222\ : Span4Mux_h
    port map (
            O => \N__22114\,
            I => \N__22032\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__22111\,
            I => \N__22032\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__22108\,
            I => \N__22027\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__22105\,
            I => \N__22027\
        );

    \I__5218\ : ClkMux
    port map (
            O => \N__22104\,
            I => \N__22024\
        );

    \I__5217\ : ClkMux
    port map (
            O => \N__22103\,
            I => \N__22021\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__22100\,
            I => \N__22018\
        );

    \I__5215\ : ClkMux
    port map (
            O => \N__22099\,
            I => \N__22015\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__22096\,
            I => \N__22011\
        );

    \I__5213\ : ClkMux
    port map (
            O => \N__22095\,
            I => \N__22008\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__22092\,
            I => \N__22004\
        );

    \I__5211\ : ClkMux
    port map (
            O => \N__22091\,
            I => \N__22001\
        );

    \I__5210\ : ClkMux
    port map (
            O => \N__22090\,
            I => \N__21998\
        );

    \I__5209\ : ClkMux
    port map (
            O => \N__22089\,
            I => \N__21994\
        );

    \I__5208\ : ClkMux
    port map (
            O => \N__22088\,
            I => \N__21991\
        );

    \I__5207\ : ClkMux
    port map (
            O => \N__22087\,
            I => \N__21988\
        );

    \I__5206\ : ClkMux
    port map (
            O => \N__22086\,
            I => \N__21984\
        );

    \I__5205\ : ClkMux
    port map (
            O => \N__22085\,
            I => \N__21980\
        );

    \I__5204\ : ClkMux
    port map (
            O => \N__22084\,
            I => \N__21977\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__22081\,
            I => \N__21973\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__21970\
        );

    \I__5201\ : ClkMux
    port map (
            O => \N__22077\,
            I => \N__21967\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__22074\,
            I => \N__21963\
        );

    \I__5199\ : ClkMux
    port map (
            O => \N__22073\,
            I => \N__21960\
        );

    \I__5198\ : ClkMux
    port map (
            O => \N__22072\,
            I => \N__21953\
        );

    \I__5197\ : ClkMux
    port map (
            O => \N__22071\,
            I => \N__21950\
        );

    \I__5196\ : ClkMux
    port map (
            O => \N__22070\,
            I => \N__21943\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__22063\,
            I => \N__21936\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__22060\,
            I => \N__21936\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__21936\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__22054\,
            I => \N__21933\
        );

    \I__5191\ : ClkMux
    port map (
            O => \N__22053\,
            I => \N__21930\
        );

    \I__5190\ : ClkMux
    port map (
            O => \N__22052\,
            I => \N__21927\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__22049\,
            I => \N__21921\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__22046\,
            I => \N__21918\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__22043\,
            I => \N__21915\
        );

    \I__5186\ : ClkMux
    port map (
            O => \N__22042\,
            I => \N__21912\
        );

    \I__5185\ : ClkMux
    port map (
            O => \N__22041\,
            I => \N__21909\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__21905\
        );

    \I__5183\ : ClkMux
    port map (
            O => \N__22037\,
            I => \N__21902\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__22032\,
            I => \N__21893\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__22027\,
            I => \N__21893\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__22024\,
            I => \N__21893\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__21893\
        );

    \I__5178\ : Span4Mux_v
    port map (
            O => \N__22018\,
            I => \N__21888\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__22015\,
            I => \N__21888\
        );

    \I__5176\ : ClkMux
    port map (
            O => \N__22014\,
            I => \N__21885\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__22011\,
            I => \N__21880\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__22008\,
            I => \N__21880\
        );

    \I__5173\ : ClkMux
    port map (
            O => \N__22007\,
            I => \N__21877\
        );

    \I__5172\ : Span4Mux_v
    port map (
            O => \N__22004\,
            I => \N__21870\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__22001\,
            I => \N__21870\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__21998\,
            I => \N__21867\
        );

    \I__5169\ : ClkMux
    port map (
            O => \N__21997\,
            I => \N__21864\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__21994\,
            I => \N__21859\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__21991\,
            I => \N__21859\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__21988\,
            I => \N__21856\
        );

    \I__5165\ : ClkMux
    port map (
            O => \N__21987\,
            I => \N__21853\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__21984\,
            I => \N__21850\
        );

    \I__5163\ : ClkMux
    port map (
            O => \N__21983\,
            I => \N__21847\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21842\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__21977\,
            I => \N__21842\
        );

    \I__5160\ : ClkMux
    port map (
            O => \N__21976\,
            I => \N__21839\
        );

    \I__5159\ : Span4Mux_h
    port map (
            O => \N__21973\,
            I => \N__21832\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__21970\,
            I => \N__21832\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__21967\,
            I => \N__21832\
        );

    \I__5156\ : ClkMux
    port map (
            O => \N__21966\,
            I => \N__21829\
        );

    \I__5155\ : Span4Mux_h
    port map (
            O => \N__21963\,
            I => \N__21824\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__21960\,
            I => \N__21821\
        );

    \I__5153\ : ClkMux
    port map (
            O => \N__21959\,
            I => \N__21818\
        );

    \I__5152\ : ClkMux
    port map (
            O => \N__21958\,
            I => \N__21813\
        );

    \I__5151\ : ClkMux
    port map (
            O => \N__21957\,
            I => \N__21810\
        );

    \I__5150\ : IoInMux
    port map (
            O => \N__21956\,
            I => \N__21805\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__21953\,
            I => \N__21799\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__21950\,
            I => \N__21799\
        );

    \I__5147\ : ClkMux
    port map (
            O => \N__21949\,
            I => \N__21796\
        );

    \I__5146\ : ClkMux
    port map (
            O => \N__21948\,
            I => \N__21793\
        );

    \I__5145\ : ClkMux
    port map (
            O => \N__21947\,
            I => \N__21790\
        );

    \I__5144\ : ClkMux
    port map (
            O => \N__21946\,
            I => \N__21787\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__21943\,
            I => \N__21783\
        );

    \I__5142\ : Span4Mux_v
    port map (
            O => \N__21936\,
            I => \N__21775\
        );

    \I__5141\ : Span4Mux_h
    port map (
            O => \N__21933\,
            I => \N__21775\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__21930\,
            I => \N__21775\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__21927\,
            I => \N__21772\
        );

    \I__5138\ : ClkMux
    port map (
            O => \N__21926\,
            I => \N__21769\
        );

    \I__5137\ : ClkMux
    port map (
            O => \N__21925\,
            I => \N__21766\
        );

    \I__5136\ : ClkMux
    port map (
            O => \N__21924\,
            I => \N__21762\
        );

    \I__5135\ : Span4Mux_h
    port map (
            O => \N__21921\,
            I => \N__21753\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__21918\,
            I => \N__21753\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__21915\,
            I => \N__21753\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__21912\,
            I => \N__21753\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__21909\,
            I => \N__21750\
        );

    \I__5130\ : ClkMux
    port map (
            O => \N__21908\,
            I => \N__21747\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__21905\,
            I => \N__21742\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__21902\,
            I => \N__21742\
        );

    \I__5127\ : Span4Mux_v
    port map (
            O => \N__21893\,
            I => \N__21735\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__21888\,
            I => \N__21735\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__21885\,
            I => \N__21735\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__21880\,
            I => \N__21730\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__21877\,
            I => \N__21730\
        );

    \I__5122\ : ClkMux
    port map (
            O => \N__21876\,
            I => \N__21727\
        );

    \I__5121\ : ClkMux
    port map (
            O => \N__21875\,
            I => \N__21724\
        );

    \I__5120\ : Span4Mux_v
    port map (
            O => \N__21870\,
            I => \N__21720\
        );

    \I__5119\ : Span4Mux_v
    port map (
            O => \N__21867\,
            I => \N__21715\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__21864\,
            I => \N__21715\
        );

    \I__5117\ : Span4Mux_v
    port map (
            O => \N__21859\,
            I => \N__21708\
        );

    \I__5116\ : Span4Mux_h
    port map (
            O => \N__21856\,
            I => \N__21708\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__21853\,
            I => \N__21708\
        );

    \I__5114\ : Span4Mux_v
    port map (
            O => \N__21850\,
            I => \N__21703\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21703\
        );

    \I__5112\ : Span4Mux_v
    port map (
            O => \N__21842\,
            I => \N__21698\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__21839\,
            I => \N__21698\
        );

    \I__5110\ : Span4Mux_h
    port map (
            O => \N__21832\,
            I => \N__21693\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__21829\,
            I => \N__21693\
        );

    \I__5108\ : ClkMux
    port map (
            O => \N__21828\,
            I => \N__21690\
        );

    \I__5107\ : ClkMux
    port map (
            O => \N__21827\,
            I => \N__21687\
        );

    \I__5106\ : Span4Mux_v
    port map (
            O => \N__21824\,
            I => \N__21677\
        );

    \I__5105\ : Span4Mux_h
    port map (
            O => \N__21821\,
            I => \N__21677\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__21818\,
            I => \N__21674\
        );

    \I__5103\ : ClkMux
    port map (
            O => \N__21817\,
            I => \N__21671\
        );

    \I__5102\ : ClkMux
    port map (
            O => \N__21816\,
            I => \N__21668\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__21813\,
            I => \N__21662\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21810\,
            I => \N__21662\
        );

    \I__5099\ : ClkMux
    port map (
            O => \N__21809\,
            I => \N__21659\
        );

    \I__5098\ : ClkMux
    port map (
            O => \N__21808\,
            I => \N__21656\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__21805\,
            I => \N__21653\
        );

    \I__5096\ : ClkMux
    port map (
            O => \N__21804\,
            I => \N__21650\
        );

    \I__5095\ : Span4Mux_v
    port map (
            O => \N__21799\,
            I => \N__21641\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__21796\,
            I => \N__21641\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__21793\,
            I => \N__21641\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__21790\,
            I => \N__21641\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__21787\,
            I => \N__21638\
        );

    \I__5090\ : ClkMux
    port map (
            O => \N__21786\,
            I => \N__21635\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__21783\,
            I => \N__21632\
        );

    \I__5088\ : ClkMux
    port map (
            O => \N__21782\,
            I => \N__21629\
        );

    \I__5087\ : Span4Mux_v
    port map (
            O => \N__21775\,
            I => \N__21621\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__21772\,
            I => \N__21621\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__21769\,
            I => \N__21621\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__21766\,
            I => \N__21618\
        );

    \I__5083\ : ClkMux
    port map (
            O => \N__21765\,
            I => \N__21615\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__21762\,
            I => \N__21612\
        );

    \I__5081\ : Span4Mux_v
    port map (
            O => \N__21753\,
            I => \N__21609\
        );

    \I__5080\ : Span4Mux_v
    port map (
            O => \N__21750\,
            I => \N__21604\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21747\,
            I => \N__21604\
        );

    \I__5078\ : Span4Mux_v
    port map (
            O => \N__21742\,
            I => \N__21593\
        );

    \I__5077\ : Span4Mux_h
    port map (
            O => \N__21735\,
            I => \N__21593\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__21730\,
            I => \N__21593\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21593\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__21724\,
            I => \N__21593\
        );

    \I__5073\ : ClkMux
    port map (
            O => \N__21723\,
            I => \N__21590\
        );

    \I__5072\ : Span4Mux_v
    port map (
            O => \N__21720\,
            I => \N__21585\
        );

    \I__5071\ : Span4Mux_v
    port map (
            O => \N__21715\,
            I => \N__21585\
        );

    \I__5070\ : Span4Mux_h
    port map (
            O => \N__21708\,
            I => \N__21572\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__21703\,
            I => \N__21572\
        );

    \I__5068\ : Span4Mux_v
    port map (
            O => \N__21698\,
            I => \N__21572\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__21693\,
            I => \N__21572\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__21690\,
            I => \N__21572\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21572\
        );

    \I__5064\ : ClkMux
    port map (
            O => \N__21686\,
            I => \N__21569\
        );

    \I__5063\ : ClkMux
    port map (
            O => \N__21685\,
            I => \N__21566\
        );

    \I__5062\ : ClkMux
    port map (
            O => \N__21684\,
            I => \N__21563\
        );

    \I__5061\ : ClkMux
    port map (
            O => \N__21683\,
            I => \N__21560\
        );

    \I__5060\ : ClkMux
    port map (
            O => \N__21682\,
            I => \N__21554\
        );

    \I__5059\ : Span4Mux_v
    port map (
            O => \N__21677\,
            I => \N__21548\
        );

    \I__5058\ : Span4Mux_h
    port map (
            O => \N__21674\,
            I => \N__21548\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__21671\,
            I => \N__21545\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__21668\,
            I => \N__21542\
        );

    \I__5055\ : ClkMux
    port map (
            O => \N__21667\,
            I => \N__21539\
        );

    \I__5054\ : Span4Mux_v
    port map (
            O => \N__21662\,
            I => \N__21532\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21659\,
            I => \N__21532\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__21656\,
            I => \N__21532\
        );

    \I__5051\ : Span4Mux_s2_v
    port map (
            O => \N__21653\,
            I => \N__21529\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__21650\,
            I => \N__21526\
        );

    \I__5049\ : Span4Mux_v
    port map (
            O => \N__21641\,
            I => \N__21523\
        );

    \I__5048\ : Span4Mux_v
    port map (
            O => \N__21638\,
            I => \N__21518\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__21635\,
            I => \N__21518\
        );

    \I__5046\ : Span4Mux_v
    port map (
            O => \N__21632\,
            I => \N__21513\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__21629\,
            I => \N__21513\
        );

    \I__5044\ : ClkMux
    port map (
            O => \N__21628\,
            I => \N__21510\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__21621\,
            I => \N__21502\
        );

    \I__5042\ : Span4Mux_h
    port map (
            O => \N__21618\,
            I => \N__21502\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__21615\,
            I => \N__21502\
        );

    \I__5040\ : Span4Mux_v
    port map (
            O => \N__21612\,
            I => \N__21499\
        );

    \I__5039\ : Span4Mux_v
    port map (
            O => \N__21609\,
            I => \N__21496\
        );

    \I__5038\ : Span4Mux_v
    port map (
            O => \N__21604\,
            I => \N__21491\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__21593\,
            I => \N__21491\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__21590\,
            I => \N__21487\
        );

    \I__5035\ : Span4Mux_v
    port map (
            O => \N__21585\,
            I => \N__21480\
        );

    \I__5034\ : Span4Mux_h
    port map (
            O => \N__21572\,
            I => \N__21480\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21480\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__21566\,
            I => \N__21476\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__21563\,
            I => \N__21471\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__21560\,
            I => \N__21471\
        );

    \I__5029\ : ClkMux
    port map (
            O => \N__21559\,
            I => \N__21468\
        );

    \I__5028\ : ClkMux
    port map (
            O => \N__21558\,
            I => \N__21465\
        );

    \I__5027\ : ClkMux
    port map (
            O => \N__21557\,
            I => \N__21462\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__21554\,
            I => \N__21459\
        );

    \I__5025\ : ClkMux
    port map (
            O => \N__21553\,
            I => \N__21456\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__21548\,
            I => \N__21447\
        );

    \I__5023\ : Span4Mux_h
    port map (
            O => \N__21545\,
            I => \N__21447\
        );

    \I__5022\ : Span4Mux_h
    port map (
            O => \N__21542\,
            I => \N__21447\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__21539\,
            I => \N__21447\
        );

    \I__5020\ : Span4Mux_v
    port map (
            O => \N__21532\,
            I => \N__21439\
        );

    \I__5019\ : Span4Mux_h
    port map (
            O => \N__21529\,
            I => \N__21439\
        );

    \I__5018\ : Span4Mux_s2_v
    port map (
            O => \N__21526\,
            I => \N__21439\
        );

    \I__5017\ : Span4Mux_v
    port map (
            O => \N__21523\,
            I => \N__21434\
        );

    \I__5016\ : Span4Mux_v
    port map (
            O => \N__21518\,
            I => \N__21434\
        );

    \I__5015\ : Span4Mux_v
    port map (
            O => \N__21513\,
            I => \N__21429\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__21510\,
            I => \N__21429\
        );

    \I__5013\ : ClkMux
    port map (
            O => \N__21509\,
            I => \N__21426\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__21502\,
            I => \N__21423\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__21499\,
            I => \N__21416\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__21496\,
            I => \N__21416\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__21491\,
            I => \N__21416\
        );

    \I__5008\ : ClkMux
    port map (
            O => \N__21490\,
            I => \N__21413\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__21487\,
            I => \N__21408\
        );

    \I__5006\ : Span4Mux_v
    port map (
            O => \N__21480\,
            I => \N__21408\
        );

    \I__5005\ : ClkMux
    port map (
            O => \N__21479\,
            I => \N__21405\
        );

    \I__5004\ : Span4Mux_v
    port map (
            O => \N__21476\,
            I => \N__21394\
        );

    \I__5003\ : Span4Mux_v
    port map (
            O => \N__21471\,
            I => \N__21394\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__21468\,
            I => \N__21394\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__21465\,
            I => \N__21394\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__21462\,
            I => \N__21394\
        );

    \I__4999\ : Span12Mux_h
    port map (
            O => \N__21459\,
            I => \N__21391\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__21456\,
            I => \N__21388\
        );

    \I__4997\ : Span4Mux_h
    port map (
            O => \N__21447\,
            I => \N__21385\
        );

    \I__4996\ : ClkMux
    port map (
            O => \N__21446\,
            I => \N__21382\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__21439\,
            I => \N__21379\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__21434\,
            I => \N__21376\
        );

    \I__4993\ : Span4Mux_v
    port map (
            O => \N__21429\,
            I => \N__21371\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__21426\,
            I => \N__21371\
        );

    \I__4991\ : Sp12to4
    port map (
            O => \N__21423\,
            I => \N__21366\
        );

    \I__4990\ : Sp12to4
    port map (
            O => \N__21416\,
            I => \N__21366\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__21413\,
            I => \N__21361\
        );

    \I__4988\ : Sp12to4
    port map (
            O => \N__21408\,
            I => \N__21361\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__21405\,
            I => \N__21356\
        );

    \I__4986\ : Sp12to4
    port map (
            O => \N__21394\,
            I => \N__21356\
        );

    \I__4985\ : Span12Mux_v
    port map (
            O => \N__21391\,
            I => \N__21349\
        );

    \I__4984\ : Span12Mux_h
    port map (
            O => \N__21388\,
            I => \N__21349\
        );

    \I__4983\ : Sp12to4
    port map (
            O => \N__21385\,
            I => \N__21349\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__21382\,
            I => \N__21346\
        );

    \I__4981\ : IoSpan4Mux
    port map (
            O => \N__21379\,
            I => \N__21343\
        );

    \I__4980\ : Span4Mux_v
    port map (
            O => \N__21376\,
            I => \N__21340\
        );

    \I__4979\ : Span4Mux_h
    port map (
            O => \N__21371\,
            I => \N__21337\
        );

    \I__4978\ : Span12Mux_h
    port map (
            O => \N__21366\,
            I => \N__21330\
        );

    \I__4977\ : Span12Mux_h
    port map (
            O => \N__21361\,
            I => \N__21330\
        );

    \I__4976\ : Span12Mux_v
    port map (
            O => \N__21356\,
            I => \N__21330\
        );

    \I__4975\ : Span12Mux_v
    port map (
            O => \N__21349\,
            I => \N__21325\
        );

    \I__4974\ : Span12Mux_h
    port map (
            O => \N__21346\,
            I => \N__21325\
        );

    \I__4973\ : IoSpan4Mux
    port map (
            O => \N__21343\,
            I => \N__21322\
        );

    \I__4972\ : Span4Mux_h
    port map (
            O => \N__21340\,
            I => \N__21317\
        );

    \I__4971\ : Span4Mux_h
    port map (
            O => \N__21337\,
            I => \N__21317\
        );

    \I__4970\ : Odrv12
    port map (
            O => \N__21330\,
            I => \ADV_CLK_c\
        );

    \I__4969\ : Odrv12
    port map (
            O => \N__21325\,
            I => \ADV_CLK_c\
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__21322\,
            I => \ADV_CLK_c\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__21317\,
            I => \ADV_CLK_c\
        );

    \I__4966\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21305\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21302\
        );

    \I__4964\ : Span12Mux_v
    port map (
            O => \N__21302\,
            I => \N__21299\
        );

    \I__4963\ : Odrv12
    port map (
            O => \N__21299\,
            I => \line_buffer.n3699\
        );

    \I__4962\ : IoInMux
    port map (
            O => \N__21296\,
            I => \N__21292\
        );

    \I__4961\ : CascadeMux
    port map (
            O => \N__21295\,
            I => \N__21285\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__21292\,
            I => \N__21281\
        );

    \I__4959\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21278\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__21290\,
            I => \N__21273\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__21289\,
            I => \N__21268\
        );

    \I__4956\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21265\
        );

    \I__4955\ : InMux
    port map (
            O => \N__21285\,
            I => \N__21262\
        );

    \I__4954\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21258\
        );

    \I__4953\ : Span4Mux_s3_h
    port map (
            O => \N__21281\,
            I => \N__21254\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__21278\,
            I => \N__21250\
        );

    \I__4951\ : InMux
    port map (
            O => \N__21277\,
            I => \N__21247\
        );

    \I__4950\ : InMux
    port map (
            O => \N__21276\,
            I => \N__21242\
        );

    \I__4949\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21242\
        );

    \I__4948\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21235\
        );

    \I__4947\ : InMux
    port map (
            O => \N__21271\,
            I => \N__21235\
        );

    \I__4946\ : InMux
    port map (
            O => \N__21268\,
            I => \N__21235\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__21265\,
            I => \N__21230\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__21262\,
            I => \N__21230\
        );

    \I__4943\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21227\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__21258\,
            I => \N__21224\
        );

    \I__4941\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21221\
        );

    \I__4940\ : Span4Mux_v
    port map (
            O => \N__21254\,
            I => \N__21218\
        );

    \I__4939\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21215\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__21250\,
            I => \N__21211\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__21247\,
            I => \N__21208\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__21242\,
            I => \N__21203\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21203\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__21230\,
            I => \N__21200\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__21227\,
            I => \N__21197\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__21224\,
            I => \N__21192\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21192\
        );

    \I__4930\ : Sp12to4
    port map (
            O => \N__21218\,
            I => \N__21189\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21186\
        );

    \I__4928\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21183\
        );

    \I__4927\ : Span4Mux_h
    port map (
            O => \N__21211\,
            I => \N__21176\
        );

    \I__4926\ : Span4Mux_v
    port map (
            O => \N__21208\,
            I => \N__21176\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__21203\,
            I => \N__21176\
        );

    \I__4924\ : Span4Mux_h
    port map (
            O => \N__21200\,
            I => \N__21173\
        );

    \I__4923\ : Span4Mux_v
    port map (
            O => \N__21197\,
            I => \N__21168\
        );

    \I__4922\ : Span4Mux_v
    port map (
            O => \N__21192\,
            I => \N__21168\
        );

    \I__4921\ : Odrv12
    port map (
            O => \N__21189\,
            I => \DEBUG_c_2\
        );

    \I__4920\ : Odrv4
    port map (
            O => \N__21186\,
            I => \DEBUG_c_2\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__21183\,
            I => \DEBUG_c_2\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__21176\,
            I => \DEBUG_c_2\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__21173\,
            I => \DEBUG_c_2\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__21168\,
            I => \DEBUG_c_2\
        );

    \I__4915\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__21152\,
            I => \N__21149\
        );

    \I__4913\ : Odrv4
    port map (
            O => \N__21149\,
            I => \line_buffer.n3797\
        );

    \I__4912\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__4910\ : Span4Mux_v
    port map (
            O => \N__21140\,
            I => \N__21137\
        );

    \I__4909\ : Span4Mux_v
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__4908\ : Sp12to4
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__4907\ : Odrv12
    port map (
            O => \N__21131\,
            I => \line_buffer.n636\
        );

    \I__4906\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21125\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__4903\ : Span4Mux_v
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__4901\ : Span4Mux_h
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__21110\,
            I => \line_buffer.n628\
        );

    \I__4899\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__4897\ : Odrv4
    port map (
            O => \N__21101\,
            I => \line_buffer.n3700\
        );

    \I__4896\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21093\
        );

    \I__4895\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21088\
        );

    \I__4894\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21088\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__21093\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__21088\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__4891\ : InMux
    port map (
            O => \N__21083\,
            I => \receive_module.rx_counter.n3363\
        );

    \I__4890\ : InMux
    port map (
            O => \N__21080\,
            I => \N__21076\
        );

    \I__4889\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21073\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__21076\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__21073\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__4886\ : InMux
    port map (
            O => \N__21068\,
            I => \bfn_17_10_0_\
        );

    \I__4885\ : InMux
    port map (
            O => \N__21065\,
            I => \receive_module.rx_counter.n3365\
        );

    \I__4884\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21058\
        );

    \I__4883\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21055\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__21058\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__21055\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__4880\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__21047\,
            I => \N__21036\
        );

    \I__4878\ : ClkMux
    port map (
            O => \N__21046\,
            I => \N__20909\
        );

    \I__4877\ : ClkMux
    port map (
            O => \N__21045\,
            I => \N__20909\
        );

    \I__4876\ : ClkMux
    port map (
            O => \N__21044\,
            I => \N__20909\
        );

    \I__4875\ : ClkMux
    port map (
            O => \N__21043\,
            I => \N__20909\
        );

    \I__4874\ : ClkMux
    port map (
            O => \N__21042\,
            I => \N__20909\
        );

    \I__4873\ : ClkMux
    port map (
            O => \N__21041\,
            I => \N__20909\
        );

    \I__4872\ : ClkMux
    port map (
            O => \N__21040\,
            I => \N__20909\
        );

    \I__4871\ : ClkMux
    port map (
            O => \N__21039\,
            I => \N__20909\
        );

    \I__4870\ : Glb2LocalMux
    port map (
            O => \N__21036\,
            I => \N__20909\
        );

    \I__4869\ : ClkMux
    port map (
            O => \N__21035\,
            I => \N__20909\
        );

    \I__4868\ : ClkMux
    port map (
            O => \N__21034\,
            I => \N__20909\
        );

    \I__4867\ : ClkMux
    port map (
            O => \N__21033\,
            I => \N__20909\
        );

    \I__4866\ : ClkMux
    port map (
            O => \N__21032\,
            I => \N__20909\
        );

    \I__4865\ : ClkMux
    port map (
            O => \N__21031\,
            I => \N__20909\
        );

    \I__4864\ : ClkMux
    port map (
            O => \N__21030\,
            I => \N__20909\
        );

    \I__4863\ : ClkMux
    port map (
            O => \N__21029\,
            I => \N__20909\
        );

    \I__4862\ : ClkMux
    port map (
            O => \N__21028\,
            I => \N__20909\
        );

    \I__4861\ : ClkMux
    port map (
            O => \N__21027\,
            I => \N__20909\
        );

    \I__4860\ : ClkMux
    port map (
            O => \N__21026\,
            I => \N__20909\
        );

    \I__4859\ : ClkMux
    port map (
            O => \N__21025\,
            I => \N__20909\
        );

    \I__4858\ : ClkMux
    port map (
            O => \N__21024\,
            I => \N__20909\
        );

    \I__4857\ : ClkMux
    port map (
            O => \N__21023\,
            I => \N__20909\
        );

    \I__4856\ : ClkMux
    port map (
            O => \N__21022\,
            I => \N__20909\
        );

    \I__4855\ : ClkMux
    port map (
            O => \N__21021\,
            I => \N__20909\
        );

    \I__4854\ : ClkMux
    port map (
            O => \N__21020\,
            I => \N__20909\
        );

    \I__4853\ : ClkMux
    port map (
            O => \N__21019\,
            I => \N__20909\
        );

    \I__4852\ : ClkMux
    port map (
            O => \N__21018\,
            I => \N__20909\
        );

    \I__4851\ : ClkMux
    port map (
            O => \N__21017\,
            I => \N__20909\
        );

    \I__4850\ : ClkMux
    port map (
            O => \N__21016\,
            I => \N__20909\
        );

    \I__4849\ : ClkMux
    port map (
            O => \N__21015\,
            I => \N__20909\
        );

    \I__4848\ : ClkMux
    port map (
            O => \N__21014\,
            I => \N__20909\
        );

    \I__4847\ : ClkMux
    port map (
            O => \N__21013\,
            I => \N__20909\
        );

    \I__4846\ : ClkMux
    port map (
            O => \N__21012\,
            I => \N__20909\
        );

    \I__4845\ : ClkMux
    port map (
            O => \N__21011\,
            I => \N__20909\
        );

    \I__4844\ : ClkMux
    port map (
            O => \N__21010\,
            I => \N__20909\
        );

    \I__4843\ : ClkMux
    port map (
            O => \N__21009\,
            I => \N__20909\
        );

    \I__4842\ : ClkMux
    port map (
            O => \N__21008\,
            I => \N__20909\
        );

    \I__4841\ : ClkMux
    port map (
            O => \N__21007\,
            I => \N__20909\
        );

    \I__4840\ : ClkMux
    port map (
            O => \N__21006\,
            I => \N__20909\
        );

    \I__4839\ : ClkMux
    port map (
            O => \N__21005\,
            I => \N__20909\
        );

    \I__4838\ : ClkMux
    port map (
            O => \N__21004\,
            I => \N__20909\
        );

    \I__4837\ : ClkMux
    port map (
            O => \N__21003\,
            I => \N__20909\
        );

    \I__4836\ : ClkMux
    port map (
            O => \N__21002\,
            I => \N__20909\
        );

    \I__4835\ : ClkMux
    port map (
            O => \N__21001\,
            I => \N__20909\
        );

    \I__4834\ : ClkMux
    port map (
            O => \N__21000\,
            I => \N__20909\
        );

    \I__4833\ : GlobalMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__4832\ : gio2CtrlBuf
    port map (
            O => \N__20906\,
            I => \TVP_CLK_c\
        );

    \I__4831\ : SRMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__20900\,
            I => \N__20896\
        );

    \I__4829\ : SRMux
    port map (
            O => \N__20899\,
            I => \N__20893\
        );

    \I__4828\ : Span4Mux_v
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__20893\,
            I => \N__20887\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__20890\,
            I => n3860
        );

    \I__4825\ : Odrv12
    port map (
            O => \N__20887\,
            I => n3860
        );

    \I__4824\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__20876\,
            I => \line_buffer.n597\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__4820\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__20867\,
            I => \N__20864\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__4817\ : Span4Mux_h
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__4816\ : Span4Mux_h
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__20855\,
            I => \line_buffer.n605\
        );

    \I__4814\ : InMux
    port map (
            O => \N__20852\,
            I => \N__20849\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__4812\ : Span4Mux_v
    port map (
            O => \N__20846\,
            I => \N__20843\
        );

    \I__4811\ : Span4Mux_h
    port map (
            O => \N__20843\,
            I => \N__20840\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__20840\,
            I => \N__20837\
        );

    \I__4809\ : Odrv4
    port map (
            O => \N__20837\,
            I => \line_buffer.n604\
        );

    \I__4808\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__4806\ : Span12Mux_v
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__4805\ : Odrv12
    port map (
            O => \N__20825\,
            I => \line_buffer.n596\
        );

    \I__4804\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20819\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__4802\ : Span4Mux_h
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__4801\ : Span4Mux_v
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__4800\ : Span4Mux_h
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__20807\,
            I => \line_buffer.n508\
        );

    \I__4798\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20801\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__20801\,
            I => \line_buffer.n3833\
        );

    \I__4796\ : CascadeMux
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20792\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__20792\,
            I => \N__20789\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__20789\,
            I => \N__20786\
        );

    \I__4792\ : Span4Mux_v
    port map (
            O => \N__20786\,
            I => \N__20783\
        );

    \I__4791\ : Sp12to4
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__4790\ : Span12Mux_h
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__4789\ : Odrv12
    port map (
            O => \N__20777\,
            I => \line_buffer.n500\
        );

    \I__4788\ : InMux
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__20771\,
            I => \line_buffer.n3836\
        );

    \I__4786\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__4784\ : Odrv12
    port map (
            O => \N__20762\,
            I => \line_buffer.n3721\
        );

    \I__4783\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__20750\,
            I => \TX_DATA_4\
        );

    \I__4779\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20743\
        );

    \I__4778\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20740\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__20743\,
            I => \N__20737\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__20740\,
            I => \transmit_module.n179\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__20737\,
            I => \transmit_module.n179\
        );

    \I__4774\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__20729\,
            I => \N__20725\
        );

    \I__4772\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20722\
        );

    \I__4771\ : Odrv4
    port map (
            O => \N__20725\,
            I => \transmit_module.n211\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__20722\,
            I => \transmit_module.n211\
        );

    \I__4769\ : SRMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__20714\,
            I => \N__20708\
        );

    \I__4767\ : SRMux
    port map (
            O => \N__20713\,
            I => \N__20705\
        );

    \I__4766\ : CascadeMux
    port map (
            O => \N__20712\,
            I => \N__20702\
        );

    \I__4765\ : SRMux
    port map (
            O => \N__20711\,
            I => \N__20687\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__20708\,
            I => \N__20676\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20676\
        );

    \I__4762\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20673\
        );

    \I__4761\ : CascadeMux
    port map (
            O => \N__20701\,
            I => \N__20670\
        );

    \I__4760\ : CascadeMux
    port map (
            O => \N__20700\,
            I => \N__20667\
        );

    \I__4759\ : IoInMux
    port map (
            O => \N__20699\,
            I => \N__20662\
        );

    \I__4758\ : SRMux
    port map (
            O => \N__20698\,
            I => \N__20657\
        );

    \I__4757\ : SRMux
    port map (
            O => \N__20697\,
            I => \N__20653\
        );

    \I__4756\ : SRMux
    port map (
            O => \N__20696\,
            I => \N__20650\
        );

    \I__4755\ : SRMux
    port map (
            O => \N__20695\,
            I => \N__20646\
        );

    \I__4754\ : SRMux
    port map (
            O => \N__20694\,
            I => \N__20643\
        );

    \I__4753\ : SRMux
    port map (
            O => \N__20693\,
            I => \N__20640\
        );

    \I__4752\ : SRMux
    port map (
            O => \N__20692\,
            I => \N__20637\
        );

    \I__4751\ : SRMux
    port map (
            O => \N__20691\,
            I => \N__20634\
        );

    \I__4750\ : SRMux
    port map (
            O => \N__20690\,
            I => \N__20631\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__20687\,
            I => \N__20627\
        );

    \I__4748\ : SRMux
    port map (
            O => \N__20686\,
            I => \N__20624\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__20685\,
            I => \N__20621\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__20684\,
            I => \N__20614\
        );

    \I__4745\ : SRMux
    port map (
            O => \N__20683\,
            I => \N__20610\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__20682\,
            I => \N__20606\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__20681\,
            I => \N__20602\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__20676\,
            I => \N__20593\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__20673\,
            I => \N__20593\
        );

    \I__4740\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20588\
        );

    \I__4739\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20588\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__20666\,
            I => \N__20584\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__20665\,
            I => \N__20581\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__20662\,
            I => \N__20578\
        );

    \I__4735\ : SRMux
    port map (
            O => \N__20661\,
            I => \N__20574\
        );

    \I__4734\ : SRMux
    port map (
            O => \N__20660\,
            I => \N__20569\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__20657\,
            I => \N__20565\
        );

    \I__4732\ : SRMux
    port map (
            O => \N__20656\,
            I => \N__20562\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__20653\,
            I => \N__20557\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__20650\,
            I => \N__20557\
        );

    \I__4729\ : SRMux
    port map (
            O => \N__20649\,
            I => \N__20554\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__20646\,
            I => \N__20545\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20545\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__20640\,
            I => \N__20545\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__20637\,
            I => \N__20545\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__20634\,
            I => \N__20540\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20631\,
            I => \N__20540\
        );

    \I__4722\ : SRMux
    port map (
            O => \N__20630\,
            I => \N__20537\
        );

    \I__4721\ : Span4Mux_h
    port map (
            O => \N__20627\,
            I => \N__20532\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__20624\,
            I => \N__20532\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20525\
        );

    \I__4718\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20525\
        );

    \I__4717\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20525\
        );

    \I__4716\ : SRMux
    port map (
            O => \N__20618\,
            I => \N__20522\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__20617\,
            I => \N__20519\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20513\
        );

    \I__4713\ : SRMux
    port map (
            O => \N__20613\,
            I => \N__20509\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__20610\,
            I => \N__20505\
        );

    \I__4711\ : SRMux
    port map (
            O => \N__20609\,
            I => \N__20502\
        );

    \I__4710\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20495\
        );

    \I__4709\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20495\
        );

    \I__4708\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20495\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__20601\,
            I => \N__20492\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__20600\,
            I => \N__20486\
        );

    \I__4705\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20481\
        );

    \I__4704\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20481\
        );

    \I__4703\ : Span4Mux_h
    port map (
            O => \N__20593\,
            I => \N__20476\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__20588\,
            I => \N__20476\
        );

    \I__4701\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20471\
        );

    \I__4700\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20471\
        );

    \I__4699\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20468\
        );

    \I__4698\ : Span4Mux_s3_h
    port map (
            O => \N__20578\,
            I => \N__20465\
        );

    \I__4697\ : SRMux
    port map (
            O => \N__20577\,
            I => \N__20462\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20459\
        );

    \I__4695\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20456\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__20572\,
            I => \N__20453\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__20569\,
            I => \N__20449\
        );

    \I__4692\ : SRMux
    port map (
            O => \N__20568\,
            I => \N__20446\
        );

    \I__4691\ : Span4Mux_v
    port map (
            O => \N__20565\,
            I => \N__20431\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__20562\,
            I => \N__20431\
        );

    \I__4689\ : Span4Mux_v
    port map (
            O => \N__20557\,
            I => \N__20431\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__20554\,
            I => \N__20431\
        );

    \I__4687\ : Span4Mux_v
    port map (
            O => \N__20545\,
            I => \N__20431\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__20540\,
            I => \N__20431\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__20537\,
            I => \N__20431\
        );

    \I__4684\ : Span4Mux_v
    port map (
            O => \N__20532\,
            I => \N__20424\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__20525\,
            I => \N__20424\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__20522\,
            I => \N__20424\
        );

    \I__4681\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20421\
        );

    \I__4680\ : SRMux
    port map (
            O => \N__20518\,
            I => \N__20418\
        );

    \I__4679\ : SRMux
    port map (
            O => \N__20517\,
            I => \N__20415\
        );

    \I__4678\ : SRMux
    port map (
            O => \N__20516\,
            I => \N__20412\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__20513\,
            I => \N__20409\
        );

    \I__4676\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20406\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__20509\,
            I => \N__20403\
        );

    \I__4674\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20400\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__20505\,
            I => \N__20395\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__20502\,
            I => \N__20395\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__20495\,
            I => \N__20392\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20385\
        );

    \I__4669\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20385\
        );

    \I__4668\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20385\
        );

    \I__4667\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20378\
        );

    \I__4666\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20378\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__20481\,
            I => \N__20369\
        );

    \I__4664\ : Span4Mux_h
    port map (
            O => \N__20476\,
            I => \N__20369\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__20471\,
            I => \N__20369\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20369\
        );

    \I__4661\ : Sp12to4
    port map (
            O => \N__20465\,
            I => \N__20363\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20360\
        );

    \I__4659\ : Span4Mux_v
    port map (
            O => \N__20459\,
            I => \N__20357\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__20456\,
            I => \N__20354\
        );

    \I__4657\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20349\
        );

    \I__4656\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20349\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__20449\,
            I => \N__20342\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20342\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__20431\,
            I => \N__20342\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__20424\,
            I => \N__20337\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__20421\,
            I => \N__20337\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__20418\,
            I => \N__20328\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__20415\,
            I => \N__20328\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__20412\,
            I => \N__20328\
        );

    \I__4647\ : Span4Mux_v
    port map (
            O => \N__20409\,
            I => \N__20328\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__20406\,
            I => \N__20315\
        );

    \I__4645\ : Span4Mux_v
    port map (
            O => \N__20403\,
            I => \N__20315\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__20400\,
            I => \N__20315\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__20395\,
            I => \N__20315\
        );

    \I__4642\ : Span4Mux_h
    port map (
            O => \N__20392\,
            I => \N__20315\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__20385\,
            I => \N__20315\
        );

    \I__4640\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20310\
        );

    \I__4639\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20310\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__20378\,
            I => \N__20305\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__20369\,
            I => \N__20305\
        );

    \I__4636\ : SRMux
    port map (
            O => \N__20368\,
            I => \N__20302\
        );

    \I__4635\ : SRMux
    port map (
            O => \N__20367\,
            I => \N__20299\
        );

    \I__4634\ : SRMux
    port map (
            O => \N__20366\,
            I => \N__20296\
        );

    \I__4633\ : Span12Mux_v
    port map (
            O => \N__20363\,
            I => \N__20291\
        );

    \I__4632\ : Span12Mux_v
    port map (
            O => \N__20360\,
            I => \N__20291\
        );

    \I__4631\ : Span4Mux_h
    port map (
            O => \N__20357\,
            I => \N__20284\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__20354\,
            I => \N__20284\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__20349\,
            I => \N__20284\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__20342\,
            I => \N__20277\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__20337\,
            I => \N__20277\
        );

    \I__4626\ : Span4Mux_v
    port map (
            O => \N__20328\,
            I => \N__20277\
        );

    \I__4625\ : Span4Mux_v
    port map (
            O => \N__20315\,
            I => \N__20270\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__20310\,
            I => \N__20270\
        );

    \I__4623\ : Span4Mux_h
    port map (
            O => \N__20305\,
            I => \N__20270\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__20302\,
            I => \ADV_VSYNC_c\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__20299\,
            I => \ADV_VSYNC_c\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__20296\,
            I => \ADV_VSYNC_c\
        );

    \I__4619\ : Odrv12
    port map (
            O => \N__20291\,
            I => \ADV_VSYNC_c\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__20284\,
            I => \ADV_VSYNC_c\
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__20277\,
            I => \ADV_VSYNC_c\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__20270\,
            I => \ADV_VSYNC_c\
        );

    \I__4615\ : InMux
    port map (
            O => \N__20255\,
            I => \N__20246\
        );

    \I__4614\ : InMux
    port map (
            O => \N__20254\,
            I => \N__20241\
        );

    \I__4613\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20241\
        );

    \I__4612\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20229\
        );

    \I__4611\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20222\
        );

    \I__4610\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20222\
        );

    \I__4609\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20222\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__20246\,
            I => \N__20217\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__20241\,
            I => \N__20217\
        );

    \I__4606\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20212\
        );

    \I__4605\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20212\
        );

    \I__4604\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20207\
        );

    \I__4603\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20207\
        );

    \I__4602\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20197\
        );

    \I__4601\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20197\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20197\
        );

    \I__4599\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20197\
        );

    \I__4598\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20190\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__20229\,
            I => \N__20187\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__20222\,
            I => \N__20180\
        );

    \I__4595\ : Span4Mux_h
    port map (
            O => \N__20217\,
            I => \N__20180\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__20212\,
            I => \N__20180\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__20207\,
            I => \N__20175\
        );

    \I__4592\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20172\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__20197\,
            I => \N__20169\
        );

    \I__4590\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20160\
        );

    \I__4589\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20160\
        );

    \I__4588\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20160\
        );

    \I__4587\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20160\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__20190\,
            I => \N__20157\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__20187\,
            I => \N__20152\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__20180\,
            I => \N__20152\
        );

    \I__4583\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20147\
        );

    \I__4582\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20147\
        );

    \I__4581\ : Span4Mux_h
    port map (
            O => \N__20175\,
            I => \N__20136\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20136\
        );

    \I__4579\ : Span4Mux_v
    port map (
            O => \N__20169\,
            I => \N__20136\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20136\
        );

    \I__4577\ : Span4Mux_h
    port map (
            O => \N__20157\,
            I => \N__20136\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__20152\,
            I => \transmit_module.n3853\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__20147\,
            I => \transmit_module.n3853\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__20136\,
            I => \transmit_module.n3853\
        );

    \I__4573\ : CascadeMux
    port map (
            O => \N__20129\,
            I => \N__20125\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__20128\,
            I => \N__20122\
        );

    \I__4571\ : CascadeBuf
    port map (
            O => \N__20125\,
            I => \N__20119\
        );

    \I__4570\ : CascadeBuf
    port map (
            O => \N__20122\,
            I => \N__20116\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__20119\,
            I => \N__20113\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__20116\,
            I => \N__20110\
        );

    \I__4567\ : CascadeBuf
    port map (
            O => \N__20113\,
            I => \N__20107\
        );

    \I__4566\ : CascadeBuf
    port map (
            O => \N__20110\,
            I => \N__20104\
        );

    \I__4565\ : CascadeMux
    port map (
            O => \N__20107\,
            I => \N__20101\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__20104\,
            I => \N__20098\
        );

    \I__4563\ : CascadeBuf
    port map (
            O => \N__20101\,
            I => \N__20095\
        );

    \I__4562\ : CascadeBuf
    port map (
            O => \N__20098\,
            I => \N__20092\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__20095\,
            I => \N__20089\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__20092\,
            I => \N__20086\
        );

    \I__4559\ : CascadeBuf
    port map (
            O => \N__20089\,
            I => \N__20083\
        );

    \I__4558\ : CascadeBuf
    port map (
            O => \N__20086\,
            I => \N__20080\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__20083\,
            I => \N__20077\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__20080\,
            I => \N__20074\
        );

    \I__4555\ : CascadeBuf
    port map (
            O => \N__20077\,
            I => \N__20071\
        );

    \I__4554\ : CascadeBuf
    port map (
            O => \N__20074\,
            I => \N__20068\
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__20071\,
            I => \N__20065\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__20068\,
            I => \N__20062\
        );

    \I__4551\ : CascadeBuf
    port map (
            O => \N__20065\,
            I => \N__20059\
        );

    \I__4550\ : CascadeBuf
    port map (
            O => \N__20062\,
            I => \N__20056\
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__20059\,
            I => \N__20053\
        );

    \I__4548\ : CascadeMux
    port map (
            O => \N__20056\,
            I => \N__20050\
        );

    \I__4547\ : CascadeBuf
    port map (
            O => \N__20053\,
            I => \N__20047\
        );

    \I__4546\ : CascadeBuf
    port map (
            O => \N__20050\,
            I => \N__20044\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__20047\,
            I => \N__20041\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__20044\,
            I => \N__20038\
        );

    \I__4543\ : CascadeBuf
    port map (
            O => \N__20041\,
            I => \N__20035\
        );

    \I__4542\ : CascadeBuf
    port map (
            O => \N__20038\,
            I => \N__20032\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__20035\,
            I => \N__20029\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__20032\,
            I => \N__20026\
        );

    \I__4539\ : CascadeBuf
    port map (
            O => \N__20029\,
            I => \N__20023\
        );

    \I__4538\ : CascadeBuf
    port map (
            O => \N__20026\,
            I => \N__20020\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__20023\,
            I => \N__20017\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__20020\,
            I => \N__20014\
        );

    \I__4535\ : CascadeBuf
    port map (
            O => \N__20017\,
            I => \N__20011\
        );

    \I__4534\ : CascadeBuf
    port map (
            O => \N__20014\,
            I => \N__20008\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__20011\,
            I => \N__20005\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__20008\,
            I => \N__20002\
        );

    \I__4531\ : CascadeBuf
    port map (
            O => \N__20005\,
            I => \N__19999\
        );

    \I__4530\ : CascadeBuf
    port map (
            O => \N__20002\,
            I => \N__19996\
        );

    \I__4529\ : CascadeMux
    port map (
            O => \N__19999\,
            I => \N__19993\
        );

    \I__4528\ : CascadeMux
    port map (
            O => \N__19996\,
            I => \N__19990\
        );

    \I__4527\ : CascadeBuf
    port map (
            O => \N__19993\,
            I => \N__19987\
        );

    \I__4526\ : CascadeBuf
    port map (
            O => \N__19990\,
            I => \N__19984\
        );

    \I__4525\ : CascadeMux
    port map (
            O => \N__19987\,
            I => \N__19981\
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__19984\,
            I => \N__19978\
        );

    \I__4523\ : CascadeBuf
    port map (
            O => \N__19981\,
            I => \N__19975\
        );

    \I__4522\ : CascadeBuf
    port map (
            O => \N__19978\,
            I => \N__19972\
        );

    \I__4521\ : CascadeMux
    port map (
            O => \N__19975\,
            I => \N__19969\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__19972\,
            I => \N__19966\
        );

    \I__4519\ : CascadeBuf
    port map (
            O => \N__19969\,
            I => \N__19963\
        );

    \I__4518\ : CascadeBuf
    port map (
            O => \N__19966\,
            I => \N__19960\
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__19963\,
            I => \N__19957\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__19960\,
            I => \N__19954\
        );

    \I__4515\ : CascadeBuf
    port map (
            O => \N__19957\,
            I => \N__19951\
        );

    \I__4514\ : CascadeBuf
    port map (
            O => \N__19954\,
            I => \N__19948\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__19951\,
            I => \N__19945\
        );

    \I__4512\ : CascadeMux
    port map (
            O => \N__19948\,
            I => \N__19942\
        );

    \I__4511\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19939\
        );

    \I__4510\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19936\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__19939\,
            I => \N__19933\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19936\,
            I => \N__19930\
        );

    \I__4507\ : Span12Mux_h
    port map (
            O => \N__19933\,
            I => \N__19927\
        );

    \I__4506\ : Span12Mux_s11_h
    port map (
            O => \N__19930\,
            I => \N__19924\
        );

    \I__4505\ : Span12Mux_v
    port map (
            O => \N__19927\,
            I => \N__19921\
        );

    \I__4504\ : Span12Mux_v
    port map (
            O => \N__19924\,
            I => \N__19918\
        );

    \I__4503\ : Odrv12
    port map (
            O => \N__19921\,
            I => n19
        );

    \I__4502\ : Odrv12
    port map (
            O => \N__19918\,
            I => n19
        );

    \I__4501\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19907\
        );

    \I__4500\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19907\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19903\
        );

    \I__4498\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19900\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__19903\,
            I => \N__19897\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__19900\,
            I => \N__19894\
        );

    \I__4495\ : Span4Mux_h
    port map (
            O => \N__19897\,
            I => \N__19891\
        );

    \I__4494\ : Span4Mux_h
    port map (
            O => \N__19894\,
            I => \N__19888\
        );

    \I__4493\ : Span4Mux_h
    port map (
            O => \N__19891\,
            I => \N__19883\
        );

    \I__4492\ : Span4Mux_v
    port map (
            O => \N__19888\,
            I => \N__19883\
        );

    \I__4491\ : Odrv4
    port map (
            O => \N__19883\,
            I => \TVP_HSYNC_c\
        );

    \I__4490\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__19877\,
            I => \receive_module.rx_counter.n10\
        );

    \I__4488\ : InMux
    port map (
            O => \N__19874\,
            I => \bfn_17_9_0_\
        );

    \I__4487\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__19868\,
            I => \receive_module.rx_counter.n9\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19865\,
            I => \receive_module.rx_counter.n3357\
        );

    \I__4484\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19859\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__19859\,
            I => \receive_module.rx_counter.n8\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19856\,
            I => \receive_module.rx_counter.n3358\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19849\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19846\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19849\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__19846\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19841\,
            I => \receive_module.rx_counter.n3359\
        );

    \I__4476\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19834\
        );

    \I__4475\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__19834\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__19831\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19826\,
            I => \receive_module.rx_counter.n3360\
        );

    \I__4471\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19819\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19816\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__19819\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19816\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__4467\ : InMux
    port map (
            O => \N__19811\,
            I => \receive_module.rx_counter.n3361\
        );

    \I__4466\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19803\
        );

    \I__4465\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19798\
        );

    \I__4464\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19798\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__19803\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__19798\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__4461\ : InMux
    port map (
            O => \N__19793\,
            I => \receive_module.rx_counter.n3362\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__19790\,
            I => \transmit_module.n210_cascade_\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__4458\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__19778\,
            I => \transmit_module.n201\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__19775\,
            I => \transmit_module.n217_cascade_\
        );

    \I__4454\ : InMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__19769\,
            I => \N__19765\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19760\
        );

    \I__4451\ : Span4Mux_h
    port map (
            O => \N__19765\,
            I => \N__19757\
        );

    \I__4450\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19754\
        );

    \I__4449\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19751\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19748\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__19757\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__19754\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__19751\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__19748\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__4443\ : CascadeMux
    port map (
            O => \N__19739\,
            I => \N__19734\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__19738\,
            I => \N__19731\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__19737\,
            I => \N__19724\
        );

    \I__4440\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19716\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19716\
        );

    \I__4438\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19709\
        );

    \I__4437\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19709\
        );

    \I__4436\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19709\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__19727\,
            I => \N__19704\
        );

    \I__4434\ : InMux
    port map (
            O => \N__19724\,
            I => \N__19701\
        );

    \I__4433\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19698\
        );

    \I__4432\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19693\
        );

    \I__4431\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19693\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__19716\,
            I => \N__19688\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__19709\,
            I => \N__19688\
        );

    \I__4428\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19685\
        );

    \I__4427\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19682\
        );

    \I__4426\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19679\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__19701\,
            I => \N__19674\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19674\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__19693\,
            I => \N__19669\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__19688\,
            I => \N__19669\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__19685\,
            I => \transmit_module.n3855\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__19682\,
            I => \transmit_module.n3855\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__19679\,
            I => \transmit_module.n3855\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__19674\,
            I => \transmit_module.n3855\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__19669\,
            I => \transmit_module.n3855\
        );

    \I__4416\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__4414\ : Span4Mux_v
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__19649\,
            I => \transmit_module.n195\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__4409\ : Span4Mux_h
    port map (
            O => \N__19637\,
            I => \N__19631\
        );

    \I__4408\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19628\
        );

    \I__4407\ : InMux
    port map (
            O => \N__19635\,
            I => \N__19623\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19623\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__19631\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__19628\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19623\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19610\
        );

    \I__4401\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19610\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19602\
        );

    \I__4399\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19597\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19608\,
            I => \N__19597\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19594\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19586\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19583\
        );

    \I__4394\ : Span4Mux_v
    port map (
            O => \N__19602\,
            I => \N__19576\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__19597\,
            I => \N__19576\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__19594\,
            I => \N__19576\
        );

    \I__4391\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19569\
        );

    \I__4390\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19569\
        );

    \I__4389\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19569\
        );

    \I__4388\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19564\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19561\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__19586\,
            I => \N__19558\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19583\,
            I => \N__19555\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__19576\,
            I => \N__19550\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__19569\,
            I => \N__19550\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19537\
        );

    \I__4381\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19537\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__19564\,
            I => \N__19530\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__19561\,
            I => \N__19530\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__19558\,
            I => \N__19530\
        );

    \I__4377\ : Span4Mux_v
    port map (
            O => \N__19555\,
            I => \N__19525\
        );

    \I__4376\ : Span4Mux_v
    port map (
            O => \N__19550\,
            I => \N__19525\
        );

    \I__4375\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19516\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19516\
        );

    \I__4373\ : InMux
    port map (
            O => \N__19547\,
            I => \N__19516\
        );

    \I__4372\ : InMux
    port map (
            O => \N__19546\,
            I => \N__19516\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19507\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19507\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19507\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19542\,
            I => \N__19507\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__19537\,
            I => \transmit_module.n3549\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__19530\,
            I => \transmit_module.n3549\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__19525\,
            I => \transmit_module.n3549\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19516\,
            I => \transmit_module.n3549\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19507\,
            I => \transmit_module.n3549\
        );

    \I__4362\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__19493\,
            I => \transmit_module.n217\
        );

    \I__4360\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19486\
        );

    \I__4359\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19483\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__19486\,
            I => \transmit_module.n185\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__19483\,
            I => \transmit_module.n185\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__19478\,
            I => \N__19474\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__19477\,
            I => \N__19471\
        );

    \I__4354\ : CascadeBuf
    port map (
            O => \N__19474\,
            I => \N__19468\
        );

    \I__4353\ : CascadeBuf
    port map (
            O => \N__19471\,
            I => \N__19465\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__19468\,
            I => \N__19462\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__19465\,
            I => \N__19459\
        );

    \I__4350\ : CascadeBuf
    port map (
            O => \N__19462\,
            I => \N__19456\
        );

    \I__4349\ : CascadeBuf
    port map (
            O => \N__19459\,
            I => \N__19453\
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__19456\,
            I => \N__19450\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__19453\,
            I => \N__19447\
        );

    \I__4346\ : CascadeBuf
    port map (
            O => \N__19450\,
            I => \N__19444\
        );

    \I__4345\ : CascadeBuf
    port map (
            O => \N__19447\,
            I => \N__19441\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__19444\,
            I => \N__19438\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__4342\ : CascadeBuf
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__4341\ : CascadeBuf
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__4340\ : CascadeMux
    port map (
            O => \N__19432\,
            I => \N__19426\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__19429\,
            I => \N__19423\
        );

    \I__4338\ : CascadeBuf
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__4337\ : CascadeBuf
    port map (
            O => \N__19423\,
            I => \N__19417\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__19420\,
            I => \N__19414\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__19417\,
            I => \N__19411\
        );

    \I__4334\ : CascadeBuf
    port map (
            O => \N__19414\,
            I => \N__19408\
        );

    \I__4333\ : CascadeBuf
    port map (
            O => \N__19411\,
            I => \N__19405\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__19408\,
            I => \N__19402\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__19405\,
            I => \N__19399\
        );

    \I__4330\ : CascadeBuf
    port map (
            O => \N__19402\,
            I => \N__19396\
        );

    \I__4329\ : CascadeBuf
    port map (
            O => \N__19399\,
            I => \N__19393\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__19396\,
            I => \N__19390\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__19393\,
            I => \N__19387\
        );

    \I__4326\ : CascadeBuf
    port map (
            O => \N__19390\,
            I => \N__19384\
        );

    \I__4325\ : CascadeBuf
    port map (
            O => \N__19387\,
            I => \N__19381\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__19384\,
            I => \N__19378\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__19381\,
            I => \N__19375\
        );

    \I__4322\ : CascadeBuf
    port map (
            O => \N__19378\,
            I => \N__19372\
        );

    \I__4321\ : CascadeBuf
    port map (
            O => \N__19375\,
            I => \N__19369\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__19372\,
            I => \N__19366\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__4318\ : CascadeBuf
    port map (
            O => \N__19366\,
            I => \N__19360\
        );

    \I__4317\ : CascadeBuf
    port map (
            O => \N__19363\,
            I => \N__19357\
        );

    \I__4316\ : CascadeMux
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__19357\,
            I => \N__19351\
        );

    \I__4314\ : CascadeBuf
    port map (
            O => \N__19354\,
            I => \N__19348\
        );

    \I__4313\ : CascadeBuf
    port map (
            O => \N__19351\,
            I => \N__19345\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__19348\,
            I => \N__19342\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__19345\,
            I => \N__19339\
        );

    \I__4310\ : CascadeBuf
    port map (
            O => \N__19342\,
            I => \N__19336\
        );

    \I__4309\ : CascadeBuf
    port map (
            O => \N__19339\,
            I => \N__19333\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__19336\,
            I => \N__19330\
        );

    \I__4307\ : CascadeMux
    port map (
            O => \N__19333\,
            I => \N__19327\
        );

    \I__4306\ : CascadeBuf
    port map (
            O => \N__19330\,
            I => \N__19324\
        );

    \I__4305\ : CascadeBuf
    port map (
            O => \N__19327\,
            I => \N__19321\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__19324\,
            I => \N__19318\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__19321\,
            I => \N__19315\
        );

    \I__4302\ : CascadeBuf
    port map (
            O => \N__19318\,
            I => \N__19312\
        );

    \I__4301\ : CascadeBuf
    port map (
            O => \N__19315\,
            I => \N__19309\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__19312\,
            I => \N__19306\
        );

    \I__4299\ : CascadeMux
    port map (
            O => \N__19309\,
            I => \N__19303\
        );

    \I__4298\ : CascadeBuf
    port map (
            O => \N__19306\,
            I => \N__19300\
        );

    \I__4297\ : CascadeBuf
    port map (
            O => \N__19303\,
            I => \N__19297\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__19300\,
            I => \N__19294\
        );

    \I__4295\ : CascadeMux
    port map (
            O => \N__19297\,
            I => \N__19291\
        );

    \I__4294\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19288\
        );

    \I__4293\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19285\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__19288\,
            I => \N__19282\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__19285\,
            I => \N__19279\
        );

    \I__4290\ : Span4Mux_h
    port map (
            O => \N__19282\,
            I => \N__19276\
        );

    \I__4289\ : Span4Mux_h
    port map (
            O => \N__19279\,
            I => \N__19273\
        );

    \I__4288\ : Sp12to4
    port map (
            O => \N__19276\,
            I => \N__19270\
        );

    \I__4287\ : Sp12to4
    port map (
            O => \N__19273\,
            I => \N__19267\
        );

    \I__4286\ : Span12Mux_v
    port map (
            O => \N__19270\,
            I => \N__19262\
        );

    \I__4285\ : Span12Mux_v
    port map (
            O => \N__19267\,
            I => \N__19262\
        );

    \I__4284\ : Odrv12
    port map (
            O => \N__19262\,
            I => n25
        );

    \I__4283\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19254\
        );

    \I__4282\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19246\
        );

    \I__4281\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19242\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__19254\,
            I => \N__19239\
        );

    \I__4279\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19236\
        );

    \I__4278\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19233\
        );

    \I__4277\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19228\
        );

    \I__4276\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19228\
        );

    \I__4275\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19223\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__19246\,
            I => \N__19218\
        );

    \I__4273\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19215\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__19242\,
            I => \N__19212\
        );

    \I__4271\ : Span4Mux_h
    port map (
            O => \N__19239\,
            I => \N__19207\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19207\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19202\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__19228\,
            I => \N__19202\
        );

    \I__4267\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19197\
        );

    \I__4266\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19197\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__19223\,
            I => \N__19194\
        );

    \I__4264\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19189\
        );

    \I__4263\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19189\
        );

    \I__4262\ : Sp12to4
    port map (
            O => \N__19218\,
            I => \N__19183\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__19215\,
            I => \N__19183\
        );

    \I__4260\ : Span4Mux_v
    port map (
            O => \N__19212\,
            I => \N__19180\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__19207\,
            I => \N__19177\
        );

    \I__4258\ : Span4Mux_v
    port map (
            O => \N__19202\,
            I => \N__19172\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__19197\,
            I => \N__19172\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__19194\,
            I => \N__19167\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19167\
        );

    \I__4254\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19164\
        );

    \I__4253\ : Span12Mux_v
    port map (
            O => \N__19183\,
            I => \N__19161\
        );

    \I__4252\ : Span4Mux_v
    port map (
            O => \N__19180\,
            I => \N__19158\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__19177\,
            I => \N__19155\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__19172\,
            I => \N__19150\
        );

    \I__4249\ : Span4Mux_v
    port map (
            O => \N__19167\,
            I => \N__19150\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__19164\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4247\ : Odrv12
    port map (
            O => \N__19161\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__19158\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__19155\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__19150\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4243\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__19136\,
            I => \transmit_module.ADDR_Y_COMPONENT_10\
        );

    \I__4241\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19129\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__19132\,
            I => \N__19124\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__19129\,
            I => \N__19121\
        );

    \I__4238\ : InMux
    port map (
            O => \N__19128\,
            I => \N__19118\
        );

    \I__4237\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19115\
        );

    \I__4236\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19112\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__19121\,
            I => \N__19109\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__19118\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__19115\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__19112\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__4231\ : Odrv4
    port map (
            O => \N__19109\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__4230\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__19097\,
            I => \transmit_module.n178\
        );

    \I__4228\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__19091\,
            I => \transmit_module.n210\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__19088\,
            I => \transmit_module.n178_cascade_\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__4224\ : CascadeBuf
    port map (
            O => \N__19082\,
            I => \N__19078\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__19081\,
            I => \N__19075\
        );

    \I__4222\ : CascadeMux
    port map (
            O => \N__19078\,
            I => \N__19072\
        );

    \I__4221\ : CascadeBuf
    port map (
            O => \N__19075\,
            I => \N__19069\
        );

    \I__4220\ : CascadeBuf
    port map (
            O => \N__19072\,
            I => \N__19066\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__19069\,
            I => \N__19063\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__19066\,
            I => \N__19060\
        );

    \I__4217\ : CascadeBuf
    port map (
            O => \N__19063\,
            I => \N__19057\
        );

    \I__4216\ : CascadeBuf
    port map (
            O => \N__19060\,
            I => \N__19054\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__19057\,
            I => \N__19051\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__19054\,
            I => \N__19048\
        );

    \I__4213\ : CascadeBuf
    port map (
            O => \N__19051\,
            I => \N__19045\
        );

    \I__4212\ : CascadeBuf
    port map (
            O => \N__19048\,
            I => \N__19042\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__19045\,
            I => \N__19039\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__19042\,
            I => \N__19036\
        );

    \I__4209\ : CascadeBuf
    port map (
            O => \N__19039\,
            I => \N__19033\
        );

    \I__4208\ : CascadeBuf
    port map (
            O => \N__19036\,
            I => \N__19030\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__19033\,
            I => \N__19027\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__19030\,
            I => \N__19024\
        );

    \I__4205\ : CascadeBuf
    port map (
            O => \N__19027\,
            I => \N__19021\
        );

    \I__4204\ : CascadeBuf
    port map (
            O => \N__19024\,
            I => \N__19018\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__19021\,
            I => \N__19015\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__19018\,
            I => \N__19012\
        );

    \I__4201\ : CascadeBuf
    port map (
            O => \N__19015\,
            I => \N__19009\
        );

    \I__4200\ : CascadeBuf
    port map (
            O => \N__19012\,
            I => \N__19006\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__19009\,
            I => \N__19003\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__19006\,
            I => \N__19000\
        );

    \I__4197\ : CascadeBuf
    port map (
            O => \N__19003\,
            I => \N__18997\
        );

    \I__4196\ : CascadeBuf
    port map (
            O => \N__19000\,
            I => \N__18994\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__18997\,
            I => \N__18991\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__18994\,
            I => \N__18988\
        );

    \I__4193\ : CascadeBuf
    port map (
            O => \N__18991\,
            I => \N__18985\
        );

    \I__4192\ : CascadeBuf
    port map (
            O => \N__18988\,
            I => \N__18982\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__18985\,
            I => \N__18979\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__18982\,
            I => \N__18976\
        );

    \I__4189\ : CascadeBuf
    port map (
            O => \N__18979\,
            I => \N__18973\
        );

    \I__4188\ : CascadeBuf
    port map (
            O => \N__18976\,
            I => \N__18970\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__18973\,
            I => \N__18967\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__18970\,
            I => \N__18964\
        );

    \I__4185\ : CascadeBuf
    port map (
            O => \N__18967\,
            I => \N__18961\
        );

    \I__4184\ : CascadeBuf
    port map (
            O => \N__18964\,
            I => \N__18958\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__18961\,
            I => \N__18955\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__18958\,
            I => \N__18952\
        );

    \I__4181\ : CascadeBuf
    port map (
            O => \N__18955\,
            I => \N__18949\
        );

    \I__4180\ : CascadeBuf
    port map (
            O => \N__18952\,
            I => \N__18946\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__18949\,
            I => \N__18943\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__18946\,
            I => \N__18940\
        );

    \I__4177\ : CascadeBuf
    port map (
            O => \N__18943\,
            I => \N__18937\
        );

    \I__4176\ : CascadeBuf
    port map (
            O => \N__18940\,
            I => \N__18934\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__18937\,
            I => \N__18931\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__18934\,
            I => \N__18928\
        );

    \I__4173\ : CascadeBuf
    port map (
            O => \N__18931\,
            I => \N__18925\
        );

    \I__4172\ : CascadeBuf
    port map (
            O => \N__18928\,
            I => \N__18922\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__18925\,
            I => \N__18919\
        );

    \I__4170\ : CascadeMux
    port map (
            O => \N__18922\,
            I => \N__18916\
        );

    \I__4169\ : CascadeBuf
    port map (
            O => \N__18919\,
            I => \N__18913\
        );

    \I__4168\ : CascadeBuf
    port map (
            O => \N__18916\,
            I => \N__18910\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__18913\,
            I => \N__18907\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__18910\,
            I => \N__18904\
        );

    \I__4165\ : CascadeBuf
    port map (
            O => \N__18907\,
            I => \N__18901\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18904\,
            I => \N__18898\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__18901\,
            I => \N__18895\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18892\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18895\,
            I => \N__18889\
        );

    \I__4160\ : Span12Mux_h
    port map (
            O => \N__18892\,
            I => \N__18886\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__18889\,
            I => \N__18883\
        );

    \I__4158\ : Span12Mux_v
    port map (
            O => \N__18886\,
            I => \N__18878\
        );

    \I__4157\ : Span12Mux_v
    port map (
            O => \N__18883\,
            I => \N__18878\
        );

    \I__4156\ : Odrv12
    port map (
            O => \N__18878\,
            I => n18
        );

    \I__4155\ : IoInMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__4153\ : Span4Mux_s0_v
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__18866\,
            I => \GB_BUFFER_TVP_CLK_c_THRU_CO\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__18863\,
            I => \receive_module.rx_counter.n3547_cascade_\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__18857\,
            I => \receive_module.rx_counter.n3547\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__18854\,
            I => \receive_module.rx_counter.n3646_cascade_\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18848\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__18848\,
            I => \receive_module.rx_counter.n3613\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__18839\,
            I => \receive_module.rx_counter.n28\
        );

    \I__4142\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__4140\ : Span4Mux_h
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__4139\ : Sp12to4
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__4138\ : Span12Mux_v
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__4137\ : Odrv12
    port map (
            O => \N__18821\,
            I => \line_buffer.n629\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__4133\ : Odrv12
    port map (
            O => \N__18809\,
            I => \line_buffer.n637\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__4130\ : Span4Mux_v
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__4129\ : Span4Mux_h
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__4127\ : Odrv4
    port map (
            O => \N__18791\,
            I => \line_buffer.n565\
        );

    \I__4126\ : CascadeMux
    port map (
            O => \N__18788\,
            I => \line_buffer.n3761_cascade_\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4123\ : Span4Mux_h
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__4122\ : Sp12to4
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__4121\ : Span12Mux_v
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__4120\ : Odrv12
    port map (
            O => \N__18770\,
            I => \line_buffer.n573\
        );

    \I__4119\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__18764\,
            I => \line_buffer.n3764\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__4115\ : Span4Mux_h
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__18752\,
            I => \TX_DATA_5\
        );

    \I__4113\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__18746\,
            I => \transmit_module.Y_DELTA_PATTERN_33\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__4109\ : Span12Mux_v
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__4108\ : Odrv12
    port map (
            O => \N__18734\,
            I => \transmit_module.Y_DELTA_PATTERN_32\
        );

    \I__4107\ : CEMux
    port map (
            O => \N__18731\,
            I => \N__18727\
        );

    \I__4106\ : CEMux
    port map (
            O => \N__18730\,
            I => \N__18721\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18727\,
            I => \N__18717\
        );

    \I__4104\ : CEMux
    port map (
            O => \N__18726\,
            I => \N__18714\
        );

    \I__4103\ : CEMux
    port map (
            O => \N__18725\,
            I => \N__18709\
        );

    \I__4102\ : SRMux
    port map (
            O => \N__18724\,
            I => \N__18704\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__18721\,
            I => \N__18698\
        );

    \I__4100\ : CEMux
    port map (
            O => \N__18720\,
            I => \N__18695\
        );

    \I__4099\ : Span4Mux_h
    port map (
            O => \N__18717\,
            I => \N__18688\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__18714\,
            I => \N__18688\
        );

    \I__4097\ : CEMux
    port map (
            O => \N__18713\,
            I => \N__18685\
        );

    \I__4096\ : CEMux
    port map (
            O => \N__18712\,
            I => \N__18682\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18709\,
            I => \N__18679\
        );

    \I__4094\ : CEMux
    port map (
            O => \N__18708\,
            I => \N__18676\
        );

    \I__4093\ : CEMux
    port map (
            O => \N__18707\,
            I => \N__18673\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__18704\,
            I => \N__18670\
        );

    \I__4091\ : SRMux
    port map (
            O => \N__18703\,
            I => \N__18667\
        );

    \I__4090\ : SRMux
    port map (
            O => \N__18702\,
            I => \N__18664\
        );

    \I__4089\ : SRMux
    port map (
            O => \N__18701\,
            I => \N__18661\
        );

    \I__4088\ : Span4Mux_h
    port map (
            O => \N__18698\,
            I => \N__18656\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18695\,
            I => \N__18656\
        );

    \I__4086\ : SRMux
    port map (
            O => \N__18694\,
            I => \N__18653\
        );

    \I__4085\ : SRMux
    port map (
            O => \N__18693\,
            I => \N__18650\
        );

    \I__4084\ : Span4Mux_v
    port map (
            O => \N__18688\,
            I => \N__18647\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__18685\,
            I => \N__18644\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__18682\,
            I => \N__18641\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__18679\,
            I => \N__18638\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18676\,
            I => \N__18635\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__18673\,
            I => \N__18632\
        );

    \I__4078\ : Span4Mux_h
    port map (
            O => \N__18670\,
            I => \N__18627\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__18667\,
            I => \N__18627\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__18664\,
            I => \N__18624\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__18661\,
            I => \N__18621\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__18656\,
            I => \N__18618\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__18653\,
            I => \N__18613\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__18650\,
            I => \N__18613\
        );

    \I__4071\ : Span4Mux_h
    port map (
            O => \N__18647\,
            I => \N__18610\
        );

    \I__4070\ : Span4Mux_h
    port map (
            O => \N__18644\,
            I => \N__18603\
        );

    \I__4069\ : Span4Mux_v
    port map (
            O => \N__18641\,
            I => \N__18603\
        );

    \I__4068\ : Span4Mux_h
    port map (
            O => \N__18638\,
            I => \N__18603\
        );

    \I__4067\ : Span4Mux_h
    port map (
            O => \N__18635\,
            I => \N__18598\
        );

    \I__4066\ : Span4Mux_v
    port map (
            O => \N__18632\,
            I => \N__18598\
        );

    \I__4065\ : Span4Mux_v
    port map (
            O => \N__18627\,
            I => \N__18595\
        );

    \I__4064\ : Span4Mux_v
    port map (
            O => \N__18624\,
            I => \N__18592\
        );

    \I__4063\ : Span12Mux_s11_h
    port map (
            O => \N__18621\,
            I => \N__18589\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__18618\,
            I => \N__18584\
        );

    \I__4061\ : Span4Mux_v
    port map (
            O => \N__18613\,
            I => \N__18584\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__18610\,
            I => \transmit_module.n3864\
        );

    \I__4059\ : Odrv4
    port map (
            O => \N__18603\,
            I => \transmit_module.n3864\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__18598\,
            I => \transmit_module.n3864\
        );

    \I__4057\ : Odrv4
    port map (
            O => \N__18595\,
            I => \transmit_module.n3864\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__18592\,
            I => \transmit_module.n3864\
        );

    \I__4055\ : Odrv12
    port map (
            O => \N__18589\,
            I => \transmit_module.n3864\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__18584\,
            I => \transmit_module.n3864\
        );

    \I__4053\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__4051\ : Span4Mux_h
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__4050\ : Span4Mux_v
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__18554\,
            I => \line_buffer.n607\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__4045\ : Span4Mux_v
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__4044\ : Sp12to4
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__4043\ : Span12Mux_v
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__4042\ : Odrv12
    port map (
            O => \N__18536\,
            I => \line_buffer.n599\
        );

    \I__4041\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__18530\,
            I => \line_buffer.n3718\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__4037\ : Span4Mux_h
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__18518\,
            I => \transmit_module.n194\
        );

    \I__4035\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__4033\ : Span4Mux_v
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__4032\ : Span4Mux_h
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__18503\,
            I => \line_buffer.n575\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__4028\ : Span4Mux_v
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__4027\ : Sp12to4
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__4026\ : Span12Mux_h
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__4025\ : Span12Mux_v
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__4024\ : Odrv12
    port map (
            O => \N__18482\,
            I => \line_buffer.n567\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__18476\,
            I => \line_buffer.n3702\
        );

    \I__4021\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__18470\,
            I => \transmit_module.ADDR_Y_COMPONENT_3\
        );

    \I__4019\ : CEMux
    port map (
            O => \N__18467\,
            I => \N__18463\
        );

    \I__4018\ : CEMux
    port map (
            O => \N__18466\,
            I => \N__18460\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__18463\,
            I => \N__18455\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__18460\,
            I => \N__18452\
        );

    \I__4015\ : CEMux
    port map (
            O => \N__18459\,
            I => \N__18449\
        );

    \I__4014\ : CEMux
    port map (
            O => \N__18458\,
            I => \N__18446\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__18455\,
            I => \N__18443\
        );

    \I__4012\ : Sp12to4
    port map (
            O => \N__18452\,
            I => \N__18438\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__18449\,
            I => \N__18438\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18435\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__18443\,
            I => \transmit_module.n2321\
        );

    \I__4008\ : Odrv12
    port map (
            O => \N__18438\,
            I => \transmit_module.n2321\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__18435\,
            I => \transmit_module.n2321\
        );

    \I__4006\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__4004\ : Span4Mux_v
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__4003\ : Span4Mux_v
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__4002\ : Span4Mux_v
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__4001\ : Sp12to4
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__4000\ : Odrv12
    port map (
            O => \N__18410\,
            I => \line_buffer.n625\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__3995\ : Span4Mux_h
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__18392\,
            I => \line_buffer.n633\
        );

    \I__3993\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__3991\ : Span4Mux_v
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__3990\ : Odrv4
    port map (
            O => \N__18380\,
            I => \line_buffer.n3827\
        );

    \I__3989\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__3986\ : Sp12to4
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__3985\ : Span12Mux_h
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__3984\ : Span12Mux_v
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__3983\ : Odrv12
    port map (
            O => \N__18359\,
            I => \line_buffer.n598\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__3981\ : InMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__18341\,
            I => \line_buffer.n606\
        );

    \I__3976\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18335\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__18335\,
            I => \line_buffer.n3767\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__3972\ : Span4Mux_v
    port map (
            O => \N__18326\,
            I => \N__18323\
        );

    \I__3971\ : Sp12to4
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__3970\ : Odrv12
    port map (
            O => \N__18320\,
            I => \line_buffer.n506\
        );

    \I__3969\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18314\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__18314\,
            I => \N__18311\
        );

    \I__3967\ : Span4Mux_v
    port map (
            O => \N__18311\,
            I => \N__18308\
        );

    \I__3966\ : Sp12to4
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__3965\ : Span12Mux_h
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__3964\ : Odrv12
    port map (
            O => \N__18302\,
            I => \line_buffer.n498\
        );

    \I__3963\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18296\,
            I => \N__18293\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__18290\,
            I => \line_buffer.n3714\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18284\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__3957\ : Span12Mux_h
    port map (
            O => \N__18281\,
            I => \N__18278\
        );

    \I__3956\ : Odrv12
    port map (
            O => \N__18278\,
            I => \line_buffer.n510\
        );

    \I__3955\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__18272\,
            I => \N__18269\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__18269\,
            I => \N__18266\
        );

    \I__3952\ : Span4Mux_h
    port map (
            O => \N__18266\,
            I => \N__18263\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__18263\,
            I => \line_buffer.n502\
        );

    \I__3950\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__3948\ : Span4Mux_v
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__18251\,
            I => \line_buffer.n3717\
        );

    \I__3946\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18245\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__18242\,
            I => \line_buffer.n3715\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__18239\,
            I => \line_buffer.n3773_cascade_\
        );

    \I__3942\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__18230\,
            I => \TX_DATA_3\
        );

    \I__3939\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18224\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__18224\,
            I => \N__18221\
        );

    \I__3937\ : Span12Mux_h
    port map (
            O => \N__18221\,
            I => \N__18218\
        );

    \I__3936\ : Odrv12
    port map (
            O => \N__18218\,
            I => \line_buffer.n594\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__18215\,
            I => \N__18212\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__3932\ : Span4Mux_v
    port map (
            O => \N__18206\,
            I => \N__18203\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__3930\ : Span4Mux_h
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__18197\,
            I => \line_buffer.n602\
        );

    \I__3928\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18191\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__3926\ : Span4Mux_h
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__3925\ : Span4Mux_v
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__3924\ : Sp12to4
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__3923\ : Span12Mux_v
    port map (
            O => \N__18179\,
            I => \N__18176\
        );

    \I__3922\ : Odrv12
    port map (
            O => \N__18176\,
            I => \line_buffer.n497\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__18173\,
            I => \line_buffer.n3803_cascade_\
        );

    \I__3920\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__3918\ : Span4Mux_v
    port map (
            O => \N__18164\,
            I => \N__18161\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__3916\ : Sp12to4
    port map (
            O => \N__18158\,
            I => \N__18155\
        );

    \I__3915\ : Odrv12
    port map (
            O => \N__18155\,
            I => \line_buffer.n505\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__18152\,
            I => \line_buffer.n3806_cascade_\
        );

    \I__3913\ : InMux
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__18146\,
            I => \line_buffer.n3782\
        );

    \I__3911\ : InMux
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__18140\,
            I => \N__18137\
        );

    \I__3909\ : Odrv12
    port map (
            O => \N__18137\,
            I => \TX_DATA_2\
        );

    \I__3908\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__3906\ : Odrv12
    port map (
            O => \N__18128\,
            I => \line_buffer.n635\
        );

    \I__3905\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__3903\ : Span12Mux_h
    port map (
            O => \N__18119\,
            I => \N__18116\
        );

    \I__3902\ : Span12Mux_v
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__3901\ : Odrv12
    port map (
            O => \N__18113\,
            I => \line_buffer.n627\
        );

    \I__3900\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__18107\,
            I => \line_buffer.n3706\
        );

    \I__3898\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__3896\ : Span4Mux_v
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__3895\ : Sp12to4
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__3894\ : Span12Mux_h
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__3893\ : Span12Mux_v
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__3892\ : Odrv12
    port map (
            O => \N__18086\,
            I => \line_buffer.n626\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__3890\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__18077\,
            I => \N__18074\
        );

    \I__3888\ : Span4Mux_h
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__3887\ : Span4Mux_h
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__18068\,
            I => \line_buffer.n634\
        );

    \I__3885\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__18062\,
            I => \line_buffer.n3779\
        );

    \I__3883\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__3881\ : Odrv12
    port map (
            O => \N__18053\,
            I => \line_buffer.n3703\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \line_buffer.n3791_cascade_\
        );

    \I__3879\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__3876\ : Odrv4
    port map (
            O => \N__18038\,
            I => \TX_DATA_7\
        );

    \I__3875\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__18032\,
            I => \transmit_module.Y_DELTA_PATTERN_38\
        );

    \I__3873\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18026\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__18026\,
            I => \transmit_module.Y_DELTA_PATTERN_35\
        );

    \I__3871\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18020\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__18020\,
            I => \transmit_module.Y_DELTA_PATTERN_37\
        );

    \I__3869\ : InMux
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__18014\,
            I => \transmit_module.Y_DELTA_PATTERN_36\
        );

    \I__3867\ : InMux
    port map (
            O => \N__18011\,
            I => \N__18008\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__3865\ : Span4Mux_h
    port map (
            O => \N__18005\,
            I => \N__18002\
        );

    \I__3864\ : Span4Mux_h
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__17999\,
            I => \transmit_module.Y_DELTA_PATTERN_40\
        );

    \I__3862\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17993\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__17993\,
            I => \transmit_module.Y_DELTA_PATTERN_39\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17987\,
            I => \transmit_module.Y_DELTA_PATTERN_34\
        );

    \I__3858\ : CEMux
    port map (
            O => \N__17984\,
            I => \N__17977\
        );

    \I__3857\ : CEMux
    port map (
            O => \N__17983\,
            I => \N__17974\
        );

    \I__3856\ : CEMux
    port map (
            O => \N__17982\,
            I => \N__17971\
        );

    \I__3855\ : CEMux
    port map (
            O => \N__17981\,
            I => \N__17966\
        );

    \I__3854\ : CEMux
    port map (
            O => \N__17980\,
            I => \N__17963\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17977\,
            I => \N__17959\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__17974\,
            I => \N__17954\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__17971\,
            I => \N__17954\
        );

    \I__3850\ : CEMux
    port map (
            O => \N__17970\,
            I => \N__17951\
        );

    \I__3849\ : CEMux
    port map (
            O => \N__17969\,
            I => \N__17948\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__17966\,
            I => \N__17943\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__17963\,
            I => \N__17943\
        );

    \I__3846\ : CEMux
    port map (
            O => \N__17962\,
            I => \N__17940\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__17959\,
            I => \N__17936\
        );

    \I__3844\ : Span4Mux_v
    port map (
            O => \N__17954\,
            I => \N__17931\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17951\,
            I => \N__17931\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17948\,
            I => \N__17928\
        );

    \I__3841\ : Span4Mux_v
    port map (
            O => \N__17943\,
            I => \N__17925\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__17940\,
            I => \N__17922\
        );

    \I__3839\ : CEMux
    port map (
            O => \N__17939\,
            I => \N__17919\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__17936\,
            I => \N__17914\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__17931\,
            I => \N__17914\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__17928\,
            I => \N__17910\
        );

    \I__3835\ : Span4Mux_h
    port map (
            O => \N__17925\,
            I => \N__17905\
        );

    \I__3834\ : Span4Mux_v
    port map (
            O => \N__17922\,
            I => \N__17905\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__17919\,
            I => \N__17902\
        );

    \I__3832\ : Span4Mux_h
    port map (
            O => \N__17914\,
            I => \N__17899\
        );

    \I__3831\ : CEMux
    port map (
            O => \N__17913\,
            I => \N__17896\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__17910\,
            I => \transmit_module.n3865\
        );

    \I__3829\ : Odrv4
    port map (
            O => \N__17905\,
            I => \transmit_module.n3865\
        );

    \I__3828\ : Odrv12
    port map (
            O => \N__17902\,
            I => \transmit_module.n3865\
        );

    \I__3827\ : Odrv4
    port map (
            O => \N__17899\,
            I => \transmit_module.n3865\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__17896\,
            I => \transmit_module.n3865\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17882\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__17882\,
            I => \N__17879\
        );

    \I__3823\ : Span12Mux_h
    port map (
            O => \N__17879\,
            I => \N__17876\
        );

    \I__3822\ : Span12Mux_v
    port map (
            O => \N__17876\,
            I => \N__17873\
        );

    \I__3821\ : Odrv12
    port map (
            O => \N__17873\,
            I => \line_buffer.n570\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__17870\,
            I => \N__17867\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__17864\,
            I => \N__17861\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__17861\,
            I => \N__17858\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__17858\,
            I => \N__17855\
        );

    \I__3815\ : Sp12to4
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__3814\ : Odrv12
    port map (
            O => \N__17852\,
            I => \line_buffer.n562\
        );

    \I__3813\ : InMux
    port map (
            O => \N__17849\,
            I => \N__17846\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__3811\ : Odrv12
    port map (
            O => \N__17843\,
            I => \line_buffer.n3705\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__17840\,
            I => \N__17829\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__17839\,
            I => \N__17826\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__17838\,
            I => \N__17823\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__17837\,
            I => \N__17820\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__17836\,
            I => \N__17817\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__17835\,
            I => \N__17814\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__17834\,
            I => \N__17808\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__17833\,
            I => \N__17805\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__17832\,
            I => \N__17802\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17829\,
            I => \N__17792\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17792\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17792\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17792\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17785\
        );

    \I__3796\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17785\
        );

    \I__3795\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17785\
        );

    \I__3794\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17774\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17774\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17774\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17774\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17802\,
            I => \N__17774\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17767\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17792\,
            I => \N__17762\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__17785\,
            I => \N__17762\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__17774\,
            I => \N__17759\
        );

    \I__3785\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17753\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17772\,
            I => \N__17753\
        );

    \I__3783\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17750\
        );

    \I__3782\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17747\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__17767\,
            I => \N__17742\
        );

    \I__3780\ : Span4Mux_h
    port map (
            O => \N__17762\,
            I => \N__17742\
        );

    \I__3779\ : Span4Mux_h
    port map (
            O => \N__17759\,
            I => \N__17739\
        );

    \I__3778\ : InMux
    port map (
            O => \N__17758\,
            I => \N__17736\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17731\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__17750\,
            I => \N__17731\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__17747\,
            I => \N__17728\
        );

    \I__3774\ : Span4Mux_v
    port map (
            O => \N__17742\,
            I => \N__17723\
        );

    \I__3773\ : Span4Mux_v
    port map (
            O => \N__17739\,
            I => \N__17723\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17736\,
            I => \N__17720\
        );

    \I__3771\ : Span4Mux_v
    port map (
            O => \N__17731\,
            I => \N__17715\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__17728\,
            I => \N__17715\
        );

    \I__3769\ : Sp12to4
    port map (
            O => \N__17723\,
            I => \N__17710\
        );

    \I__3768\ : Span12Mux_h
    port map (
            O => \N__17720\,
            I => \N__17710\
        );

    \I__3767\ : Span4Mux_v
    port map (
            O => \N__17715\,
            I => \N__17707\
        );

    \I__3766\ : Odrv12
    port map (
            O => \N__17710\,
            I => \TVP_VSYNC_c\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__17707\,
            I => \TVP_VSYNC_c\
        );

    \I__3764\ : SRMux
    port map (
            O => \N__17702\,
            I => \N__17699\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__17699\,
            I => \N__17694\
        );

    \I__3762\ : SRMux
    port map (
            O => \N__17698\,
            I => \N__17691\
        );

    \I__3761\ : SRMux
    port map (
            O => \N__17697\,
            I => \N__17687\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__17694\,
            I => \N__17682\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__17691\,
            I => \N__17682\
        );

    \I__3758\ : SRMux
    port map (
            O => \N__17690\,
            I => \N__17679\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17676\
        );

    \I__3756\ : Span4Mux_v
    port map (
            O => \N__17682\,
            I => \N__17670\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__17679\,
            I => \N__17670\
        );

    \I__3754\ : Span4Mux_v
    port map (
            O => \N__17676\,
            I => \N__17667\
        );

    \I__3753\ : SRMux
    port map (
            O => \N__17675\,
            I => \N__17664\
        );

    \I__3752\ : Span4Mux_h
    port map (
            O => \N__17670\,
            I => \N__17661\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__17667\,
            I => \N__17656\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__17664\,
            I => \N__17656\
        );

    \I__3749\ : Span4Mux_v
    port map (
            O => \N__17661\,
            I => \N__17653\
        );

    \I__3748\ : Span4Mux_v
    port map (
            O => \N__17656\,
            I => \N__17650\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__17653\,
            I => \receive_module.BRAM_ADDR_13__N_31\
        );

    \I__3746\ : Odrv4
    port map (
            O => \N__17650\,
            I => \receive_module.BRAM_ADDR_13__N_31\
        );

    \I__3745\ : SRMux
    port map (
            O => \N__17645\,
            I => \N__17640\
        );

    \I__3744\ : SRMux
    port map (
            O => \N__17644\,
            I => \N__17635\
        );

    \I__3743\ : CEMux
    port map (
            O => \N__17643\,
            I => \N__17632\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__17640\,
            I => \N__17629\
        );

    \I__3741\ : InMux
    port map (
            O => \N__17639\,
            I => \N__17626\
        );

    \I__3740\ : CEMux
    port map (
            O => \N__17638\,
            I => \N__17623\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17635\,
            I => \N__17620\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__17632\,
            I => \N__17617\
        );

    \I__3737\ : Span4Mux_v
    port map (
            O => \N__17629\,
            I => \N__17612\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__17626\,
            I => \N__17612\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__17623\,
            I => \N__17609\
        );

    \I__3734\ : Sp12to4
    port map (
            O => \N__17620\,
            I => \N__17606\
        );

    \I__3733\ : Span4Mux_h
    port map (
            O => \N__17617\,
            I => \N__17601\
        );

    \I__3732\ : Span4Mux_h
    port map (
            O => \N__17612\,
            I => \N__17601\
        );

    \I__3731\ : Odrv12
    port map (
            O => \N__17609\,
            I => \transmit_module.video_signal_controller.n2030\
        );

    \I__3730\ : Odrv12
    port map (
            O => \N__17606\,
            I => \transmit_module.video_signal_controller.n2030\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__17601\,
            I => \transmit_module.video_signal_controller.n2030\
        );

    \I__3728\ : SRMux
    port map (
            O => \N__17594\,
            I => \N__17590\
        );

    \I__3727\ : SRMux
    port map (
            O => \N__17593\,
            I => \N__17587\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17590\,
            I => \N__17584\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__17587\,
            I => \N__17581\
        );

    \I__3724\ : Span4Mux_h
    port map (
            O => \N__17584\,
            I => \N__17578\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__17581\,
            I => \transmit_module.video_signal_controller.n2551\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__17578\,
            I => \transmit_module.video_signal_controller.n2551\
        );

    \I__3721\ : IoInMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3719\ : Span4Mux_s2_h
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__3718\ : Span4Mux_h
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__3717\ : Span4Mux_h
    port map (
            O => \N__17561\,
            I => \N__17557\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17560\,
            I => \N__17554\
        );

    \I__3715\ : Span4Mux_v
    port map (
            O => \N__17557\,
            I => \N__17551\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__17554\,
            I => \N__17548\
        );

    \I__3713\ : Span4Mux_v
    port map (
            O => \N__17551\,
            I => \N__17543\
        );

    \I__3712\ : Span4Mux_v
    port map (
            O => \N__17548\,
            I => \N__17543\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__17543\,
            I => \DEBUG_c_6\
        );

    \I__3710\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__17537\,
            I => \transmit_module.video_signal_controller.SYNC_BUFF1\
        );

    \I__3708\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17531\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__17531\,
            I => \transmit_module.video_signal_controller.SYNC_BUFF2\
        );

    \I__3706\ : IoInMux
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__17525\,
            I => \N__17522\
        );

    \I__3704\ : IoSpan4Mux
    port map (
            O => \N__17522\,
            I => \N__17519\
        );

    \I__3703\ : Span4Mux_s3_h
    port map (
            O => \N__17519\,
            I => \N__17515\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17512\
        );

    \I__3701\ : Span4Mux_h
    port map (
            O => \N__17515\,
            I => \N__17509\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17512\,
            I => \N__17506\
        );

    \I__3699\ : Span4Mux_h
    port map (
            O => \N__17509\,
            I => \N__17501\
        );

    \I__3698\ : Span4Mux_v
    port map (
            O => \N__17506\,
            I => \N__17501\
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__17501\,
            I => n3852
        );

    \I__3696\ : CEMux
    port map (
            O => \N__17498\,
            I => \N__17494\
        );

    \I__3695\ : CEMux
    port map (
            O => \N__17497\,
            I => \N__17491\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__17494\,
            I => \N__17487\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__17491\,
            I => \N__17484\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17481\
        );

    \I__3691\ : Span4Mux_h
    port map (
            O => \N__17487\,
            I => \N__17478\
        );

    \I__3690\ : Span4Mux_h
    port map (
            O => \N__17484\,
            I => \N__17475\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__17481\,
            I => \N__17472\
        );

    \I__3688\ : Span4Mux_h
    port map (
            O => \N__17478\,
            I => \N__17469\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__17475\,
            I => \N__17464\
        );

    \I__3686\ : Span4Mux_h
    port map (
            O => \N__17472\,
            I => \N__17464\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__17469\,
            I => \transmit_module.n2039\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__17464\,
            I => \transmit_module.n2039\
        );

    \I__3683\ : InMux
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__17456\,
            I => \N__17453\
        );

    \I__3681\ : Span4Mux_v
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__3680\ : Span4Mux_h
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__3679\ : Span4Mux_h
    port map (
            O => \N__17447\,
            I => \N__17444\
        );

    \I__3678\ : Odrv4
    port map (
            O => \N__17444\,
            I => \line_buffer.n603\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17438\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__3675\ : Span4Mux_v
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3674\ : Sp12to4
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__3673\ : Odrv12
    port map (
            O => \N__17429\,
            I => \line_buffer.n595\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17426\,
            I => \N__17423\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__17420\,
            I => \N__17417\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__3668\ : Span4Mux_h
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__3667\ : Span4Mux_v
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__17408\,
            I => \line_buffer.n569\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__3664\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3661\ : Span4Mux_h
    port map (
            O => \N__17393\,
            I => \N__17390\
        );

    \I__3660\ : Span4Mux_h
    port map (
            O => \N__17390\,
            I => \N__17387\
        );

    \I__3659\ : Odrv4
    port map (
            O => \N__17387\,
            I => \line_buffer.n561\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__17384\,
            I => \line_buffer.n3830_cascade_\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17381\,
            I => \N__17378\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__17378\,
            I => \N__17375\
        );

    \I__3655\ : Span4Mux_h
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__17372\,
            I => \TX_DATA_1\
        );

    \I__3653\ : InMux
    port map (
            O => \N__17369\,
            I => \N__17365\
        );

    \I__3652\ : InMux
    port map (
            O => \N__17368\,
            I => \N__17361\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__17365\,
            I => \N__17358\
        );

    \I__3650\ : InMux
    port map (
            O => \N__17364\,
            I => \N__17355\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__17361\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__17358\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__17355\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__3646\ : InMux
    port map (
            O => \N__17348\,
            I => \N__17343\
        );

    \I__3645\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17340\
        );

    \I__3644\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17337\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__17343\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__17340\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__17337\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__3640\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17327\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__17324\,
            I => \transmit_module.video_signal_controller.n3858\
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__17321\,
            I => \transmit_module.n213_cascade_\
        );

    \I__3636\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17312\
        );

    \I__3635\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17307\
        );

    \I__3634\ : InMux
    port map (
            O => \N__17316\,
            I => \N__17307\
        );

    \I__3633\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17304\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__17312\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__17307\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__17304\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17297\,
            I => \N__17294\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__17294\,
            I => \transmit_module.n184\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17291\,
            I => \N__17287\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17290\,
            I => \N__17284\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__17287\,
            I => \transmit_module.n216\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__17284\,
            I => \transmit_module.n216\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__17279\,
            I => \N__17275\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__17278\,
            I => \N__17272\
        );

    \I__3621\ : CascadeBuf
    port map (
            O => \N__17275\,
            I => \N__17269\
        );

    \I__3620\ : CascadeBuf
    port map (
            O => \N__17272\,
            I => \N__17266\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__17269\,
            I => \N__17263\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__17266\,
            I => \N__17260\
        );

    \I__3617\ : CascadeBuf
    port map (
            O => \N__17263\,
            I => \N__17257\
        );

    \I__3616\ : CascadeBuf
    port map (
            O => \N__17260\,
            I => \N__17254\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__17257\,
            I => \N__17251\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__17254\,
            I => \N__17248\
        );

    \I__3613\ : CascadeBuf
    port map (
            O => \N__17251\,
            I => \N__17245\
        );

    \I__3612\ : CascadeBuf
    port map (
            O => \N__17248\,
            I => \N__17242\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__17245\,
            I => \N__17239\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__17242\,
            I => \N__17236\
        );

    \I__3609\ : CascadeBuf
    port map (
            O => \N__17239\,
            I => \N__17233\
        );

    \I__3608\ : CascadeBuf
    port map (
            O => \N__17236\,
            I => \N__17230\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__17233\,
            I => \N__17227\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__17230\,
            I => \N__17224\
        );

    \I__3605\ : CascadeBuf
    port map (
            O => \N__17227\,
            I => \N__17221\
        );

    \I__3604\ : CascadeBuf
    port map (
            O => \N__17224\,
            I => \N__17218\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__17221\,
            I => \N__17215\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__17218\,
            I => \N__17212\
        );

    \I__3601\ : CascadeBuf
    port map (
            O => \N__17215\,
            I => \N__17209\
        );

    \I__3600\ : CascadeBuf
    port map (
            O => \N__17212\,
            I => \N__17206\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__17209\,
            I => \N__17203\
        );

    \I__3598\ : CascadeMux
    port map (
            O => \N__17206\,
            I => \N__17200\
        );

    \I__3597\ : CascadeBuf
    port map (
            O => \N__17203\,
            I => \N__17197\
        );

    \I__3596\ : CascadeBuf
    port map (
            O => \N__17200\,
            I => \N__17194\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__17197\,
            I => \N__17191\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__17194\,
            I => \N__17188\
        );

    \I__3593\ : CascadeBuf
    port map (
            O => \N__17191\,
            I => \N__17185\
        );

    \I__3592\ : CascadeBuf
    port map (
            O => \N__17188\,
            I => \N__17182\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__17185\,
            I => \N__17179\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__17182\,
            I => \N__17176\
        );

    \I__3589\ : CascadeBuf
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__3588\ : CascadeBuf
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__17173\,
            I => \N__17167\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__17170\,
            I => \N__17164\
        );

    \I__3585\ : CascadeBuf
    port map (
            O => \N__17167\,
            I => \N__17161\
        );

    \I__3584\ : CascadeBuf
    port map (
            O => \N__17164\,
            I => \N__17158\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__17161\,
            I => \N__17155\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__17158\,
            I => \N__17152\
        );

    \I__3581\ : CascadeBuf
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__3580\ : CascadeBuf
    port map (
            O => \N__17152\,
            I => \N__17146\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__17149\,
            I => \N__17143\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__17146\,
            I => \N__17140\
        );

    \I__3577\ : CascadeBuf
    port map (
            O => \N__17143\,
            I => \N__17137\
        );

    \I__3576\ : CascadeBuf
    port map (
            O => \N__17140\,
            I => \N__17134\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__17134\,
            I => \N__17128\
        );

    \I__3573\ : CascadeBuf
    port map (
            O => \N__17131\,
            I => \N__17125\
        );

    \I__3572\ : CascadeBuf
    port map (
            O => \N__17128\,
            I => \N__17122\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__17125\,
            I => \N__17119\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__17122\,
            I => \N__17116\
        );

    \I__3569\ : CascadeBuf
    port map (
            O => \N__17119\,
            I => \N__17113\
        );

    \I__3568\ : CascadeBuf
    port map (
            O => \N__17116\,
            I => \N__17110\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__17113\,
            I => \N__17107\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__17110\,
            I => \N__17104\
        );

    \I__3565\ : CascadeBuf
    port map (
            O => \N__17107\,
            I => \N__17101\
        );

    \I__3564\ : CascadeBuf
    port map (
            O => \N__17104\,
            I => \N__17098\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__17101\,
            I => \N__17095\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__17098\,
            I => \N__17092\
        );

    \I__3561\ : InMux
    port map (
            O => \N__17095\,
            I => \N__17089\
        );

    \I__3560\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17086\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__17089\,
            I => \N__17083\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__17086\,
            I => \N__17080\
        );

    \I__3557\ : Span12Mux_s10_h
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__3556\ : Span12Mux_s9_h
    port map (
            O => \N__17080\,
            I => \N__17074\
        );

    \I__3555\ : Span12Mux_v
    port map (
            O => \N__17077\,
            I => \N__17069\
        );

    \I__3554\ : Span12Mux_v
    port map (
            O => \N__17074\,
            I => \N__17069\
        );

    \I__3553\ : Odrv12
    port map (
            O => \N__17069\,
            I => n24
        );

    \I__3552\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17063\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__17063\,
            I => \transmit_module.ADDR_Y_COMPONENT_9\
        );

    \I__3550\ : InMux
    port map (
            O => \N__17060\,
            I => \N__17056\
        );

    \I__3549\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17053\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__17056\,
            I => \transmit_module.n181\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__17053\,
            I => \transmit_module.n181\
        );

    \I__3546\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__17045\,
            I => \transmit_module.n213\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__17042\,
            I => \N__17038\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__17041\,
            I => \N__17035\
        );

    \I__3542\ : CascadeBuf
    port map (
            O => \N__17038\,
            I => \N__17032\
        );

    \I__3541\ : CascadeBuf
    port map (
            O => \N__17035\,
            I => \N__17029\
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__17032\,
            I => \N__17026\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__17029\,
            I => \N__17023\
        );

    \I__3538\ : CascadeBuf
    port map (
            O => \N__17026\,
            I => \N__17020\
        );

    \I__3537\ : CascadeBuf
    port map (
            O => \N__17023\,
            I => \N__17017\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__17020\,
            I => \N__17014\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__17017\,
            I => \N__17011\
        );

    \I__3534\ : CascadeBuf
    port map (
            O => \N__17014\,
            I => \N__17008\
        );

    \I__3533\ : CascadeBuf
    port map (
            O => \N__17011\,
            I => \N__17005\
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__17008\,
            I => \N__17002\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__17005\,
            I => \N__16999\
        );

    \I__3530\ : CascadeBuf
    port map (
            O => \N__17002\,
            I => \N__16996\
        );

    \I__3529\ : CascadeBuf
    port map (
            O => \N__16999\,
            I => \N__16993\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__16996\,
            I => \N__16990\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__16993\,
            I => \N__16987\
        );

    \I__3526\ : CascadeBuf
    port map (
            O => \N__16990\,
            I => \N__16984\
        );

    \I__3525\ : CascadeBuf
    port map (
            O => \N__16987\,
            I => \N__16981\
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__16984\,
            I => \N__16978\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__16981\,
            I => \N__16975\
        );

    \I__3522\ : CascadeBuf
    port map (
            O => \N__16978\,
            I => \N__16972\
        );

    \I__3521\ : CascadeBuf
    port map (
            O => \N__16975\,
            I => \N__16969\
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__16972\,
            I => \N__16966\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__16969\,
            I => \N__16963\
        );

    \I__3518\ : CascadeBuf
    port map (
            O => \N__16966\,
            I => \N__16960\
        );

    \I__3517\ : CascadeBuf
    port map (
            O => \N__16963\,
            I => \N__16957\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__16960\,
            I => \N__16954\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__16957\,
            I => \N__16951\
        );

    \I__3514\ : CascadeBuf
    port map (
            O => \N__16954\,
            I => \N__16948\
        );

    \I__3513\ : CascadeBuf
    port map (
            O => \N__16951\,
            I => \N__16945\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__16948\,
            I => \N__16942\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__16945\,
            I => \N__16939\
        );

    \I__3510\ : CascadeBuf
    port map (
            O => \N__16942\,
            I => \N__16936\
        );

    \I__3509\ : CascadeBuf
    port map (
            O => \N__16939\,
            I => \N__16933\
        );

    \I__3508\ : CascadeMux
    port map (
            O => \N__16936\,
            I => \N__16930\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__16933\,
            I => \N__16927\
        );

    \I__3506\ : CascadeBuf
    port map (
            O => \N__16930\,
            I => \N__16924\
        );

    \I__3505\ : CascadeBuf
    port map (
            O => \N__16927\,
            I => \N__16921\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__16924\,
            I => \N__16918\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__16921\,
            I => \N__16915\
        );

    \I__3502\ : CascadeBuf
    port map (
            O => \N__16918\,
            I => \N__16912\
        );

    \I__3501\ : CascadeBuf
    port map (
            O => \N__16915\,
            I => \N__16909\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__16912\,
            I => \N__16906\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__16909\,
            I => \N__16903\
        );

    \I__3498\ : CascadeBuf
    port map (
            O => \N__16906\,
            I => \N__16900\
        );

    \I__3497\ : CascadeBuf
    port map (
            O => \N__16903\,
            I => \N__16897\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__16900\,
            I => \N__16894\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__16897\,
            I => \N__16891\
        );

    \I__3494\ : CascadeBuf
    port map (
            O => \N__16894\,
            I => \N__16888\
        );

    \I__3493\ : CascadeBuf
    port map (
            O => \N__16891\,
            I => \N__16885\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__16888\,
            I => \N__16882\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__16885\,
            I => \N__16879\
        );

    \I__3490\ : CascadeBuf
    port map (
            O => \N__16882\,
            I => \N__16876\
        );

    \I__3489\ : CascadeBuf
    port map (
            O => \N__16879\,
            I => \N__16873\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__16876\,
            I => \N__16870\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__16873\,
            I => \N__16867\
        );

    \I__3486\ : CascadeBuf
    port map (
            O => \N__16870\,
            I => \N__16864\
        );

    \I__3485\ : CascadeBuf
    port map (
            O => \N__16867\,
            I => \N__16861\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__16864\,
            I => \N__16858\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__16861\,
            I => \N__16855\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16858\,
            I => \N__16852\
        );

    \I__3481\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16849\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16852\,
            I => \N__16846\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__16849\,
            I => \N__16843\
        );

    \I__3478\ : Span12Mux_h
    port map (
            O => \N__16846\,
            I => \N__16838\
        );

    \I__3477\ : Span12Mux_h
    port map (
            O => \N__16843\,
            I => \N__16838\
        );

    \I__3476\ : Span12Mux_v
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__3475\ : Odrv12
    port map (
            O => \N__16835\,
            I => n21
        );

    \I__3474\ : InMux
    port map (
            O => \N__16832\,
            I => \N__16829\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__16829\,
            I => \N__16826\
        );

    \I__3472\ : Span4Mux_h
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__3471\ : Span4Mux_v
    port map (
            O => \N__16823\,
            I => \N__16820\
        );

    \I__3470\ : Span4Mux_h
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__3469\ : Span4Mux_h
    port map (
            O => \N__16817\,
            I => \N__16814\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__16814\,
            I => \line_buffer.n509\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__16811\,
            I => \N__16808\
        );

    \I__3466\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__16805\,
            I => \N__16802\
        );

    \I__3464\ : Span4Mux_v
    port map (
            O => \N__16802\,
            I => \N__16799\
        );

    \I__3463\ : Span4Mux_v
    port map (
            O => \N__16799\,
            I => \N__16796\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__16796\,
            I => \N__16793\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__16793\,
            I => \line_buffer.n501\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16787\,
            I => \line_buffer.n3770\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__16778\,
            I => \N__16775\
        );

    \I__3455\ : Span4Mux_h
    port map (
            O => \N__16775\,
            I => \N__16772\
        );

    \I__3454\ : Span4Mux_h
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__16769\,
            I => \line_buffer.n571\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__3450\ : Span12Mux_h
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__3449\ : Odrv12
    port map (
            O => \N__16757\,
            I => \line_buffer.n563\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__16751\,
            I => \receive_module.rx_counter.n11\
        );

    \I__3446\ : IoInMux
    port map (
            O => \N__16748\,
            I => \N__16745\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__3444\ : Span4Mux_s1_v
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__3443\ : Span4Mux_v
    port map (
            O => \N__16739\,
            I => \N__16736\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__16736\,
            I => \N__16733\
        );

    \I__3441\ : Span4Mux_h
    port map (
            O => \N__16733\,
            I => \N__16729\
        );

    \I__3440\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16726\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__16729\,
            I => \LED_c\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__16726\,
            I => \LED_c\
        );

    \I__3437\ : CEMux
    port map (
            O => \N__16721\,
            I => \N__16717\
        );

    \I__3436\ : CEMux
    port map (
            O => \N__16720\,
            I => \N__16714\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__16717\,
            I => \receive_module.rx_counter.n3862\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__16714\,
            I => \receive_module.rx_counter.n3862\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16709\,
            I => \N__16706\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16706\,
            I => \N__16703\
        );

    \I__3431\ : Span4Mux_h
    port map (
            O => \N__16703\,
            I => \N__16697\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16692\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16692\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16689\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__16697\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__16692\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__16689\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__16679\,
            I => \N__16676\
        );

    \I__3422\ : Span4Mux_h
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__16673\,
            I => \transmit_module.ADDR_Y_COMPONENT_6\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16664\
        );

    \I__3419\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16659\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16659\
        );

    \I__3417\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16656\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__16664\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16659\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__16656\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__3413\ : InMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16646\,
            I => \transmit_module.ADDR_Y_COMPONENT_2\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__16640\,
            I => \transmit_module.ADDR_Y_COMPONENT_7\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__16634\,
            I => \transmit_module.ADDR_Y_COMPONENT_4\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__16631\,
            I => \transmit_module.n184_cascade_\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16625\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__16625\,
            I => \transmit_module.n200\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16616\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16621\,
            I => \N__16611\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16620\,
            I => \N__16611\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16608\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__16616\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16611\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16608\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__16598\,
            I => \transmit_module.n197\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__16589\,
            I => \N__16585\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16582\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__16585\,
            I => \transmit_module.n188\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__16582\,
            I => \transmit_module.n188\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16572\
        );

    \I__3388\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16569\
        );

    \I__3387\ : InMux
    port map (
            O => \N__16575\,
            I => \N__16565\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__16572\,
            I => \N__16560\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16560\
        );

    \I__3384\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16557\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__16565\,
            I => \N__16554\
        );

    \I__3382\ : Span4Mux_v
    port map (
            O => \N__16560\,
            I => \N__16551\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__16557\,
            I => \transmit_module.n3859\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__16554\,
            I => \transmit_module.n3859\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__16551\,
            I => \transmit_module.n3859\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16540\
        );

    \I__3377\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16535\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16540\,
            I => \N__16532\
        );

    \I__3375\ : InMux
    port map (
            O => \N__16539\,
            I => \N__16529\
        );

    \I__3374\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16526\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__16535\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__16532\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__16529\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__16526\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3369\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__16514\,
            I => \transmit_module.ADDR_Y_COMPONENT_1\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__16511\,
            I => \N__16508\
        );

    \I__3366\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3364\ : Span4Mux_h
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__16499\,
            I => \transmit_module.ADDR_Y_COMPONENT_11\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__16496\,
            I => \N__16493\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16493\,
            I => \N__16490\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__3359\ : Span4Mux_h
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__3358\ : Odrv4
    port map (
            O => \N__16484\,
            I => \transmit_module.ADDR_Y_COMPONENT_12\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16478\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__3355\ : Odrv12
    port map (
            O => \N__16475\,
            I => \transmit_module.ADDR_Y_COMPONENT_13\
        );

    \I__3354\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16467\
        );

    \I__3353\ : InMux
    port map (
            O => \N__16471\,
            I => \N__16464\
        );

    \I__3352\ : InMux
    port map (
            O => \N__16470\,
            I => \N__16460\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__16467\,
            I => \N__16455\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__16464\,
            I => \N__16455\
        );

    \I__3349\ : InMux
    port map (
            O => \N__16463\,
            I => \N__16452\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__16460\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__16455\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__16452\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3345\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16442\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__16442\,
            I => \transmit_module.ADDR_Y_COMPONENT_0\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__16436\,
            I => \N__16432\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16428\
        );

    \I__3340\ : Span4Mux_h
    port map (
            O => \N__16432\,
            I => \N__16424\
        );

    \I__3339\ : InMux
    port map (
            O => \N__16431\,
            I => \N__16421\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__16428\,
            I => \N__16418\
        );

    \I__3337\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16415\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__16424\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__16421\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__16418\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__16415\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__3332\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__16403\,
            I => \N__16400\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__16400\,
            I => \transmit_module.ADDR_Y_COMPONENT_5\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__3328\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16390\
        );

    \I__3327\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16385\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__16390\,
            I => \N__16382\
        );

    \I__3325\ : InMux
    port map (
            O => \N__16389\,
            I => \N__16377\
        );

    \I__3324\ : InMux
    port map (
            O => \N__16388\,
            I => \N__16377\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__16385\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__16382\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__16377\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16370\,
            I => \transmit_module.video_signal_controller.n3369\
        );

    \I__3319\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16362\
        );

    \I__3318\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16359\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16356\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__16362\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__16359\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__16356\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__3313\ : InMux
    port map (
            O => \N__16349\,
            I => \transmit_module.video_signal_controller.n3370\
        );

    \I__3312\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16341\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16338\
        );

    \I__3310\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16335\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__16341\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__16338\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__16335\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__3306\ : InMux
    port map (
            O => \N__16328\,
            I => \transmit_module.video_signal_controller.n3371\
        );

    \I__3305\ : InMux
    port map (
            O => \N__16325\,
            I => \N__16321\
        );

    \I__3304\ : InMux
    port map (
            O => \N__16324\,
            I => \N__16318\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__16321\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__16318\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__3301\ : InMux
    port map (
            O => \N__16313\,
            I => \transmit_module.video_signal_controller.n3372\
        );

    \I__3300\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16306\
        );

    \I__3299\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16303\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__16306\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__16303\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16298\,
            I => \bfn_14_14_0_\
        );

    \I__3295\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16290\
        );

    \I__3294\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16285\
        );

    \I__3293\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16285\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__16290\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__16285\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__3290\ : InMux
    port map (
            O => \N__16280\,
            I => \transmit_module.video_signal_controller.n3374\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16277\,
            I => \transmit_module.video_signal_controller.n3375\
        );

    \I__3288\ : InMux
    port map (
            O => \N__16274\,
            I => \transmit_module.video_signal_controller.n3376\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__16271\,
            I => \N__16268\
        );

    \I__3286\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16265\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__16265\,
            I => \N__16262\
        );

    \I__3284\ : Span4Mux_v
    port map (
            O => \N__16262\,
            I => \N__16255\
        );

    \I__3283\ : InMux
    port map (
            O => \N__16261\,
            I => \N__16250\
        );

    \I__3282\ : InMux
    port map (
            O => \N__16260\,
            I => \N__16250\
        );

    \I__3281\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16247\
        );

    \I__3280\ : InMux
    port map (
            O => \N__16258\,
            I => \N__16244\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__16255\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__16250\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__16247\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__16244\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3275\ : IoInMux
    port map (
            O => \N__16235\,
            I => \N__16232\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__16232\,
            I => \N__16229\
        );

    \I__3273\ : Span4Mux_s0_h
    port map (
            O => \N__16229\,
            I => \N__16225\
        );

    \I__3272\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16222\
        );

    \I__3271\ : Sp12to4
    port map (
            O => \N__16225\,
            I => \N__16217\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__16222\,
            I => \N__16214\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__16221\,
            I => \N__16210\
        );

    \I__3268\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16205\
        );

    \I__3267\ : Span12Mux_v
    port map (
            O => \N__16217\,
            I => \N__16202\
        );

    \I__3266\ : Span4Mux_h
    port map (
            O => \N__16214\,
            I => \N__16199\
        );

    \I__3265\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16194\
        );

    \I__3264\ : InMux
    port map (
            O => \N__16210\,
            I => \N__16194\
        );

    \I__3263\ : InMux
    port map (
            O => \N__16209\,
            I => \N__16189\
        );

    \I__3262\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16189\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__16205\,
            I => \N__16186\
        );

    \I__3260\ : Odrv12
    port map (
            O => \N__16202\,
            I => \ADV_HSYNC_c\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__16199\,
            I => \ADV_HSYNC_c\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__16194\,
            I => \ADV_HSYNC_c\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__16189\,
            I => \ADV_HSYNC_c\
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__16186\,
            I => \ADV_HSYNC_c\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__16175\,
            I => \N__16171\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__16174\,
            I => \N__16168\
        );

    \I__3253\ : CascadeBuf
    port map (
            O => \N__16171\,
            I => \N__16165\
        );

    \I__3252\ : CascadeBuf
    port map (
            O => \N__16168\,
            I => \N__16162\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__16165\,
            I => \N__16159\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__16162\,
            I => \N__16156\
        );

    \I__3249\ : CascadeBuf
    port map (
            O => \N__16159\,
            I => \N__16153\
        );

    \I__3248\ : CascadeBuf
    port map (
            O => \N__16156\,
            I => \N__16150\
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__16153\,
            I => \N__16147\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__16150\,
            I => \N__16144\
        );

    \I__3245\ : CascadeBuf
    port map (
            O => \N__16147\,
            I => \N__16141\
        );

    \I__3244\ : CascadeBuf
    port map (
            O => \N__16144\,
            I => \N__16138\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__16141\,
            I => \N__16135\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__16138\,
            I => \N__16132\
        );

    \I__3241\ : CascadeBuf
    port map (
            O => \N__16135\,
            I => \N__16129\
        );

    \I__3240\ : CascadeBuf
    port map (
            O => \N__16132\,
            I => \N__16126\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__16129\,
            I => \N__16123\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__16126\,
            I => \N__16120\
        );

    \I__3237\ : CascadeBuf
    port map (
            O => \N__16123\,
            I => \N__16117\
        );

    \I__3236\ : CascadeBuf
    port map (
            O => \N__16120\,
            I => \N__16114\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__16117\,
            I => \N__16111\
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__16114\,
            I => \N__16108\
        );

    \I__3233\ : CascadeBuf
    port map (
            O => \N__16111\,
            I => \N__16105\
        );

    \I__3232\ : CascadeBuf
    port map (
            O => \N__16108\,
            I => \N__16102\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__16105\,
            I => \N__16099\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__16102\,
            I => \N__16096\
        );

    \I__3229\ : CascadeBuf
    port map (
            O => \N__16099\,
            I => \N__16093\
        );

    \I__3228\ : CascadeBuf
    port map (
            O => \N__16096\,
            I => \N__16090\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__16093\,
            I => \N__16087\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__16090\,
            I => \N__16084\
        );

    \I__3225\ : CascadeBuf
    port map (
            O => \N__16087\,
            I => \N__16081\
        );

    \I__3224\ : CascadeBuf
    port map (
            O => \N__16084\,
            I => \N__16078\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__16081\,
            I => \N__16075\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__16078\,
            I => \N__16072\
        );

    \I__3221\ : CascadeBuf
    port map (
            O => \N__16075\,
            I => \N__16069\
        );

    \I__3220\ : CascadeBuf
    port map (
            O => \N__16072\,
            I => \N__16066\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__16069\,
            I => \N__16063\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__16066\,
            I => \N__16060\
        );

    \I__3217\ : CascadeBuf
    port map (
            O => \N__16063\,
            I => \N__16057\
        );

    \I__3216\ : CascadeBuf
    port map (
            O => \N__16060\,
            I => \N__16054\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__16057\,
            I => \N__16051\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__16054\,
            I => \N__16048\
        );

    \I__3213\ : CascadeBuf
    port map (
            O => \N__16051\,
            I => \N__16045\
        );

    \I__3212\ : CascadeBuf
    port map (
            O => \N__16048\,
            I => \N__16042\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__16045\,
            I => \N__16039\
        );

    \I__3210\ : CascadeMux
    port map (
            O => \N__16042\,
            I => \N__16036\
        );

    \I__3209\ : CascadeBuf
    port map (
            O => \N__16039\,
            I => \N__16033\
        );

    \I__3208\ : CascadeBuf
    port map (
            O => \N__16036\,
            I => \N__16030\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__16033\,
            I => \N__16027\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__16030\,
            I => \N__16024\
        );

    \I__3205\ : CascadeBuf
    port map (
            O => \N__16027\,
            I => \N__16021\
        );

    \I__3204\ : CascadeBuf
    port map (
            O => \N__16024\,
            I => \N__16018\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__16021\,
            I => \N__16015\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__16018\,
            I => \N__16012\
        );

    \I__3201\ : CascadeBuf
    port map (
            O => \N__16015\,
            I => \N__16009\
        );

    \I__3200\ : CascadeBuf
    port map (
            O => \N__16012\,
            I => \N__16006\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__16009\,
            I => \N__16003\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__16006\,
            I => \N__16000\
        );

    \I__3197\ : CascadeBuf
    port map (
            O => \N__16003\,
            I => \N__15997\
        );

    \I__3196\ : CascadeBuf
    port map (
            O => \N__16000\,
            I => \N__15994\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__15997\,
            I => \N__15991\
        );

    \I__3194\ : CascadeMux
    port map (
            O => \N__15994\,
            I => \N__15988\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15985\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15982\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__15985\,
            I => \N__15979\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__15982\,
            I => \N__15976\
        );

    \I__3189\ : Span4Mux_h
    port map (
            O => \N__15979\,
            I => \N__15972\
        );

    \I__3188\ : Span4Mux_h
    port map (
            O => \N__15976\,
            I => \N__15969\
        );

    \I__3187\ : InMux
    port map (
            O => \N__15975\,
            I => \N__15966\
        );

    \I__3186\ : Sp12to4
    port map (
            O => \N__15972\,
            I => \N__15963\
        );

    \I__3185\ : Sp12to4
    port map (
            O => \N__15969\,
            I => \N__15960\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__15966\,
            I => \N__15957\
        );

    \I__3183\ : Span12Mux_s9_v
    port map (
            O => \N__15963\,
            I => \N__15953\
        );

    \I__3182\ : Span12Mux_s9_v
    port map (
            O => \N__15960\,
            I => \N__15950\
        );

    \I__3181\ : Span4Mux_v
    port map (
            O => \N__15957\,
            I => \N__15947\
        );

    \I__3180\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15944\
        );

    \I__3179\ : Span12Mux_v
    port map (
            O => \N__15953\,
            I => \N__15939\
        );

    \I__3178\ : Span12Mux_v
    port map (
            O => \N__15950\,
            I => \N__15939\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__15947\,
            I => \RX_ADDR_10\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__15944\,
            I => \RX_ADDR_10\
        );

    \I__3175\ : Odrv12
    port map (
            O => \N__15939\,
            I => \RX_ADDR_10\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15929\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__15929\,
            I => \N__15926\
        );

    \I__3172\ : Span4Mux_h
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__15923\,
            I => \receive_module.n126\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15920\,
            I => \receive_module.n3332\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15900\
        );

    \I__3168\ : InMux
    port map (
            O => \N__15916\,
            I => \N__15900\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15915\,
            I => \N__15900\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15914\,
            I => \N__15900\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15913\,
            I => \N__15895\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15912\,
            I => \N__15895\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15911\,
            I => \N__15892\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15889\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15909\,
            I => \N__15886\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__15900\,
            I => \N__15879\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__15895\,
            I => \N__15879\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__15892\,
            I => \N__15879\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__15889\,
            I => \N__15876\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__15886\,
            I => \N__15871\
        );

    \I__3155\ : Span4Mux_v
    port map (
            O => \N__15879\,
            I => \N__15871\
        );

    \I__3154\ : Span4Mux_h
    port map (
            O => \N__15876\,
            I => \N__15868\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__15871\,
            I => \RX_ADDR_11\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__15868\,
            I => \RX_ADDR_11\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15863\,
            I => \receive_module.n3333\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__15860\,
            I => \N__15856\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15848\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15848\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__15855\,
            I => \N__15844\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__15854\,
            I => \N__15841\
        );

    \I__3145\ : InMux
    port map (
            O => \N__15853\,
            I => \N__15836\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__15848\,
            I => \N__15833\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15830\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15820\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15820\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15820\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15820\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15836\,
            I => \N__15817\
        );

    \I__3137\ : Span4Mux_v
    port map (
            O => \N__15833\,
            I => \N__15814\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__15830\,
            I => \N__15811\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15829\,
            I => \N__15808\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__15820\,
            I => \N__15805\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__15817\,
            I => \N__15802\
        );

    \I__3132\ : Span4Mux_h
    port map (
            O => \N__15814\,
            I => \N__15797\
        );

    \I__3131\ : Span4Mux_v
    port map (
            O => \N__15811\,
            I => \N__15797\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__15808\,
            I => \RX_ADDR_12\
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__15805\,
            I => \RX_ADDR_12\
        );

    \I__3128\ : Odrv4
    port map (
            O => \N__15802\,
            I => \RX_ADDR_12\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__15797\,
            I => \RX_ADDR_12\
        );

    \I__3126\ : InMux
    port map (
            O => \N__15788\,
            I => \receive_module.n3334\
        );

    \I__3125\ : CEMux
    port map (
            O => \N__15785\,
            I => \N__15782\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__15776\,
            I => \receive_module.n3854\
        );

    \I__3121\ : IoInMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__15770\,
            I => \N__15767\
        );

    \I__3119\ : Span4Mux_s2_h
    port map (
            O => \N__15767\,
            I => \N__15761\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15766\,
            I => \N__15756\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__15765\,
            I => \N__15753\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__15764\,
            I => \N__15748\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__15761\,
            I => \N__15743\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__15760\,
            I => \N__15740\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__15759\,
            I => \N__15736\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__15756\,
            I => \N__15733\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15753\,
            I => \N__15728\
        );

    \I__3110\ : InMux
    port map (
            O => \N__15752\,
            I => \N__15728\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15751\,
            I => \N__15719\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15748\,
            I => \N__15719\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15719\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15719\
        );

    \I__3105\ : Span4Mux_h
    port map (
            O => \N__15743\,
            I => \N__15716\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15713\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15739\,
            I => \N__15708\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15708\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__15733\,
            I => \N__15701\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__15728\,
            I => \N__15701\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__15719\,
            I => \N__15701\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__15716\,
            I => \DEBUG_c_3\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__15713\,
            I => \DEBUG_c_3\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__15708\,
            I => \DEBUG_c_3\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__15701\,
            I => \DEBUG_c_3\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15692\,
            I => \receive_module.n3335\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__3091\ : Span4Mux_h
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__15680\,
            I => \receive_module.n123\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15673\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15670\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15673\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15670\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15665\,
            I => \bfn_14_13_0_\
        );

    \I__3084\ : InMux
    port map (
            O => \N__15662\,
            I => \N__15656\
        );

    \I__3083\ : InMux
    port map (
            O => \N__15661\,
            I => \N__15649\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15660\,
            I => \N__15649\
        );

    \I__3081\ : InMux
    port map (
            O => \N__15659\,
            I => \N__15649\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__15656\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__15649\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__3078\ : InMux
    port map (
            O => \N__15644\,
            I => \transmit_module.video_signal_controller.n3366\
        );

    \I__3077\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15635\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15628\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15639\,
            I => \N__15628\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15628\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15635\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__15628\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15623\,
            I => \transmit_module.video_signal_controller.n3367\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__15620\,
            I => \N__15615\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15619\,
            I => \N__15611\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15604\
        );

    \I__3067\ : InMux
    port map (
            O => \N__15615\,
            I => \N__15604\
        );

    \I__3066\ : InMux
    port map (
            O => \N__15614\,
            I => \N__15604\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__15611\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__15604\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15599\,
            I => \transmit_module.video_signal_controller.n3368\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__15596\,
            I => \N__15592\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__15595\,
            I => \N__15589\
        );

    \I__3060\ : CascadeBuf
    port map (
            O => \N__15592\,
            I => \N__15586\
        );

    \I__3059\ : CascadeBuf
    port map (
            O => \N__15589\,
            I => \N__15583\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__15586\,
            I => \N__15580\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__15583\,
            I => \N__15577\
        );

    \I__3056\ : CascadeBuf
    port map (
            O => \N__15580\,
            I => \N__15574\
        );

    \I__3055\ : CascadeBuf
    port map (
            O => \N__15577\,
            I => \N__15571\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__15574\,
            I => \N__15568\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__15571\,
            I => \N__15565\
        );

    \I__3052\ : CascadeBuf
    port map (
            O => \N__15568\,
            I => \N__15562\
        );

    \I__3051\ : CascadeBuf
    port map (
            O => \N__15565\,
            I => \N__15559\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__15562\,
            I => \N__15556\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__15559\,
            I => \N__15553\
        );

    \I__3048\ : CascadeBuf
    port map (
            O => \N__15556\,
            I => \N__15550\
        );

    \I__3047\ : CascadeBuf
    port map (
            O => \N__15553\,
            I => \N__15547\
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__15550\,
            I => \N__15544\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__15547\,
            I => \N__15541\
        );

    \I__3044\ : CascadeBuf
    port map (
            O => \N__15544\,
            I => \N__15538\
        );

    \I__3043\ : CascadeBuf
    port map (
            O => \N__15541\,
            I => \N__15535\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__15538\,
            I => \N__15532\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__15535\,
            I => \N__15529\
        );

    \I__3040\ : CascadeBuf
    port map (
            O => \N__15532\,
            I => \N__15526\
        );

    \I__3039\ : CascadeBuf
    port map (
            O => \N__15529\,
            I => \N__15523\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__15526\,
            I => \N__15520\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__15523\,
            I => \N__15517\
        );

    \I__3036\ : CascadeBuf
    port map (
            O => \N__15520\,
            I => \N__15514\
        );

    \I__3035\ : CascadeBuf
    port map (
            O => \N__15517\,
            I => \N__15511\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__15514\,
            I => \N__15508\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__15511\,
            I => \N__15505\
        );

    \I__3032\ : CascadeBuf
    port map (
            O => \N__15508\,
            I => \N__15502\
        );

    \I__3031\ : CascadeBuf
    port map (
            O => \N__15505\,
            I => \N__15499\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__15502\,
            I => \N__15496\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__15499\,
            I => \N__15493\
        );

    \I__3028\ : CascadeBuf
    port map (
            O => \N__15496\,
            I => \N__15490\
        );

    \I__3027\ : CascadeBuf
    port map (
            O => \N__15493\,
            I => \N__15487\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__15490\,
            I => \N__15484\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__15487\,
            I => \N__15481\
        );

    \I__3024\ : CascadeBuf
    port map (
            O => \N__15484\,
            I => \N__15478\
        );

    \I__3023\ : CascadeBuf
    port map (
            O => \N__15481\,
            I => \N__15475\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__15478\,
            I => \N__15472\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__15475\,
            I => \N__15469\
        );

    \I__3020\ : CascadeBuf
    port map (
            O => \N__15472\,
            I => \N__15466\
        );

    \I__3019\ : CascadeBuf
    port map (
            O => \N__15469\,
            I => \N__15463\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__15466\,
            I => \N__15460\
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__15463\,
            I => \N__15457\
        );

    \I__3016\ : CascadeBuf
    port map (
            O => \N__15460\,
            I => \N__15454\
        );

    \I__3015\ : CascadeBuf
    port map (
            O => \N__15457\,
            I => \N__15451\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__15454\,
            I => \N__15448\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__15451\,
            I => \N__15445\
        );

    \I__3012\ : CascadeBuf
    port map (
            O => \N__15448\,
            I => \N__15442\
        );

    \I__3011\ : CascadeBuf
    port map (
            O => \N__15445\,
            I => \N__15439\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__15442\,
            I => \N__15436\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__15439\,
            I => \N__15433\
        );

    \I__3008\ : CascadeBuf
    port map (
            O => \N__15436\,
            I => \N__15430\
        );

    \I__3007\ : CascadeBuf
    port map (
            O => \N__15433\,
            I => \N__15427\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__15430\,
            I => \N__15424\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__15427\,
            I => \N__15421\
        );

    \I__3004\ : CascadeBuf
    port map (
            O => \N__15424\,
            I => \N__15418\
        );

    \I__3003\ : CascadeBuf
    port map (
            O => \N__15421\,
            I => \N__15415\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__15418\,
            I => \N__15412\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__15415\,
            I => \N__15409\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15406\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15409\,
            I => \N__15403\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__15406\,
            I => \N__15400\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__15403\,
            I => \N__15397\
        );

    \I__2996\ : Span4Mux_s2_v
    port map (
            O => \N__15400\,
            I => \N__15394\
        );

    \I__2995\ : Span4Mux_s1_v
    port map (
            O => \N__15397\,
            I => \N__15391\
        );

    \I__2994\ : Span4Mux_v
    port map (
            O => \N__15394\,
            I => \N__15388\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__15391\,
            I => \N__15384\
        );

    \I__2992\ : Span4Mux_v
    port map (
            O => \N__15388\,
            I => \N__15381\
        );

    \I__2991\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15378\
        );

    \I__2990\ : Sp12to4
    port map (
            O => \N__15384\,
            I => \N__15374\
        );

    \I__2989\ : Sp12to4
    port map (
            O => \N__15381\,
            I => \N__15371\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__15378\,
            I => \N__15368\
        );

    \I__2987\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15365\
        );

    \I__2986\ : Span12Mux_s10_v
    port map (
            O => \N__15374\,
            I => \N__15360\
        );

    \I__2985\ : Span12Mux_h
    port map (
            O => \N__15371\,
            I => \N__15360\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__15368\,
            I => \RX_ADDR_2\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__15365\,
            I => \RX_ADDR_2\
        );

    \I__2982\ : Odrv12
    port map (
            O => \N__15360\,
            I => \RX_ADDR_2\
        );

    \I__2981\ : InMux
    port map (
            O => \N__15353\,
            I => \N__15350\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__15350\,
            I => \N__15347\
        );

    \I__2979\ : Span4Mux_h
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__15344\,
            I => \receive_module.n134\
        );

    \I__2977\ : InMux
    port map (
            O => \N__15341\,
            I => \receive_module.n3324\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__15338\,
            I => \N__15334\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__15337\,
            I => \N__15331\
        );

    \I__2974\ : CascadeBuf
    port map (
            O => \N__15334\,
            I => \N__15328\
        );

    \I__2973\ : CascadeBuf
    port map (
            O => \N__15331\,
            I => \N__15325\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__15328\,
            I => \N__15322\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__15325\,
            I => \N__15319\
        );

    \I__2970\ : CascadeBuf
    port map (
            O => \N__15322\,
            I => \N__15316\
        );

    \I__2969\ : CascadeBuf
    port map (
            O => \N__15319\,
            I => \N__15313\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__15316\,
            I => \N__15310\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__15313\,
            I => \N__15307\
        );

    \I__2966\ : CascadeBuf
    port map (
            O => \N__15310\,
            I => \N__15304\
        );

    \I__2965\ : CascadeBuf
    port map (
            O => \N__15307\,
            I => \N__15301\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__15304\,
            I => \N__15298\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__15301\,
            I => \N__15295\
        );

    \I__2962\ : CascadeBuf
    port map (
            O => \N__15298\,
            I => \N__15292\
        );

    \I__2961\ : CascadeBuf
    port map (
            O => \N__15295\,
            I => \N__15289\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__15292\,
            I => \N__15286\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__15289\,
            I => \N__15283\
        );

    \I__2958\ : CascadeBuf
    port map (
            O => \N__15286\,
            I => \N__15280\
        );

    \I__2957\ : CascadeBuf
    port map (
            O => \N__15283\,
            I => \N__15277\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__15280\,
            I => \N__15274\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__15277\,
            I => \N__15271\
        );

    \I__2954\ : CascadeBuf
    port map (
            O => \N__15274\,
            I => \N__15268\
        );

    \I__2953\ : CascadeBuf
    port map (
            O => \N__15271\,
            I => \N__15265\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__15268\,
            I => \N__15262\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__15265\,
            I => \N__15259\
        );

    \I__2950\ : CascadeBuf
    port map (
            O => \N__15262\,
            I => \N__15256\
        );

    \I__2949\ : CascadeBuf
    port map (
            O => \N__15259\,
            I => \N__15253\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__15256\,
            I => \N__15250\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__15253\,
            I => \N__15247\
        );

    \I__2946\ : CascadeBuf
    port map (
            O => \N__15250\,
            I => \N__15244\
        );

    \I__2945\ : CascadeBuf
    port map (
            O => \N__15247\,
            I => \N__15241\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__15244\,
            I => \N__15238\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__15241\,
            I => \N__15235\
        );

    \I__2942\ : CascadeBuf
    port map (
            O => \N__15238\,
            I => \N__15232\
        );

    \I__2941\ : CascadeBuf
    port map (
            O => \N__15235\,
            I => \N__15229\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__15232\,
            I => \N__15226\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__15229\,
            I => \N__15223\
        );

    \I__2938\ : CascadeBuf
    port map (
            O => \N__15226\,
            I => \N__15220\
        );

    \I__2937\ : CascadeBuf
    port map (
            O => \N__15223\,
            I => \N__15217\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__15220\,
            I => \N__15214\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__15217\,
            I => \N__15211\
        );

    \I__2934\ : CascadeBuf
    port map (
            O => \N__15214\,
            I => \N__15208\
        );

    \I__2933\ : CascadeBuf
    port map (
            O => \N__15211\,
            I => \N__15205\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__15208\,
            I => \N__15202\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__15205\,
            I => \N__15199\
        );

    \I__2930\ : CascadeBuf
    port map (
            O => \N__15202\,
            I => \N__15196\
        );

    \I__2929\ : CascadeBuf
    port map (
            O => \N__15199\,
            I => \N__15193\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__15196\,
            I => \N__15190\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__15193\,
            I => \N__15187\
        );

    \I__2926\ : CascadeBuf
    port map (
            O => \N__15190\,
            I => \N__15184\
        );

    \I__2925\ : CascadeBuf
    port map (
            O => \N__15187\,
            I => \N__15181\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__15184\,
            I => \N__15178\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__15181\,
            I => \N__15175\
        );

    \I__2922\ : CascadeBuf
    port map (
            O => \N__15178\,
            I => \N__15172\
        );

    \I__2921\ : CascadeBuf
    port map (
            O => \N__15175\,
            I => \N__15169\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__15172\,
            I => \N__15166\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__15169\,
            I => \N__15163\
        );

    \I__2918\ : CascadeBuf
    port map (
            O => \N__15166\,
            I => \N__15160\
        );

    \I__2917\ : CascadeBuf
    port map (
            O => \N__15163\,
            I => \N__15157\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__15160\,
            I => \N__15154\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__15157\,
            I => \N__15151\
        );

    \I__2914\ : InMux
    port map (
            O => \N__15154\,
            I => \N__15148\
        );

    \I__2913\ : InMux
    port map (
            O => \N__15151\,
            I => \N__15145\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__15148\,
            I => \N__15142\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__15145\,
            I => \N__15139\
        );

    \I__2910\ : Span4Mux_s1_v
    port map (
            O => \N__15142\,
            I => \N__15136\
        );

    \I__2909\ : Span4Mux_s1_v
    port map (
            O => \N__15139\,
            I => \N__15133\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__15136\,
            I => \N__15130\
        );

    \I__2907\ : Span4Mux_h
    port map (
            O => \N__15133\,
            I => \N__15127\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__15130\,
            I => \N__15124\
        );

    \I__2905\ : Span4Mux_h
    port map (
            O => \N__15127\,
            I => \N__15121\
        );

    \I__2904\ : Sp12to4
    port map (
            O => \N__15124\,
            I => \N__15117\
        );

    \I__2903\ : Sp12to4
    port map (
            O => \N__15121\,
            I => \N__15114\
        );

    \I__2902\ : InMux
    port map (
            O => \N__15120\,
            I => \N__15110\
        );

    \I__2901\ : Span12Mux_h
    port map (
            O => \N__15117\,
            I => \N__15105\
        );

    \I__2900\ : Span12Mux_s9_v
    port map (
            O => \N__15114\,
            I => \N__15105\
        );

    \I__2899\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15102\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__15110\,
            I => \N__15099\
        );

    \I__2897\ : Span12Mux_v
    port map (
            O => \N__15105\,
            I => \N__15096\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__15102\,
            I => \RX_ADDR_3\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__15099\,
            I => \RX_ADDR_3\
        );

    \I__2894\ : Odrv12
    port map (
            O => \N__15096\,
            I => \RX_ADDR_3\
        );

    \I__2893\ : InMux
    port map (
            O => \N__15089\,
            I => \N__15086\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__15086\,
            I => \N__15083\
        );

    \I__2891\ : Odrv12
    port map (
            O => \N__15083\,
            I => \receive_module.n133\
        );

    \I__2890\ : InMux
    port map (
            O => \N__15080\,
            I => \receive_module.n3325\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__2888\ : CascadeBuf
    port map (
            O => \N__15074\,
            I => \N__15071\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__15071\,
            I => \N__15067\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__15070\,
            I => \N__15064\
        );

    \I__2885\ : CascadeBuf
    port map (
            O => \N__15067\,
            I => \N__15061\
        );

    \I__2884\ : CascadeBuf
    port map (
            O => \N__15064\,
            I => \N__15058\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__15061\,
            I => \N__15055\
        );

    \I__2882\ : CascadeMux
    port map (
            O => \N__15058\,
            I => \N__15052\
        );

    \I__2881\ : CascadeBuf
    port map (
            O => \N__15055\,
            I => \N__15049\
        );

    \I__2880\ : CascadeBuf
    port map (
            O => \N__15052\,
            I => \N__15046\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__15049\,
            I => \N__15043\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__15046\,
            I => \N__15040\
        );

    \I__2877\ : CascadeBuf
    port map (
            O => \N__15043\,
            I => \N__15037\
        );

    \I__2876\ : CascadeBuf
    port map (
            O => \N__15040\,
            I => \N__15034\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__15037\,
            I => \N__15031\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__15034\,
            I => \N__15028\
        );

    \I__2873\ : CascadeBuf
    port map (
            O => \N__15031\,
            I => \N__15025\
        );

    \I__2872\ : CascadeBuf
    port map (
            O => \N__15028\,
            I => \N__15022\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__15025\,
            I => \N__15019\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__15022\,
            I => \N__15016\
        );

    \I__2869\ : CascadeBuf
    port map (
            O => \N__15019\,
            I => \N__15013\
        );

    \I__2868\ : CascadeBuf
    port map (
            O => \N__15016\,
            I => \N__15010\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__15013\,
            I => \N__15007\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__15010\,
            I => \N__15004\
        );

    \I__2865\ : CascadeBuf
    port map (
            O => \N__15007\,
            I => \N__15001\
        );

    \I__2864\ : CascadeBuf
    port map (
            O => \N__15004\,
            I => \N__14998\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__15001\,
            I => \N__14995\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__14998\,
            I => \N__14992\
        );

    \I__2861\ : CascadeBuf
    port map (
            O => \N__14995\,
            I => \N__14989\
        );

    \I__2860\ : CascadeBuf
    port map (
            O => \N__14992\,
            I => \N__14986\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__14989\,
            I => \N__14983\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__14986\,
            I => \N__14980\
        );

    \I__2857\ : CascadeBuf
    port map (
            O => \N__14983\,
            I => \N__14977\
        );

    \I__2856\ : CascadeBuf
    port map (
            O => \N__14980\,
            I => \N__14974\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__14977\,
            I => \N__14971\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__14974\,
            I => \N__14968\
        );

    \I__2853\ : CascadeBuf
    port map (
            O => \N__14971\,
            I => \N__14965\
        );

    \I__2852\ : CascadeBuf
    port map (
            O => \N__14968\,
            I => \N__14962\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__14965\,
            I => \N__14959\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__14962\,
            I => \N__14956\
        );

    \I__2849\ : CascadeBuf
    port map (
            O => \N__14959\,
            I => \N__14953\
        );

    \I__2848\ : CascadeBuf
    port map (
            O => \N__14956\,
            I => \N__14950\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__14953\,
            I => \N__14947\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__14950\,
            I => \N__14944\
        );

    \I__2845\ : CascadeBuf
    port map (
            O => \N__14947\,
            I => \N__14941\
        );

    \I__2844\ : CascadeBuf
    port map (
            O => \N__14944\,
            I => \N__14938\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__14941\,
            I => \N__14935\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__14938\,
            I => \N__14932\
        );

    \I__2841\ : CascadeBuf
    port map (
            O => \N__14935\,
            I => \N__14929\
        );

    \I__2840\ : CascadeBuf
    port map (
            O => \N__14932\,
            I => \N__14926\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__14929\,
            I => \N__14923\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__14926\,
            I => \N__14920\
        );

    \I__2837\ : CascadeBuf
    port map (
            O => \N__14923\,
            I => \N__14917\
        );

    \I__2836\ : CascadeBuf
    port map (
            O => \N__14920\,
            I => \N__14914\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__14917\,
            I => \N__14911\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__14914\,
            I => \N__14908\
        );

    \I__2833\ : CascadeBuf
    port map (
            O => \N__14911\,
            I => \N__14905\
        );

    \I__2832\ : CascadeBuf
    port map (
            O => \N__14908\,
            I => \N__14902\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__14905\,
            I => \N__14899\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__14902\,
            I => \N__14896\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14899\,
            I => \N__14893\
        );

    \I__2828\ : CascadeBuf
    port map (
            O => \N__14896\,
            I => \N__14890\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__14893\,
            I => \N__14887\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__14890\,
            I => \N__14884\
        );

    \I__2825\ : Span4Mux_s1_v
    port map (
            O => \N__14887\,
            I => \N__14881\
        );

    \I__2824\ : InMux
    port map (
            O => \N__14884\,
            I => \N__14878\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__14881\,
            I => \N__14875\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14878\,
            I => \N__14872\
        );

    \I__2821\ : Sp12to4
    port map (
            O => \N__14875\,
            I => \N__14867\
        );

    \I__2820\ : Span12Mux_s10_v
    port map (
            O => \N__14872\,
            I => \N__14864\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14871\,
            I => \N__14861\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14858\
        );

    \I__2817\ : Span12Mux_s10_v
    port map (
            O => \N__14867\,
            I => \N__14853\
        );

    \I__2816\ : Span12Mux_h
    port map (
            O => \N__14864\,
            I => \N__14853\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__14861\,
            I => \RX_ADDR_4\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__14858\,
            I => \RX_ADDR_4\
        );

    \I__2813\ : Odrv12
    port map (
            O => \N__14853\,
            I => \RX_ADDR_4\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__14846\,
            I => \N__14843\
        );

    \I__2811\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14840\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__14840\,
            I => \receive_module.n132\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14837\,
            I => \receive_module.n3326\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__14834\,
            I => \N__14831\
        );

    \I__2807\ : CascadeBuf
    port map (
            O => \N__14831\,
            I => \N__14828\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__14828\,
            I => \N__14824\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__14827\,
            I => \N__14821\
        );

    \I__2804\ : CascadeBuf
    port map (
            O => \N__14824\,
            I => \N__14818\
        );

    \I__2803\ : CascadeBuf
    port map (
            O => \N__14821\,
            I => \N__14815\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__14818\,
            I => \N__14812\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__14815\,
            I => \N__14809\
        );

    \I__2800\ : CascadeBuf
    port map (
            O => \N__14812\,
            I => \N__14806\
        );

    \I__2799\ : CascadeBuf
    port map (
            O => \N__14809\,
            I => \N__14803\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__14806\,
            I => \N__14800\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__14803\,
            I => \N__14797\
        );

    \I__2796\ : CascadeBuf
    port map (
            O => \N__14800\,
            I => \N__14794\
        );

    \I__2795\ : CascadeBuf
    port map (
            O => \N__14797\,
            I => \N__14791\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__14794\,
            I => \N__14788\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__14791\,
            I => \N__14785\
        );

    \I__2792\ : CascadeBuf
    port map (
            O => \N__14788\,
            I => \N__14782\
        );

    \I__2791\ : CascadeBuf
    port map (
            O => \N__14785\,
            I => \N__14779\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__14782\,
            I => \N__14776\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__14779\,
            I => \N__14773\
        );

    \I__2788\ : CascadeBuf
    port map (
            O => \N__14776\,
            I => \N__14770\
        );

    \I__2787\ : CascadeBuf
    port map (
            O => \N__14773\,
            I => \N__14767\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__14770\,
            I => \N__14764\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__14767\,
            I => \N__14761\
        );

    \I__2784\ : CascadeBuf
    port map (
            O => \N__14764\,
            I => \N__14758\
        );

    \I__2783\ : CascadeBuf
    port map (
            O => \N__14761\,
            I => \N__14755\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__14758\,
            I => \N__14752\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__14755\,
            I => \N__14749\
        );

    \I__2780\ : CascadeBuf
    port map (
            O => \N__14752\,
            I => \N__14746\
        );

    \I__2779\ : CascadeBuf
    port map (
            O => \N__14749\,
            I => \N__14743\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__14746\,
            I => \N__14740\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__14743\,
            I => \N__14737\
        );

    \I__2776\ : CascadeBuf
    port map (
            O => \N__14740\,
            I => \N__14734\
        );

    \I__2775\ : CascadeBuf
    port map (
            O => \N__14737\,
            I => \N__14731\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__14734\,
            I => \N__14728\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__14731\,
            I => \N__14725\
        );

    \I__2772\ : CascadeBuf
    port map (
            O => \N__14728\,
            I => \N__14722\
        );

    \I__2771\ : CascadeBuf
    port map (
            O => \N__14725\,
            I => \N__14719\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__14722\,
            I => \N__14716\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__14719\,
            I => \N__14713\
        );

    \I__2768\ : CascadeBuf
    port map (
            O => \N__14716\,
            I => \N__14710\
        );

    \I__2767\ : CascadeBuf
    port map (
            O => \N__14713\,
            I => \N__14707\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__14710\,
            I => \N__14704\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__14707\,
            I => \N__14701\
        );

    \I__2764\ : CascadeBuf
    port map (
            O => \N__14704\,
            I => \N__14698\
        );

    \I__2763\ : CascadeBuf
    port map (
            O => \N__14701\,
            I => \N__14695\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__14698\,
            I => \N__14692\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__14695\,
            I => \N__14689\
        );

    \I__2760\ : CascadeBuf
    port map (
            O => \N__14692\,
            I => \N__14686\
        );

    \I__2759\ : CascadeBuf
    port map (
            O => \N__14689\,
            I => \N__14683\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__14686\,
            I => \N__14680\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__14683\,
            I => \N__14677\
        );

    \I__2756\ : CascadeBuf
    port map (
            O => \N__14680\,
            I => \N__14674\
        );

    \I__2755\ : CascadeBuf
    port map (
            O => \N__14677\,
            I => \N__14671\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__14674\,
            I => \N__14668\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__14671\,
            I => \N__14665\
        );

    \I__2752\ : CascadeBuf
    port map (
            O => \N__14668\,
            I => \N__14662\
        );

    \I__2751\ : CascadeBuf
    port map (
            O => \N__14665\,
            I => \N__14659\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__14662\,
            I => \N__14656\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__14659\,
            I => \N__14653\
        );

    \I__2748\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14650\
        );

    \I__2747\ : CascadeBuf
    port map (
            O => \N__14653\,
            I => \N__14647\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__14650\,
            I => \N__14644\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__14647\,
            I => \N__14641\
        );

    \I__2744\ : Span4Mux_s2_v
    port map (
            O => \N__14644\,
            I => \N__14638\
        );

    \I__2743\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14635\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__14638\,
            I => \N__14632\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__14635\,
            I => \N__14629\
        );

    \I__2740\ : Span4Mux_h
    port map (
            O => \N__14632\,
            I => \N__14626\
        );

    \I__2739\ : Span4Mux_s2_v
    port map (
            O => \N__14629\,
            I => \N__14623\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__14626\,
            I => \N__14618\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__14623\,
            I => \N__14618\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__14618\,
            I => \N__14615\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__14615\,
            I => \N__14612\
        );

    \I__2734\ : Span4Mux_v
    port map (
            O => \N__14612\,
            I => \N__14607\
        );

    \I__2733\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14604\
        );

    \I__2732\ : InMux
    port map (
            O => \N__14610\,
            I => \N__14601\
        );

    \I__2731\ : Span4Mux_v
    port map (
            O => \N__14607\,
            I => \N__14598\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__14604\,
            I => \RX_ADDR_5\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__14601\,
            I => \RX_ADDR_5\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__14598\,
            I => \RX_ADDR_5\
        );

    \I__2727\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14588\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__14588\,
            I => \receive_module.n131\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14585\,
            I => \receive_module.n3327\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__14582\,
            I => \N__14578\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__14581\,
            I => \N__14575\
        );

    \I__2722\ : CascadeBuf
    port map (
            O => \N__14578\,
            I => \N__14572\
        );

    \I__2721\ : CascadeBuf
    port map (
            O => \N__14575\,
            I => \N__14569\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__14572\,
            I => \N__14566\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__14569\,
            I => \N__14563\
        );

    \I__2718\ : CascadeBuf
    port map (
            O => \N__14566\,
            I => \N__14560\
        );

    \I__2717\ : CascadeBuf
    port map (
            O => \N__14563\,
            I => \N__14557\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__14560\,
            I => \N__14554\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__14557\,
            I => \N__14551\
        );

    \I__2714\ : CascadeBuf
    port map (
            O => \N__14554\,
            I => \N__14548\
        );

    \I__2713\ : CascadeBuf
    port map (
            O => \N__14551\,
            I => \N__14545\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__14548\,
            I => \N__14542\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__14545\,
            I => \N__14539\
        );

    \I__2710\ : CascadeBuf
    port map (
            O => \N__14542\,
            I => \N__14536\
        );

    \I__2709\ : CascadeBuf
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__14536\,
            I => \N__14530\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__14533\,
            I => \N__14527\
        );

    \I__2706\ : CascadeBuf
    port map (
            O => \N__14530\,
            I => \N__14524\
        );

    \I__2705\ : CascadeBuf
    port map (
            O => \N__14527\,
            I => \N__14521\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__14524\,
            I => \N__14518\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__14521\,
            I => \N__14515\
        );

    \I__2702\ : CascadeBuf
    port map (
            O => \N__14518\,
            I => \N__14512\
        );

    \I__2701\ : CascadeBuf
    port map (
            O => \N__14515\,
            I => \N__14509\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__14512\,
            I => \N__14506\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__14509\,
            I => \N__14503\
        );

    \I__2698\ : CascadeBuf
    port map (
            O => \N__14506\,
            I => \N__14500\
        );

    \I__2697\ : CascadeBuf
    port map (
            O => \N__14503\,
            I => \N__14497\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__14500\,
            I => \N__14494\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__14497\,
            I => \N__14491\
        );

    \I__2694\ : CascadeBuf
    port map (
            O => \N__14494\,
            I => \N__14488\
        );

    \I__2693\ : CascadeBuf
    port map (
            O => \N__14491\,
            I => \N__14485\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__14488\,
            I => \N__14482\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__14485\,
            I => \N__14479\
        );

    \I__2690\ : CascadeBuf
    port map (
            O => \N__14482\,
            I => \N__14476\
        );

    \I__2689\ : CascadeBuf
    port map (
            O => \N__14479\,
            I => \N__14473\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__14476\,
            I => \N__14470\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__14473\,
            I => \N__14467\
        );

    \I__2686\ : CascadeBuf
    port map (
            O => \N__14470\,
            I => \N__14464\
        );

    \I__2685\ : CascadeBuf
    port map (
            O => \N__14467\,
            I => \N__14461\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__14464\,
            I => \N__14458\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__14461\,
            I => \N__14455\
        );

    \I__2682\ : CascadeBuf
    port map (
            O => \N__14458\,
            I => \N__14452\
        );

    \I__2681\ : CascadeBuf
    port map (
            O => \N__14455\,
            I => \N__14449\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__14452\,
            I => \N__14446\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__14449\,
            I => \N__14443\
        );

    \I__2678\ : CascadeBuf
    port map (
            O => \N__14446\,
            I => \N__14440\
        );

    \I__2677\ : CascadeBuf
    port map (
            O => \N__14443\,
            I => \N__14437\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__14440\,
            I => \N__14434\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__14437\,
            I => \N__14431\
        );

    \I__2674\ : CascadeBuf
    port map (
            O => \N__14434\,
            I => \N__14428\
        );

    \I__2673\ : CascadeBuf
    port map (
            O => \N__14431\,
            I => \N__14425\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__14428\,
            I => \N__14422\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__14425\,
            I => \N__14419\
        );

    \I__2670\ : CascadeBuf
    port map (
            O => \N__14422\,
            I => \N__14416\
        );

    \I__2669\ : CascadeBuf
    port map (
            O => \N__14419\,
            I => \N__14413\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__14416\,
            I => \N__14410\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__14413\,
            I => \N__14407\
        );

    \I__2666\ : CascadeBuf
    port map (
            O => \N__14410\,
            I => \N__14404\
        );

    \I__2665\ : CascadeBuf
    port map (
            O => \N__14407\,
            I => \N__14401\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__14404\,
            I => \N__14398\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__14401\,
            I => \N__14395\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14392\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14389\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__14392\,
            I => \N__14386\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__2658\ : Span12Mux_h
    port map (
            O => \N__14386\,
            I => \N__14378\
        );

    \I__2657\ : Span12Mux_v
    port map (
            O => \N__14383\,
            I => \N__14375\
        );

    \I__2656\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14372\
        );

    \I__2655\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14369\
        );

    \I__2654\ : Span12Mux_v
    port map (
            O => \N__14378\,
            I => \N__14364\
        );

    \I__2653\ : Span12Mux_h
    port map (
            O => \N__14375\,
            I => \N__14364\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__14372\,
            I => \RX_ADDR_6\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__14369\,
            I => \RX_ADDR_6\
        );

    \I__2650\ : Odrv12
    port map (
            O => \N__14364\,
            I => \RX_ADDR_6\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__14357\,
            I => \N__14354\
        );

    \I__2648\ : InMux
    port map (
            O => \N__14354\,
            I => \N__14351\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__14351\,
            I => \receive_module.n130\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14348\,
            I => \receive_module.n3328\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__14345\,
            I => \N__14341\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__14344\,
            I => \N__14338\
        );

    \I__2643\ : CascadeBuf
    port map (
            O => \N__14341\,
            I => \N__14335\
        );

    \I__2642\ : CascadeBuf
    port map (
            O => \N__14338\,
            I => \N__14332\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__14335\,
            I => \N__14329\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__14332\,
            I => \N__14326\
        );

    \I__2639\ : CascadeBuf
    port map (
            O => \N__14329\,
            I => \N__14323\
        );

    \I__2638\ : CascadeBuf
    port map (
            O => \N__14326\,
            I => \N__14320\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__14323\,
            I => \N__14317\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__14320\,
            I => \N__14314\
        );

    \I__2635\ : CascadeBuf
    port map (
            O => \N__14317\,
            I => \N__14311\
        );

    \I__2634\ : CascadeBuf
    port map (
            O => \N__14314\,
            I => \N__14308\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__14311\,
            I => \N__14305\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__14308\,
            I => \N__14302\
        );

    \I__2631\ : CascadeBuf
    port map (
            O => \N__14305\,
            I => \N__14299\
        );

    \I__2630\ : CascadeBuf
    port map (
            O => \N__14302\,
            I => \N__14296\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__14299\,
            I => \N__14293\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__14296\,
            I => \N__14290\
        );

    \I__2627\ : CascadeBuf
    port map (
            O => \N__14293\,
            I => \N__14287\
        );

    \I__2626\ : CascadeBuf
    port map (
            O => \N__14290\,
            I => \N__14284\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__14287\,
            I => \N__14281\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__14284\,
            I => \N__14278\
        );

    \I__2623\ : CascadeBuf
    port map (
            O => \N__14281\,
            I => \N__14275\
        );

    \I__2622\ : CascadeBuf
    port map (
            O => \N__14278\,
            I => \N__14272\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__14275\,
            I => \N__14269\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__14272\,
            I => \N__14266\
        );

    \I__2619\ : CascadeBuf
    port map (
            O => \N__14269\,
            I => \N__14263\
        );

    \I__2618\ : CascadeBuf
    port map (
            O => \N__14266\,
            I => \N__14260\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__14263\,
            I => \N__14257\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__14260\,
            I => \N__14254\
        );

    \I__2615\ : CascadeBuf
    port map (
            O => \N__14257\,
            I => \N__14251\
        );

    \I__2614\ : CascadeBuf
    port map (
            O => \N__14254\,
            I => \N__14248\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__14251\,
            I => \N__14245\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__14248\,
            I => \N__14242\
        );

    \I__2611\ : CascadeBuf
    port map (
            O => \N__14245\,
            I => \N__14239\
        );

    \I__2610\ : CascadeBuf
    port map (
            O => \N__14242\,
            I => \N__14236\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__14239\,
            I => \N__14233\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__14236\,
            I => \N__14230\
        );

    \I__2607\ : CascadeBuf
    port map (
            O => \N__14233\,
            I => \N__14227\
        );

    \I__2606\ : CascadeBuf
    port map (
            O => \N__14230\,
            I => \N__14224\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__14227\,
            I => \N__14221\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__14224\,
            I => \N__14218\
        );

    \I__2603\ : CascadeBuf
    port map (
            O => \N__14221\,
            I => \N__14215\
        );

    \I__2602\ : CascadeBuf
    port map (
            O => \N__14218\,
            I => \N__14212\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__14215\,
            I => \N__14209\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__14212\,
            I => \N__14206\
        );

    \I__2599\ : CascadeBuf
    port map (
            O => \N__14209\,
            I => \N__14203\
        );

    \I__2598\ : CascadeBuf
    port map (
            O => \N__14206\,
            I => \N__14200\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__14203\,
            I => \N__14197\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__14200\,
            I => \N__14194\
        );

    \I__2595\ : CascadeBuf
    port map (
            O => \N__14197\,
            I => \N__14191\
        );

    \I__2594\ : CascadeBuf
    port map (
            O => \N__14194\,
            I => \N__14188\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__14191\,
            I => \N__14185\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__14188\,
            I => \N__14182\
        );

    \I__2591\ : CascadeBuf
    port map (
            O => \N__14185\,
            I => \N__14179\
        );

    \I__2590\ : CascadeBuf
    port map (
            O => \N__14182\,
            I => \N__14176\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__14179\,
            I => \N__14173\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__14176\,
            I => \N__14170\
        );

    \I__2587\ : CascadeBuf
    port map (
            O => \N__14173\,
            I => \N__14167\
        );

    \I__2586\ : CascadeBuf
    port map (
            O => \N__14170\,
            I => \N__14164\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__14167\,
            I => \N__14161\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__14164\,
            I => \N__14158\
        );

    \I__2583\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14155\
        );

    \I__2582\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14152\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__14155\,
            I => \N__14149\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__14152\,
            I => \N__14146\
        );

    \I__2579\ : Span4Mux_s1_v
    port map (
            O => \N__14149\,
            I => \N__14143\
        );

    \I__2578\ : Span4Mux_s1_v
    port map (
            O => \N__14146\,
            I => \N__14140\
        );

    \I__2577\ : Span4Mux_h
    port map (
            O => \N__14143\,
            I => \N__14137\
        );

    \I__2576\ : Sp12to4
    port map (
            O => \N__14140\,
            I => \N__14134\
        );

    \I__2575\ : Sp12to4
    port map (
            O => \N__14137\,
            I => \N__14131\
        );

    \I__2574\ : Span12Mux_s9_v
    port map (
            O => \N__14134\,
            I => \N__14126\
        );

    \I__2573\ : Span12Mux_s9_v
    port map (
            O => \N__14131\,
            I => \N__14123\
        );

    \I__2572\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14120\
        );

    \I__2571\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14117\
        );

    \I__2570\ : Span12Mux_v
    port map (
            O => \N__14126\,
            I => \N__14112\
        );

    \I__2569\ : Span12Mux_v
    port map (
            O => \N__14123\,
            I => \N__14112\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__14120\,
            I => \RX_ADDR_7\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__14117\,
            I => \RX_ADDR_7\
        );

    \I__2566\ : Odrv12
    port map (
            O => \N__14112\,
            I => \RX_ADDR_7\
        );

    \I__2565\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14102\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__14102\,
            I => \receive_module.n129\
        );

    \I__2563\ : InMux
    port map (
            O => \N__14099\,
            I => \receive_module.n3329\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__14096\,
            I => \N__14093\
        );

    \I__2561\ : CascadeBuf
    port map (
            O => \N__14093\,
            I => \N__14089\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__14092\,
            I => \N__14086\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__14089\,
            I => \N__14083\
        );

    \I__2558\ : CascadeBuf
    port map (
            O => \N__14086\,
            I => \N__14080\
        );

    \I__2557\ : CascadeBuf
    port map (
            O => \N__14083\,
            I => \N__14077\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__14080\,
            I => \N__14074\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__14077\,
            I => \N__14071\
        );

    \I__2554\ : CascadeBuf
    port map (
            O => \N__14074\,
            I => \N__14068\
        );

    \I__2553\ : CascadeBuf
    port map (
            O => \N__14071\,
            I => \N__14065\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__14068\,
            I => \N__14062\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__14065\,
            I => \N__14059\
        );

    \I__2550\ : CascadeBuf
    port map (
            O => \N__14062\,
            I => \N__14056\
        );

    \I__2549\ : CascadeBuf
    port map (
            O => \N__14059\,
            I => \N__14053\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__14056\,
            I => \N__14050\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__14053\,
            I => \N__14047\
        );

    \I__2546\ : CascadeBuf
    port map (
            O => \N__14050\,
            I => \N__14044\
        );

    \I__2545\ : CascadeBuf
    port map (
            O => \N__14047\,
            I => \N__14041\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__14044\,
            I => \N__14038\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__2542\ : CascadeBuf
    port map (
            O => \N__14038\,
            I => \N__14032\
        );

    \I__2541\ : CascadeBuf
    port map (
            O => \N__14035\,
            I => \N__14029\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__14032\,
            I => \N__14026\
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__14029\,
            I => \N__14023\
        );

    \I__2538\ : CascadeBuf
    port map (
            O => \N__14026\,
            I => \N__14020\
        );

    \I__2537\ : CascadeBuf
    port map (
            O => \N__14023\,
            I => \N__14017\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__14020\,
            I => \N__14014\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__14017\,
            I => \N__14011\
        );

    \I__2534\ : CascadeBuf
    port map (
            O => \N__14014\,
            I => \N__14008\
        );

    \I__2533\ : CascadeBuf
    port map (
            O => \N__14011\,
            I => \N__14005\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__14008\,
            I => \N__14002\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__14005\,
            I => \N__13999\
        );

    \I__2530\ : CascadeBuf
    port map (
            O => \N__14002\,
            I => \N__13996\
        );

    \I__2529\ : CascadeBuf
    port map (
            O => \N__13999\,
            I => \N__13993\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__13996\,
            I => \N__13990\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__13993\,
            I => \N__13987\
        );

    \I__2526\ : CascadeBuf
    port map (
            O => \N__13990\,
            I => \N__13984\
        );

    \I__2525\ : CascadeBuf
    port map (
            O => \N__13987\,
            I => \N__13981\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__13984\,
            I => \N__13978\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__13981\,
            I => \N__13975\
        );

    \I__2522\ : CascadeBuf
    port map (
            O => \N__13978\,
            I => \N__13972\
        );

    \I__2521\ : CascadeBuf
    port map (
            O => \N__13975\,
            I => \N__13969\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__13972\,
            I => \N__13966\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__13969\,
            I => \N__13963\
        );

    \I__2518\ : CascadeBuf
    port map (
            O => \N__13966\,
            I => \N__13960\
        );

    \I__2517\ : CascadeBuf
    port map (
            O => \N__13963\,
            I => \N__13957\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__13960\,
            I => \N__13954\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__13957\,
            I => \N__13951\
        );

    \I__2514\ : CascadeBuf
    port map (
            O => \N__13954\,
            I => \N__13948\
        );

    \I__2513\ : CascadeBuf
    port map (
            O => \N__13951\,
            I => \N__13945\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__13948\,
            I => \N__13942\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__13945\,
            I => \N__13939\
        );

    \I__2510\ : CascadeBuf
    port map (
            O => \N__13942\,
            I => \N__13936\
        );

    \I__2509\ : CascadeBuf
    port map (
            O => \N__13939\,
            I => \N__13933\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__13936\,
            I => \N__13930\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__13933\,
            I => \N__13927\
        );

    \I__2506\ : CascadeBuf
    port map (
            O => \N__13930\,
            I => \N__13924\
        );

    \I__2505\ : CascadeBuf
    port map (
            O => \N__13927\,
            I => \N__13921\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__13924\,
            I => \N__13918\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__13921\,
            I => \N__13915\
        );

    \I__2502\ : CascadeBuf
    port map (
            O => \N__13918\,
            I => \N__13912\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13909\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__13912\,
            I => \N__13906\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__13909\,
            I => \N__13903\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13906\,
            I => \N__13900\
        );

    \I__2497\ : Span4Mux_s2_v
    port map (
            O => \N__13903\,
            I => \N__13896\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__13900\,
            I => \N__13893\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13899\,
            I => \N__13890\
        );

    \I__2494\ : Sp12to4
    port map (
            O => \N__13896\,
            I => \N__13887\
        );

    \I__2493\ : Span12Mux_s9_v
    port map (
            O => \N__13893\,
            I => \N__13884\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13890\,
            I => \N__13881\
        );

    \I__2491\ : Span12Mux_s9_v
    port map (
            O => \N__13887\,
            I => \N__13877\
        );

    \I__2490\ : Span12Mux_v
    port map (
            O => \N__13884\,
            I => \N__13874\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__13881\,
            I => \N__13871\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13868\
        );

    \I__2487\ : Span12Mux_v
    port map (
            O => \N__13877\,
            I => \N__13865\
        );

    \I__2486\ : Span12Mux_h
    port map (
            O => \N__13874\,
            I => \N__13862\
        );

    \I__2485\ : Odrv4
    port map (
            O => \N__13871\,
            I => \RX_ADDR_8\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__13868\,
            I => \RX_ADDR_8\
        );

    \I__2483\ : Odrv12
    port map (
            O => \N__13865\,
            I => \RX_ADDR_8\
        );

    \I__2482\ : Odrv12
    port map (
            O => \N__13862\,
            I => \RX_ADDR_8\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13850\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__13850\,
            I => \N__13847\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__13844\,
            I => \receive_module.n128\
        );

    \I__2477\ : InMux
    port map (
            O => \N__13841\,
            I => \bfn_14_12_0_\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__13838\,
            I => \N__13834\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__13837\,
            I => \N__13831\
        );

    \I__2474\ : CascadeBuf
    port map (
            O => \N__13834\,
            I => \N__13828\
        );

    \I__2473\ : CascadeBuf
    port map (
            O => \N__13831\,
            I => \N__13825\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__13828\,
            I => \N__13822\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__13825\,
            I => \N__13819\
        );

    \I__2470\ : CascadeBuf
    port map (
            O => \N__13822\,
            I => \N__13816\
        );

    \I__2469\ : CascadeBuf
    port map (
            O => \N__13819\,
            I => \N__13813\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__13816\,
            I => \N__13810\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__13813\,
            I => \N__13807\
        );

    \I__2466\ : CascadeBuf
    port map (
            O => \N__13810\,
            I => \N__13804\
        );

    \I__2465\ : CascadeBuf
    port map (
            O => \N__13807\,
            I => \N__13801\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__13804\,
            I => \N__13798\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__13801\,
            I => \N__13795\
        );

    \I__2462\ : CascadeBuf
    port map (
            O => \N__13798\,
            I => \N__13792\
        );

    \I__2461\ : CascadeBuf
    port map (
            O => \N__13795\,
            I => \N__13789\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__13792\,
            I => \N__13786\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__13789\,
            I => \N__13783\
        );

    \I__2458\ : CascadeBuf
    port map (
            O => \N__13786\,
            I => \N__13780\
        );

    \I__2457\ : CascadeBuf
    port map (
            O => \N__13783\,
            I => \N__13777\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__13780\,
            I => \N__13774\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__13777\,
            I => \N__13771\
        );

    \I__2454\ : CascadeBuf
    port map (
            O => \N__13774\,
            I => \N__13768\
        );

    \I__2453\ : CascadeBuf
    port map (
            O => \N__13771\,
            I => \N__13765\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__13768\,
            I => \N__13762\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__13765\,
            I => \N__13759\
        );

    \I__2450\ : CascadeBuf
    port map (
            O => \N__13762\,
            I => \N__13756\
        );

    \I__2449\ : CascadeBuf
    port map (
            O => \N__13759\,
            I => \N__13753\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__13756\,
            I => \N__13750\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__13753\,
            I => \N__13747\
        );

    \I__2446\ : CascadeBuf
    port map (
            O => \N__13750\,
            I => \N__13744\
        );

    \I__2445\ : CascadeBuf
    port map (
            O => \N__13747\,
            I => \N__13741\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__13744\,
            I => \N__13738\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__13741\,
            I => \N__13735\
        );

    \I__2442\ : CascadeBuf
    port map (
            O => \N__13738\,
            I => \N__13732\
        );

    \I__2441\ : CascadeBuf
    port map (
            O => \N__13735\,
            I => \N__13729\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__13732\,
            I => \N__13726\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__13729\,
            I => \N__13723\
        );

    \I__2438\ : CascadeBuf
    port map (
            O => \N__13726\,
            I => \N__13720\
        );

    \I__2437\ : CascadeBuf
    port map (
            O => \N__13723\,
            I => \N__13717\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__13720\,
            I => \N__13714\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__13717\,
            I => \N__13711\
        );

    \I__2434\ : CascadeBuf
    port map (
            O => \N__13714\,
            I => \N__13708\
        );

    \I__2433\ : CascadeBuf
    port map (
            O => \N__13711\,
            I => \N__13705\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__13708\,
            I => \N__13702\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__13705\,
            I => \N__13699\
        );

    \I__2430\ : CascadeBuf
    port map (
            O => \N__13702\,
            I => \N__13696\
        );

    \I__2429\ : CascadeBuf
    port map (
            O => \N__13699\,
            I => \N__13693\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__13696\,
            I => \N__13690\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__13693\,
            I => \N__13687\
        );

    \I__2426\ : CascadeBuf
    port map (
            O => \N__13690\,
            I => \N__13684\
        );

    \I__2425\ : CascadeBuf
    port map (
            O => \N__13687\,
            I => \N__13681\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__13684\,
            I => \N__13678\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__13681\,
            I => \N__13675\
        );

    \I__2422\ : CascadeBuf
    port map (
            O => \N__13678\,
            I => \N__13672\
        );

    \I__2421\ : CascadeBuf
    port map (
            O => \N__13675\,
            I => \N__13669\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__13672\,
            I => \N__13666\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__13669\,
            I => \N__13663\
        );

    \I__2418\ : CascadeBuf
    port map (
            O => \N__13666\,
            I => \N__13660\
        );

    \I__2417\ : CascadeBuf
    port map (
            O => \N__13663\,
            I => \N__13657\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__13660\,
            I => \N__13654\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__13657\,
            I => \N__13651\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13648\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13645\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__13648\,
            I => \N__13642\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__13645\,
            I => \N__13639\
        );

    \I__2410\ : Span4Mux_s3_v
    port map (
            O => \N__13642\,
            I => \N__13635\
        );

    \I__2409\ : Span4Mux_s3_v
    port map (
            O => \N__13639\,
            I => \N__13632\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13629\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__13635\,
            I => \N__13626\
        );

    \I__2406\ : Sp12to4
    port map (
            O => \N__13632\,
            I => \N__13623\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__13629\,
            I => \N__13620\
        );

    \I__2404\ : Sp12to4
    port map (
            O => \N__13626\,
            I => \N__13614\
        );

    \I__2403\ : Span12Mux_h
    port map (
            O => \N__13623\,
            I => \N__13614\
        );

    \I__2402\ : Span4Mux_h
    port map (
            O => \N__13620\,
            I => \N__13611\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13608\
        );

    \I__2400\ : Span12Mux_v
    port map (
            O => \N__13614\,
            I => \N__13605\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__13611\,
            I => \RX_ADDR_9\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__13608\,
            I => \RX_ADDR_9\
        );

    \I__2397\ : Odrv12
    port map (
            O => \N__13605\,
            I => \RX_ADDR_9\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13598\,
            I => \N__13595\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__13595\,
            I => \N__13592\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__13592\,
            I => \N__13589\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__13589\,
            I => \receive_module.n127\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13586\,
            I => \receive_module.n3331\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13579\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13582\,
            I => \N__13576\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__13579\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__13576\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13571\,
            I => \N__13567\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13564\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__13567\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__13564\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13555\
        );

    \I__2382\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13552\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__13555\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13552\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__2379\ : InMux
    port map (
            O => \N__13547\,
            I => \N__13543\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13540\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13543\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__13540\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__2375\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13531\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13528\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13531\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__13528\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13523\,
            I => \N__13519\
        );

    \I__2370\ : InMux
    port map (
            O => \N__13522\,
            I => \N__13516\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__13519\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__13516\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__13511\,
            I => \receive_module.rx_counter.n3693_cascade_\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13505\,
            I => \receive_module.rx_counter.n7\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__13502\,
            I => \receive_module.rx_counter.n11_cascade_\
        );

    \I__2363\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13493\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13493\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__13493\,
            I => \N__13490\
        );

    \I__2360\ : Odrv12
    port map (
            O => \N__13490\,
            I => \receive_module.rx_counter.PULSE_1HZ_N_94\
        );

    \I__2359\ : SRMux
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13484\,
            I => \N__13481\
        );

    \I__2357\ : Odrv12
    port map (
            O => \N__13481\,
            I => \receive_module.rx_counter.n2562\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__2355\ : CascadeBuf
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__13472\,
            I => \N__13469\
        );

    \I__2353\ : CascadeBuf
    port map (
            O => \N__13469\,
            I => \N__13465\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__13468\,
            I => \N__13462\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__13465\,
            I => \N__13459\
        );

    \I__2350\ : CascadeBuf
    port map (
            O => \N__13462\,
            I => \N__13456\
        );

    \I__2349\ : CascadeBuf
    port map (
            O => \N__13459\,
            I => \N__13453\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__13456\,
            I => \N__13450\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__13453\,
            I => \N__13447\
        );

    \I__2346\ : CascadeBuf
    port map (
            O => \N__13450\,
            I => \N__13444\
        );

    \I__2345\ : CascadeBuf
    port map (
            O => \N__13447\,
            I => \N__13441\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__13444\,
            I => \N__13438\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__13441\,
            I => \N__13435\
        );

    \I__2342\ : CascadeBuf
    port map (
            O => \N__13438\,
            I => \N__13432\
        );

    \I__2341\ : CascadeBuf
    port map (
            O => \N__13435\,
            I => \N__13429\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__13432\,
            I => \N__13426\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__13429\,
            I => \N__13423\
        );

    \I__2338\ : CascadeBuf
    port map (
            O => \N__13426\,
            I => \N__13420\
        );

    \I__2337\ : CascadeBuf
    port map (
            O => \N__13423\,
            I => \N__13417\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__13420\,
            I => \N__13414\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__13417\,
            I => \N__13411\
        );

    \I__2334\ : CascadeBuf
    port map (
            O => \N__13414\,
            I => \N__13408\
        );

    \I__2333\ : CascadeBuf
    port map (
            O => \N__13411\,
            I => \N__13405\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__13408\,
            I => \N__13402\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__13405\,
            I => \N__13399\
        );

    \I__2330\ : CascadeBuf
    port map (
            O => \N__13402\,
            I => \N__13396\
        );

    \I__2329\ : CascadeBuf
    port map (
            O => \N__13399\,
            I => \N__13393\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__13396\,
            I => \N__13390\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__13393\,
            I => \N__13387\
        );

    \I__2326\ : CascadeBuf
    port map (
            O => \N__13390\,
            I => \N__13384\
        );

    \I__2325\ : CascadeBuf
    port map (
            O => \N__13387\,
            I => \N__13381\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__13384\,
            I => \N__13378\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__13381\,
            I => \N__13375\
        );

    \I__2322\ : CascadeBuf
    port map (
            O => \N__13378\,
            I => \N__13372\
        );

    \I__2321\ : CascadeBuf
    port map (
            O => \N__13375\,
            I => \N__13369\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__13372\,
            I => \N__13366\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__13369\,
            I => \N__13363\
        );

    \I__2318\ : CascadeBuf
    port map (
            O => \N__13366\,
            I => \N__13360\
        );

    \I__2317\ : CascadeBuf
    port map (
            O => \N__13363\,
            I => \N__13357\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__13360\,
            I => \N__13354\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__13357\,
            I => \N__13351\
        );

    \I__2314\ : CascadeBuf
    port map (
            O => \N__13354\,
            I => \N__13348\
        );

    \I__2313\ : CascadeBuf
    port map (
            O => \N__13351\,
            I => \N__13345\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__13348\,
            I => \N__13342\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__13345\,
            I => \N__13339\
        );

    \I__2310\ : CascadeBuf
    port map (
            O => \N__13342\,
            I => \N__13336\
        );

    \I__2309\ : CascadeBuf
    port map (
            O => \N__13339\,
            I => \N__13333\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__13336\,
            I => \N__13330\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__13333\,
            I => \N__13327\
        );

    \I__2306\ : CascadeBuf
    port map (
            O => \N__13330\,
            I => \N__13324\
        );

    \I__2305\ : CascadeBuf
    port map (
            O => \N__13327\,
            I => \N__13321\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__13324\,
            I => \N__13318\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__13321\,
            I => \N__13315\
        );

    \I__2302\ : CascadeBuf
    port map (
            O => \N__13318\,
            I => \N__13312\
        );

    \I__2301\ : CascadeBuf
    port map (
            O => \N__13315\,
            I => \N__13309\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__13312\,
            I => \N__13306\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__13309\,
            I => \N__13303\
        );

    \I__2298\ : CascadeBuf
    port map (
            O => \N__13306\,
            I => \N__13300\
        );

    \I__2297\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13297\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__13300\,
            I => \N__13294\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__13297\,
            I => \N__13291\
        );

    \I__2294\ : CascadeBuf
    port map (
            O => \N__13294\,
            I => \N__13288\
        );

    \I__2293\ : Span4Mux_s1_v
    port map (
            O => \N__13291\,
            I => \N__13285\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__13288\,
            I => \N__13282\
        );

    \I__2291\ : Span4Mux_h
    port map (
            O => \N__13285\,
            I => \N__13279\
        );

    \I__2290\ : InMux
    port map (
            O => \N__13282\,
            I => \N__13276\
        );

    \I__2289\ : Sp12to4
    port map (
            O => \N__13279\,
            I => \N__13273\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__13276\,
            I => \N__13270\
        );

    \I__2287\ : Span12Mux_s9_v
    port map (
            O => \N__13273\,
            I => \N__13265\
        );

    \I__2286\ : Span12Mux_s9_v
    port map (
            O => \N__13270\,
            I => \N__13262\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13269\,
            I => \N__13259\
        );

    \I__2284\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13256\
        );

    \I__2283\ : Span12Mux_v
    port map (
            O => \N__13265\,
            I => \N__13253\
        );

    \I__2282\ : Span12Mux_v
    port map (
            O => \N__13262\,
            I => \N__13250\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__13259\,
            I => \RX_ADDR_0\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__13256\,
            I => \RX_ADDR_0\
        );

    \I__2279\ : Odrv12
    port map (
            O => \N__13253\,
            I => \RX_ADDR_0\
        );

    \I__2278\ : Odrv12
    port map (
            O => \N__13250\,
            I => \RX_ADDR_0\
        );

    \I__2277\ : InMux
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__13238\,
            I => \receive_module.n136\
        );

    \I__2275\ : InMux
    port map (
            O => \N__13235\,
            I => \bfn_14_11_0_\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__13232\,
            I => \N__13228\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__13231\,
            I => \N__13225\
        );

    \I__2272\ : CascadeBuf
    port map (
            O => \N__13228\,
            I => \N__13222\
        );

    \I__2271\ : CascadeBuf
    port map (
            O => \N__13225\,
            I => \N__13219\
        );

    \I__2270\ : CascadeMux
    port map (
            O => \N__13222\,
            I => \N__13216\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__13219\,
            I => \N__13213\
        );

    \I__2268\ : CascadeBuf
    port map (
            O => \N__13216\,
            I => \N__13210\
        );

    \I__2267\ : CascadeBuf
    port map (
            O => \N__13213\,
            I => \N__13207\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__13210\,
            I => \N__13204\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__13207\,
            I => \N__13201\
        );

    \I__2264\ : CascadeBuf
    port map (
            O => \N__13204\,
            I => \N__13198\
        );

    \I__2263\ : CascadeBuf
    port map (
            O => \N__13201\,
            I => \N__13195\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__13198\,
            I => \N__13192\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__13195\,
            I => \N__13189\
        );

    \I__2260\ : CascadeBuf
    port map (
            O => \N__13192\,
            I => \N__13186\
        );

    \I__2259\ : CascadeBuf
    port map (
            O => \N__13189\,
            I => \N__13183\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__13186\,
            I => \N__13180\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__13183\,
            I => \N__13177\
        );

    \I__2256\ : CascadeBuf
    port map (
            O => \N__13180\,
            I => \N__13174\
        );

    \I__2255\ : CascadeBuf
    port map (
            O => \N__13177\,
            I => \N__13171\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__13174\,
            I => \N__13168\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__13171\,
            I => \N__13165\
        );

    \I__2252\ : CascadeBuf
    port map (
            O => \N__13168\,
            I => \N__13162\
        );

    \I__2251\ : CascadeBuf
    port map (
            O => \N__13165\,
            I => \N__13159\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__13162\,
            I => \N__13156\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__13159\,
            I => \N__13153\
        );

    \I__2248\ : CascadeBuf
    port map (
            O => \N__13156\,
            I => \N__13150\
        );

    \I__2247\ : CascadeBuf
    port map (
            O => \N__13153\,
            I => \N__13147\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__13150\,
            I => \N__13144\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__13147\,
            I => \N__13141\
        );

    \I__2244\ : CascadeBuf
    port map (
            O => \N__13144\,
            I => \N__13138\
        );

    \I__2243\ : CascadeBuf
    port map (
            O => \N__13141\,
            I => \N__13135\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__13138\,
            I => \N__13132\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__13135\,
            I => \N__13129\
        );

    \I__2240\ : CascadeBuf
    port map (
            O => \N__13132\,
            I => \N__13126\
        );

    \I__2239\ : CascadeBuf
    port map (
            O => \N__13129\,
            I => \N__13123\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__13126\,
            I => \N__13120\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__13123\,
            I => \N__13117\
        );

    \I__2236\ : CascadeBuf
    port map (
            O => \N__13120\,
            I => \N__13114\
        );

    \I__2235\ : CascadeBuf
    port map (
            O => \N__13117\,
            I => \N__13111\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__13114\,
            I => \N__13108\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__13111\,
            I => \N__13105\
        );

    \I__2232\ : CascadeBuf
    port map (
            O => \N__13108\,
            I => \N__13102\
        );

    \I__2231\ : CascadeBuf
    port map (
            O => \N__13105\,
            I => \N__13099\
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__13102\,
            I => \N__13096\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__13099\,
            I => \N__13093\
        );

    \I__2228\ : CascadeBuf
    port map (
            O => \N__13096\,
            I => \N__13090\
        );

    \I__2227\ : CascadeBuf
    port map (
            O => \N__13093\,
            I => \N__13087\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__13090\,
            I => \N__13084\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__13087\,
            I => \N__13081\
        );

    \I__2224\ : CascadeBuf
    port map (
            O => \N__13084\,
            I => \N__13078\
        );

    \I__2223\ : CascadeBuf
    port map (
            O => \N__13081\,
            I => \N__13075\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__13078\,
            I => \N__13072\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__13075\,
            I => \N__13069\
        );

    \I__2220\ : CascadeBuf
    port map (
            O => \N__13072\,
            I => \N__13066\
        );

    \I__2219\ : CascadeBuf
    port map (
            O => \N__13069\,
            I => \N__13063\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__13066\,
            I => \N__13060\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__13063\,
            I => \N__13057\
        );

    \I__2216\ : CascadeBuf
    port map (
            O => \N__13060\,
            I => \N__13054\
        );

    \I__2215\ : CascadeBuf
    port map (
            O => \N__13057\,
            I => \N__13051\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__13054\,
            I => \N__13048\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__13051\,
            I => \N__13045\
        );

    \I__2212\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13042\
        );

    \I__2211\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13039\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__13042\,
            I => \N__13036\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__13039\,
            I => \N__13032\
        );

    \I__2208\ : Span4Mux_s1_v
    port map (
            O => \N__13036\,
            I => \N__13029\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__13035\,
            I => \N__13026\
        );

    \I__2206\ : Span4Mux_s1_v
    port map (
            O => \N__13032\,
            I => \N__13023\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__13029\,
            I => \N__13020\
        );

    \I__2204\ : InMux
    port map (
            O => \N__13026\,
            I => \N__13017\
        );

    \I__2203\ : Span4Mux_h
    port map (
            O => \N__13023\,
            I => \N__13014\
        );

    \I__2202\ : Span4Mux_v
    port map (
            O => \N__13020\,
            I => \N__13011\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__13017\,
            I => \N__13007\
        );

    \I__2200\ : Sp12to4
    port map (
            O => \N__13014\,
            I => \N__13004\
        );

    \I__2199\ : Sp12to4
    port map (
            O => \N__13011\,
            I => \N__13001\
        );

    \I__2198\ : InMux
    port map (
            O => \N__13010\,
            I => \N__12998\
        );

    \I__2197\ : Sp12to4
    port map (
            O => \N__13007\,
            I => \N__12993\
        );

    \I__2196\ : Span12Mux_s9_v
    port map (
            O => \N__13004\,
            I => \N__12993\
        );

    \I__2195\ : Span12Mux_s8_h
    port map (
            O => \N__13001\,
            I => \N__12990\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__12998\,
            I => \N__12983\
        );

    \I__2193\ : Span12Mux_v
    port map (
            O => \N__12993\,
            I => \N__12983\
        );

    \I__2192\ : Span12Mux_v
    port map (
            O => \N__12990\,
            I => \N__12983\
        );

    \I__2191\ : Odrv12
    port map (
            O => \N__12983\,
            I => \RX_ADDR_1\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12977\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__12974\,
            I => \receive_module.n135\
        );

    \I__2187\ : InMux
    port map (
            O => \N__12971\,
            I => \receive_module.n3323\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12968\,
            I => \transmit_module.n3348\
        );

    \I__2185\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12962\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__12962\,
            I => \N__12959\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__12959\,
            I => \transmit_module.n191\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12956\,
            I => \N__12948\
        );

    \I__2181\ : InMux
    port map (
            O => \N__12955\,
            I => \N__12948\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12954\,
            I => \N__12943\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12943\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__12948\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__12943\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__2176\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12935\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__12935\,
            I => \transmit_module.ADDR_Y_COMPONENT_8\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__12932\,
            I => \N__12928\
        );

    \I__2173\ : InMux
    port map (
            O => \N__12931\,
            I => \N__12925\
        );

    \I__2172\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12922\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12925\,
            I => \N__12919\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12922\,
            I => \N__12916\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__12919\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__12916\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__2167\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__12908\,
            I => \transmit_module.X_DELTA_PATTERN_1\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12905\,
            I => \N__12902\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__12902\,
            I => \transmit_module.X_DELTA_PATTERN_2\
        );

    \I__2163\ : InMux
    port map (
            O => \N__12899\,
            I => \N__12896\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__12896\,
            I => \transmit_module.X_DELTA_PATTERN_5\
        );

    \I__2161\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12890\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__12890\,
            I => \transmit_module.X_DELTA_PATTERN_4\
        );

    \I__2159\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12884\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__12884\,
            I => \transmit_module.X_DELTA_PATTERN_3\
        );

    \I__2157\ : CEMux
    port map (
            O => \N__12881\,
            I => \N__12875\
        );

    \I__2156\ : CEMux
    port map (
            O => \N__12880\,
            I => \N__12871\
        );

    \I__2155\ : CEMux
    port map (
            O => \N__12879\,
            I => \N__12868\
        );

    \I__2154\ : CEMux
    port map (
            O => \N__12878\,
            I => \N__12864\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__12875\,
            I => \N__12861\
        );

    \I__2152\ : CEMux
    port map (
            O => \N__12874\,
            I => \N__12858\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__12871\,
            I => \N__12855\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__12868\,
            I => \N__12852\
        );

    \I__2149\ : CEMux
    port map (
            O => \N__12867\,
            I => \N__12849\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12864\,
            I => \N__12846\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__12861\,
            I => \N__12843\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12858\,
            I => \N__12840\
        );

    \I__2145\ : Span4Mux_v
    port map (
            O => \N__12855\,
            I => \N__12833\
        );

    \I__2144\ : Span4Mux_h
    port map (
            O => \N__12852\,
            I => \N__12833\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__12849\,
            I => \N__12833\
        );

    \I__2142\ : Span4Mux_v
    port map (
            O => \N__12846\,
            I => \N__12830\
        );

    \I__2141\ : Span4Mux_h
    port map (
            O => \N__12843\,
            I => \N__12827\
        );

    \I__2140\ : Span4Mux_h
    port map (
            O => \N__12840\,
            I => \N__12822\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__12833\,
            I => \N__12822\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__12830\,
            I => \transmit_module.n2099\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__12827\,
            I => \transmit_module.n2099\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__12822\,
            I => \transmit_module.n2099\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12815\,
            I => \N__12812\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__12812\,
            I => \line_buffer.n3788\
        );

    \I__2133\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12806\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__12806\,
            I => \N__12803\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__12800\,
            I => \TX_DATA_6\
        );

    \I__2129\ : InMux
    port map (
            O => \N__12797\,
            I => \transmit_module.n3339\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12791\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__12791\,
            I => \transmit_module.n199\
        );

    \I__2126\ : InMux
    port map (
            O => \N__12788\,
            I => \transmit_module.n3340\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12785\,
            I => \N__12782\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__12782\,
            I => \transmit_module.n198\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12779\,
            I => \transmit_module.n3341\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12776\,
            I => \transmit_module.n3342\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__12773\,
            I => \N__12770\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12767\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12767\,
            I => \transmit_module.n196\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12764\,
            I => \bfn_13_19_0_\
        );

    \I__2117\ : InMux
    port map (
            O => \N__12761\,
            I => \transmit_module.n3344\
        );

    \I__2116\ : InMux
    port map (
            O => \N__12758\,
            I => \transmit_module.n3345\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12752\,
            I => \N__12749\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__12746\,
            I => \transmit_module.n193\
        );

    \I__2111\ : InMux
    port map (
            O => \N__12743\,
            I => \transmit_module.n3346\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12737\,
            I => \N__12734\
        );

    \I__2108\ : Odrv12
    port map (
            O => \N__12734\,
            I => \transmit_module.n192\
        );

    \I__2107\ : InMux
    port map (
            O => \N__12731\,
            I => \transmit_module.n3347\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12725\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__12725\,
            I => \N__12722\
        );

    \I__2104\ : Span4Mux_v
    port map (
            O => \N__12722\,
            I => \N__12719\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__12719\,
            I => \transmit_module.n187\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__12713\,
            I => \N__12710\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__12710\,
            I => \transmit_module.n219\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__12707\,
            I => \transmit_module.n187_cascade_\
        );

    \I__2098\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12701\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__12701\,
            I => \transmit_module.n218\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__12698\,
            I => \N__12695\
        );

    \I__2095\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12689\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12694\,
            I => \N__12689\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__12689\,
            I => \transmit_module.n186\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__12686\,
            I => \N__12683\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12683\,
            I => \N__12680\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__12680\,
            I => \N__12677\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__12677\,
            I => \transmit_module.n204\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__12674\,
            I => \N__12671\
        );

    \I__2087\ : InMux
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2085\ : Span4Mux_h
    port map (
            O => \N__12665\,
            I => \N__12662\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__12662\,
            I => \transmit_module.n203\
        );

    \I__2083\ : InMux
    port map (
            O => \N__12659\,
            I => \transmit_module.n3336\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__12656\,
            I => \N__12653\
        );

    \I__2081\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12650\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__12650\,
            I => \N__12647\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__12647\,
            I => \transmit_module.n202\
        );

    \I__2078\ : InMux
    port map (
            O => \N__12644\,
            I => \transmit_module.n3337\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12641\,
            I => \transmit_module.n3338\
        );

    \I__2076\ : IoInMux
    port map (
            O => \N__12638\,
            I => \N__12633\
        );

    \I__2075\ : IoInMux
    port map (
            O => \N__12637\,
            I => \N__12630\
        );

    \I__2074\ : IoInMux
    port map (
            O => \N__12636\,
            I => \N__12627\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__12633\,
            I => \N__12624\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__12630\,
            I => \N__12621\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__12627\,
            I => \N__12618\
        );

    \I__2070\ : Span4Mux_s2_v
    port map (
            O => \N__12624\,
            I => \N__12615\
        );

    \I__2069\ : Span4Mux_s2_v
    port map (
            O => \N__12621\,
            I => \N__12612\
        );

    \I__2068\ : Span4Mux_s0_h
    port map (
            O => \N__12618\,
            I => \N__12609\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__12615\,
            I => \N__12606\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__12612\,
            I => \N__12603\
        );

    \I__2065\ : Sp12to4
    port map (
            O => \N__12609\,
            I => \N__12600\
        );

    \I__2064\ : Sp12to4
    port map (
            O => \N__12606\,
            I => \N__12597\
        );

    \I__2063\ : Sp12to4
    port map (
            O => \N__12603\,
            I => \N__12594\
        );

    \I__2062\ : Span12Mux_v
    port map (
            O => \N__12600\,
            I => \N__12591\
        );

    \I__2061\ : Span12Mux_h
    port map (
            O => \N__12597\,
            I => \N__12584\
        );

    \I__2060\ : Span12Mux_h
    port map (
            O => \N__12594\,
            I => \N__12584\
        );

    \I__2059\ : Span12Mux_h
    port map (
            O => \N__12591\,
            I => \N__12584\
        );

    \I__2058\ : Odrv12
    port map (
            O => \N__12584\,
            I => n1848
        );

    \I__2057\ : IoInMux
    port map (
            O => \N__12581\,
            I => \N__12576\
        );

    \I__2056\ : IoInMux
    port map (
            O => \N__12580\,
            I => \N__12573\
        );

    \I__2055\ : IoInMux
    port map (
            O => \N__12579\,
            I => \N__12570\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__12576\,
            I => \N__12567\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__12573\,
            I => \N__12564\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__12570\,
            I => \N__12561\
        );

    \I__2051\ : Span4Mux_s1_v
    port map (
            O => \N__12567\,
            I => \N__12558\
        );

    \I__2050\ : IoSpan4Mux
    port map (
            O => \N__12564\,
            I => \N__12555\
        );

    \I__2049\ : Span4Mux_s1_h
    port map (
            O => \N__12561\,
            I => \N__12552\
        );

    \I__2048\ : Span4Mux_v
    port map (
            O => \N__12558\,
            I => \N__12549\
        );

    \I__2047\ : Span4Mux_s3_v
    port map (
            O => \N__12555\,
            I => \N__12546\
        );

    \I__2046\ : Span4Mux_h
    port map (
            O => \N__12552\,
            I => \N__12543\
        );

    \I__2045\ : Sp12to4
    port map (
            O => \N__12549\,
            I => \N__12540\
        );

    \I__2044\ : Sp12to4
    port map (
            O => \N__12546\,
            I => \N__12535\
        );

    \I__2043\ : Sp12to4
    port map (
            O => \N__12543\,
            I => \N__12535\
        );

    \I__2042\ : Span12Mux_h
    port map (
            O => \N__12540\,
            I => \N__12532\
        );

    \I__2041\ : Span12Mux_v
    port map (
            O => \N__12535\,
            I => \N__12529\
        );

    \I__2040\ : Odrv12
    port map (
            O => \N__12532\,
            I => n1847
        );

    \I__2039\ : Odrv12
    port map (
            O => \N__12529\,
            I => n1847
        );

    \I__2038\ : IoInMux
    port map (
            O => \N__12524\,
            I => \N__12520\
        );

    \I__2037\ : IoInMux
    port map (
            O => \N__12523\,
            I => \N__12517\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__12520\,
            I => \N__12513\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__12517\,
            I => \N__12510\
        );

    \I__2034\ : IoInMux
    port map (
            O => \N__12516\,
            I => \N__12507\
        );

    \I__2033\ : Span4Mux_s0_v
    port map (
            O => \N__12513\,
            I => \N__12504\
        );

    \I__2032\ : IoSpan4Mux
    port map (
            O => \N__12510\,
            I => \N__12501\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__12507\,
            I => \N__12498\
        );

    \I__2030\ : Sp12to4
    port map (
            O => \N__12504\,
            I => \N__12495\
        );

    \I__2029\ : IoSpan4Mux
    port map (
            O => \N__12501\,
            I => \N__12492\
        );

    \I__2028\ : Span12Mux_s4_v
    port map (
            O => \N__12498\,
            I => \N__12489\
        );

    \I__2027\ : Span12Mux_h
    port map (
            O => \N__12495\,
            I => \N__12486\
        );

    \I__2026\ : Sp12to4
    port map (
            O => \N__12492\,
            I => \N__12483\
        );

    \I__2025\ : Span12Mux_v
    port map (
            O => \N__12489\,
            I => \N__12480\
        );

    \I__2024\ : Span12Mux_v
    port map (
            O => \N__12486\,
            I => \N__12475\
        );

    \I__2023\ : Span12Mux_h
    port map (
            O => \N__12483\,
            I => \N__12475\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__12480\,
            I => n1846
        );

    \I__2021\ : Odrv12
    port map (
            O => \N__12475\,
            I => n1846
        );

    \I__2020\ : IoInMux
    port map (
            O => \N__12470\,
            I => \N__12465\
        );

    \I__2019\ : IoInMux
    port map (
            O => \N__12469\,
            I => \N__12462\
        );

    \I__2018\ : IoInMux
    port map (
            O => \N__12468\,
            I => \N__12459\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__12465\,
            I => \N__12456\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12462\,
            I => \N__12453\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__12459\,
            I => \N__12450\
        );

    \I__2014\ : Span4Mux_s2_v
    port map (
            O => \N__12456\,
            I => \N__12447\
        );

    \I__2013\ : Span12Mux_s4_v
    port map (
            O => \N__12453\,
            I => \N__12444\
        );

    \I__2012\ : Span4Mux_s3_h
    port map (
            O => \N__12450\,
            I => \N__12441\
        );

    \I__2011\ : Span4Mux_h
    port map (
            O => \N__12447\,
            I => \N__12438\
        );

    \I__2010\ : Span12Mux_v
    port map (
            O => \N__12444\,
            I => \N__12435\
        );

    \I__2009\ : Sp12to4
    port map (
            O => \N__12441\,
            I => \N__12432\
        );

    \I__2008\ : Sp12to4
    port map (
            O => \N__12438\,
            I => \N__12429\
        );

    \I__2007\ : Span12Mux_h
    port map (
            O => \N__12435\,
            I => \N__12424\
        );

    \I__2006\ : Span12Mux_v
    port map (
            O => \N__12432\,
            I => \N__12424\
        );

    \I__2005\ : Span12Mux_s11_v
    port map (
            O => \N__12429\,
            I => \N__12421\
        );

    \I__2004\ : Odrv12
    port map (
            O => \N__12424\,
            I => n1845
        );

    \I__2003\ : Odrv12
    port map (
            O => \N__12421\,
            I => n1845
        );

    \I__2002\ : IoInMux
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12413\,
            I => \N__12408\
        );

    \I__2000\ : IoInMux
    port map (
            O => \N__12412\,
            I => \N__12405\
        );

    \I__1999\ : IoInMux
    port map (
            O => \N__12411\,
            I => \N__12402\
        );

    \I__1998\ : Span4Mux_s0_v
    port map (
            O => \N__12408\,
            I => \N__12399\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12405\,
            I => \N__12396\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__12402\,
            I => \N__12393\
        );

    \I__1995\ : Span4Mux_v
    port map (
            O => \N__12399\,
            I => \N__12390\
        );

    \I__1994\ : Span4Mux_s0_h
    port map (
            O => \N__12396\,
            I => \N__12387\
        );

    \I__1993\ : IoSpan4Mux
    port map (
            O => \N__12393\,
            I => \N__12384\
        );

    \I__1992\ : Sp12to4
    port map (
            O => \N__12390\,
            I => \N__12381\
        );

    \I__1991\ : Sp12to4
    port map (
            O => \N__12387\,
            I => \N__12378\
        );

    \I__1990\ : Span4Mux_s2_v
    port map (
            O => \N__12384\,
            I => \N__12375\
        );

    \I__1989\ : Span12Mux_s9_h
    port map (
            O => \N__12381\,
            I => \N__12372\
        );

    \I__1988\ : Span12Mux_s10_v
    port map (
            O => \N__12378\,
            I => \N__12369\
        );

    \I__1987\ : Sp12to4
    port map (
            O => \N__12375\,
            I => \N__12366\
        );

    \I__1986\ : Span12Mux_v
    port map (
            O => \N__12372\,
            I => \N__12363\
        );

    \I__1985\ : Span12Mux_h
    port map (
            O => \N__12369\,
            I => \N__12358\
        );

    \I__1984\ : Span12Mux_s10_v
    port map (
            O => \N__12366\,
            I => \N__12358\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__12363\,
            I => n1844
        );

    \I__1982\ : Odrv12
    port map (
            O => \N__12358\,
            I => n1844
        );

    \I__1981\ : IoInMux
    port map (
            O => \N__12353\,
            I => \N__12350\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__12350\,
            I => \N__12346\
        );

    \I__1979\ : IoInMux
    port map (
            O => \N__12349\,
            I => \N__12342\
        );

    \I__1978\ : IoSpan4Mux
    port map (
            O => \N__12346\,
            I => \N__12339\
        );

    \I__1977\ : IoInMux
    port map (
            O => \N__12345\,
            I => \N__12336\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__12342\,
            I => \N__12333\
        );

    \I__1975\ : Span4Mux_s0_v
    port map (
            O => \N__12339\,
            I => \N__12330\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__12336\,
            I => \N__12327\
        );

    \I__1973\ : Span4Mux_s0_h
    port map (
            O => \N__12333\,
            I => \N__12324\
        );

    \I__1972\ : Span4Mux_v
    port map (
            O => \N__12330\,
            I => \N__12321\
        );

    \I__1971\ : IoSpan4Mux
    port map (
            O => \N__12327\,
            I => \N__12318\
        );

    \I__1970\ : Sp12to4
    port map (
            O => \N__12324\,
            I => \N__12315\
        );

    \I__1969\ : Sp12to4
    port map (
            O => \N__12321\,
            I => \N__12312\
        );

    \I__1968\ : Span4Mux_s3_v
    port map (
            O => \N__12318\,
            I => \N__12309\
        );

    \I__1967\ : Span12Mux_s9_v
    port map (
            O => \N__12315\,
            I => \N__12306\
        );

    \I__1966\ : Span12Mux_h
    port map (
            O => \N__12312\,
            I => \N__12301\
        );

    \I__1965\ : Sp12to4
    port map (
            O => \N__12309\,
            I => \N__12301\
        );

    \I__1964\ : Span12Mux_h
    port map (
            O => \N__12306\,
            I => \N__12298\
        );

    \I__1963\ : Span12Mux_v
    port map (
            O => \N__12301\,
            I => \N__12295\
        );

    \I__1962\ : Odrv12
    port map (
            O => \N__12298\,
            I => \ADV_B_c\
        );

    \I__1961\ : Odrv12
    port map (
            O => \N__12295\,
            I => \ADV_B_c\
        );

    \I__1960\ : SRMux
    port map (
            O => \N__12290\,
            I => \N__12287\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__12287\,
            I => \N__12284\
        );

    \I__1958\ : Span4Mux_h
    port map (
            O => \N__12284\,
            I => \N__12281\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__12281\,
            I => n2404
        );

    \I__1956\ : InMux
    port map (
            O => \N__12278\,
            I => \N__12275\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__12275\,
            I => \N__12272\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__12272\,
            I => \transmit_module.n220\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__12269\,
            I => \transmit_module.n218_cascade_\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__12266\,
            I => \N__12263\
        );

    \I__1951\ : CascadeBuf
    port map (
            O => \N__12263\,
            I => \N__12259\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__12262\,
            I => \N__12256\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__12259\,
            I => \N__12253\
        );

    \I__1948\ : CascadeBuf
    port map (
            O => \N__12256\,
            I => \N__12250\
        );

    \I__1947\ : CascadeBuf
    port map (
            O => \N__12253\,
            I => \N__12247\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__12250\,
            I => \N__12244\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__12247\,
            I => \N__12241\
        );

    \I__1944\ : CascadeBuf
    port map (
            O => \N__12244\,
            I => \N__12238\
        );

    \I__1943\ : CascadeBuf
    port map (
            O => \N__12241\,
            I => \N__12235\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__12238\,
            I => \N__12232\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__12235\,
            I => \N__12229\
        );

    \I__1940\ : CascadeBuf
    port map (
            O => \N__12232\,
            I => \N__12226\
        );

    \I__1939\ : CascadeBuf
    port map (
            O => \N__12229\,
            I => \N__12223\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \N__12220\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__12223\,
            I => \N__12217\
        );

    \I__1936\ : CascadeBuf
    port map (
            O => \N__12220\,
            I => \N__12214\
        );

    \I__1935\ : CascadeBuf
    port map (
            O => \N__12217\,
            I => \N__12211\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__12214\,
            I => \N__12208\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__12211\,
            I => \N__12205\
        );

    \I__1932\ : CascadeBuf
    port map (
            O => \N__12208\,
            I => \N__12202\
        );

    \I__1931\ : CascadeBuf
    port map (
            O => \N__12205\,
            I => \N__12199\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__12202\,
            I => \N__12196\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__12199\,
            I => \N__12193\
        );

    \I__1928\ : CascadeBuf
    port map (
            O => \N__12196\,
            I => \N__12190\
        );

    \I__1927\ : CascadeBuf
    port map (
            O => \N__12193\,
            I => \N__12187\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__12190\,
            I => \N__12184\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__12187\,
            I => \N__12181\
        );

    \I__1924\ : CascadeBuf
    port map (
            O => \N__12184\,
            I => \N__12178\
        );

    \I__1923\ : CascadeBuf
    port map (
            O => \N__12181\,
            I => \N__12175\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__12178\,
            I => \N__12172\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__12175\,
            I => \N__12169\
        );

    \I__1920\ : CascadeBuf
    port map (
            O => \N__12172\,
            I => \N__12166\
        );

    \I__1919\ : CascadeBuf
    port map (
            O => \N__12169\,
            I => \N__12163\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__12166\,
            I => \N__12160\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__12163\,
            I => \N__12157\
        );

    \I__1916\ : CascadeBuf
    port map (
            O => \N__12160\,
            I => \N__12154\
        );

    \I__1915\ : CascadeBuf
    port map (
            O => \N__12157\,
            I => \N__12151\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__12154\,
            I => \N__12148\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__12151\,
            I => \N__12145\
        );

    \I__1912\ : CascadeBuf
    port map (
            O => \N__12148\,
            I => \N__12142\
        );

    \I__1911\ : CascadeBuf
    port map (
            O => \N__12145\,
            I => \N__12139\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__12142\,
            I => \N__12136\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__12139\,
            I => \N__12133\
        );

    \I__1908\ : CascadeBuf
    port map (
            O => \N__12136\,
            I => \N__12130\
        );

    \I__1907\ : CascadeBuf
    port map (
            O => \N__12133\,
            I => \N__12127\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__12130\,
            I => \N__12124\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__12127\,
            I => \N__12121\
        );

    \I__1904\ : CascadeBuf
    port map (
            O => \N__12124\,
            I => \N__12118\
        );

    \I__1903\ : CascadeBuf
    port map (
            O => \N__12121\,
            I => \N__12115\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__12118\,
            I => \N__12112\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__12115\,
            I => \N__12109\
        );

    \I__1900\ : CascadeBuf
    port map (
            O => \N__12112\,
            I => \N__12106\
        );

    \I__1899\ : CascadeBuf
    port map (
            O => \N__12109\,
            I => \N__12103\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__12106\,
            I => \N__12100\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__12103\,
            I => \N__12097\
        );

    \I__1896\ : CascadeBuf
    port map (
            O => \N__12100\,
            I => \N__12094\
        );

    \I__1895\ : CascadeBuf
    port map (
            O => \N__12097\,
            I => \N__12091\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__12094\,
            I => \N__12088\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__12091\,
            I => \N__12085\
        );

    \I__1892\ : CascadeBuf
    port map (
            O => \N__12088\,
            I => \N__12082\
        );

    \I__1891\ : InMux
    port map (
            O => \N__12085\,
            I => \N__12079\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__12082\,
            I => \N__12076\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__12079\,
            I => \N__12073\
        );

    \I__1888\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12070\
        );

    \I__1887\ : Span12Mux_v
    port map (
            O => \N__12073\,
            I => \N__12067\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__12070\,
            I => \N__12064\
        );

    \I__1885\ : Span12Mux_h
    port map (
            O => \N__12067\,
            I => \N__12059\
        );

    \I__1884\ : Span12Mux_h
    port map (
            O => \N__12064\,
            I => \N__12059\
        );

    \I__1883\ : Span12Mux_v
    port map (
            O => \N__12059\,
            I => \N__12056\
        );

    \I__1882\ : Odrv12
    port map (
            O => \N__12056\,
            I => n26
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__12053\,
            I => \N__12050\
        );

    \I__1880\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12046\
        );

    \I__1879\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12041\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__12046\,
            I => \N__12038\
        );

    \I__1877\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12035\
        );

    \I__1876\ : InMux
    port map (
            O => \N__12044\,
            I => \N__12032\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__12041\,
            I => \transmit_module.video_signal_controller.n3857\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__12038\,
            I => \transmit_module.video_signal_controller.n3857\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__12035\,
            I => \transmit_module.video_signal_controller.n3857\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__12032\,
            I => \transmit_module.video_signal_controller.n3857\
        );

    \I__1871\ : InMux
    port map (
            O => \N__12023\,
            I => \N__12020\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__12020\,
            I => \N__12013\
        );

    \I__1869\ : InMux
    port map (
            O => \N__12019\,
            I => \N__12006\
        );

    \I__1868\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12006\
        );

    \I__1867\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12003\
        );

    \I__1866\ : InMux
    port map (
            O => \N__12016\,
            I => \N__12000\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__12013\,
            I => \N__11997\
        );

    \I__1864\ : InMux
    port map (
            O => \N__12012\,
            I => \N__11994\
        );

    \I__1863\ : InMux
    port map (
            O => \N__12011\,
            I => \N__11991\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__12006\,
            I => \N__11988\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__12003\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__12000\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__11997\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__11994\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__11991\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__11988\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__11975\,
            I => \N__11971\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__11974\,
            I => \N__11968\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11965\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11968\,
            I => \N__11962\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__11965\,
            I => \transmit_module.video_signal_controller.n3856\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__11962\,
            I => \transmit_module.video_signal_controller.n3856\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__11957\,
            I => \transmit_module.n220_cascade_\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__11954\,
            I => \N__11951\
        );

    \I__1847\ : CascadeBuf
    port map (
            O => \N__11951\,
            I => \N__11947\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__11950\,
            I => \N__11944\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__11947\,
            I => \N__11941\
        );

    \I__1844\ : CascadeBuf
    port map (
            O => \N__11944\,
            I => \N__11938\
        );

    \I__1843\ : CascadeBuf
    port map (
            O => \N__11941\,
            I => \N__11935\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__11938\,
            I => \N__11932\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__11935\,
            I => \N__11929\
        );

    \I__1840\ : CascadeBuf
    port map (
            O => \N__11932\,
            I => \N__11926\
        );

    \I__1839\ : CascadeBuf
    port map (
            O => \N__11929\,
            I => \N__11923\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__11926\,
            I => \N__11920\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__11923\,
            I => \N__11917\
        );

    \I__1836\ : CascadeBuf
    port map (
            O => \N__11920\,
            I => \N__11914\
        );

    \I__1835\ : CascadeBuf
    port map (
            O => \N__11917\,
            I => \N__11911\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__11914\,
            I => \N__11908\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__11911\,
            I => \N__11905\
        );

    \I__1832\ : CascadeBuf
    port map (
            O => \N__11908\,
            I => \N__11902\
        );

    \I__1831\ : CascadeBuf
    port map (
            O => \N__11905\,
            I => \N__11899\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__11902\,
            I => \N__11896\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__11899\,
            I => \N__11893\
        );

    \I__1828\ : CascadeBuf
    port map (
            O => \N__11896\,
            I => \N__11890\
        );

    \I__1827\ : CascadeBuf
    port map (
            O => \N__11893\,
            I => \N__11887\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__11890\,
            I => \N__11884\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__11887\,
            I => \N__11881\
        );

    \I__1824\ : CascadeBuf
    port map (
            O => \N__11884\,
            I => \N__11878\
        );

    \I__1823\ : CascadeBuf
    port map (
            O => \N__11881\,
            I => \N__11875\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__11878\,
            I => \N__11872\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__11875\,
            I => \N__11869\
        );

    \I__1820\ : CascadeBuf
    port map (
            O => \N__11872\,
            I => \N__11866\
        );

    \I__1819\ : CascadeBuf
    port map (
            O => \N__11869\,
            I => \N__11863\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__11866\,
            I => \N__11860\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__11863\,
            I => \N__11857\
        );

    \I__1816\ : CascadeBuf
    port map (
            O => \N__11860\,
            I => \N__11854\
        );

    \I__1815\ : CascadeBuf
    port map (
            O => \N__11857\,
            I => \N__11851\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__11854\,
            I => \N__11848\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__11851\,
            I => \N__11845\
        );

    \I__1812\ : CascadeBuf
    port map (
            O => \N__11848\,
            I => \N__11842\
        );

    \I__1811\ : CascadeBuf
    port map (
            O => \N__11845\,
            I => \N__11839\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__11842\,
            I => \N__11836\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__11839\,
            I => \N__11833\
        );

    \I__1808\ : CascadeBuf
    port map (
            O => \N__11836\,
            I => \N__11830\
        );

    \I__1807\ : CascadeBuf
    port map (
            O => \N__11833\,
            I => \N__11827\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__11830\,
            I => \N__11824\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__11827\,
            I => \N__11821\
        );

    \I__1804\ : CascadeBuf
    port map (
            O => \N__11824\,
            I => \N__11818\
        );

    \I__1803\ : CascadeBuf
    port map (
            O => \N__11821\,
            I => \N__11815\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__11818\,
            I => \N__11812\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__11815\,
            I => \N__11809\
        );

    \I__1800\ : CascadeBuf
    port map (
            O => \N__11812\,
            I => \N__11806\
        );

    \I__1799\ : CascadeBuf
    port map (
            O => \N__11809\,
            I => \N__11803\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__11806\,
            I => \N__11800\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__11803\,
            I => \N__11797\
        );

    \I__1796\ : CascadeBuf
    port map (
            O => \N__11800\,
            I => \N__11794\
        );

    \I__1795\ : CascadeBuf
    port map (
            O => \N__11797\,
            I => \N__11791\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__11794\,
            I => \N__11788\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__11791\,
            I => \N__11785\
        );

    \I__1792\ : CascadeBuf
    port map (
            O => \N__11788\,
            I => \N__11782\
        );

    \I__1791\ : CascadeBuf
    port map (
            O => \N__11785\,
            I => \N__11779\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__11782\,
            I => \N__11776\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__11779\,
            I => \N__11773\
        );

    \I__1788\ : CascadeBuf
    port map (
            O => \N__11776\,
            I => \N__11770\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11773\,
            I => \N__11767\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__11770\,
            I => \N__11764\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11767\,
            I => \N__11761\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11764\,
            I => \N__11758\
        );

    \I__1783\ : Span4Mux_h
    port map (
            O => \N__11761\,
            I => \N__11755\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11758\,
            I => \N__11752\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__11755\,
            I => \N__11749\
        );

    \I__1780\ : Span12Mux_s7_v
    port map (
            O => \N__11752\,
            I => \N__11746\
        );

    \I__1779\ : Sp12to4
    port map (
            O => \N__11749\,
            I => \N__11743\
        );

    \I__1778\ : Span12Mux_h
    port map (
            O => \N__11746\,
            I => \N__11738\
        );

    \I__1777\ : Span12Mux_s7_v
    port map (
            O => \N__11743\,
            I => \N__11738\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__11738\,
            I => n28
        );

    \I__1775\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11732\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__11732\,
            I => \transmit_module.BRAM_ADDR_13_N_256_13\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__11729\,
            I => \transmit_module.n219_cascade_\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__11726\,
            I => \N__11722\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__11725\,
            I => \N__11719\
        );

    \I__1770\ : CascadeBuf
    port map (
            O => \N__11722\,
            I => \N__11716\
        );

    \I__1769\ : CascadeBuf
    port map (
            O => \N__11719\,
            I => \N__11713\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__11716\,
            I => \N__11710\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__11713\,
            I => \N__11707\
        );

    \I__1766\ : CascadeBuf
    port map (
            O => \N__11710\,
            I => \N__11704\
        );

    \I__1765\ : CascadeBuf
    port map (
            O => \N__11707\,
            I => \N__11701\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__11704\,
            I => \N__11698\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__11701\,
            I => \N__11695\
        );

    \I__1762\ : CascadeBuf
    port map (
            O => \N__11698\,
            I => \N__11692\
        );

    \I__1761\ : CascadeBuf
    port map (
            O => \N__11695\,
            I => \N__11689\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__11692\,
            I => \N__11686\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__11689\,
            I => \N__11683\
        );

    \I__1758\ : CascadeBuf
    port map (
            O => \N__11686\,
            I => \N__11680\
        );

    \I__1757\ : CascadeBuf
    port map (
            O => \N__11683\,
            I => \N__11677\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__11680\,
            I => \N__11674\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__11677\,
            I => \N__11671\
        );

    \I__1754\ : CascadeBuf
    port map (
            O => \N__11674\,
            I => \N__11668\
        );

    \I__1753\ : CascadeBuf
    port map (
            O => \N__11671\,
            I => \N__11665\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__11668\,
            I => \N__11662\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__11665\,
            I => \N__11659\
        );

    \I__1750\ : CascadeBuf
    port map (
            O => \N__11662\,
            I => \N__11656\
        );

    \I__1749\ : CascadeBuf
    port map (
            O => \N__11659\,
            I => \N__11653\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__11656\,
            I => \N__11650\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__11653\,
            I => \N__11647\
        );

    \I__1746\ : CascadeBuf
    port map (
            O => \N__11650\,
            I => \N__11644\
        );

    \I__1745\ : CascadeBuf
    port map (
            O => \N__11647\,
            I => \N__11641\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11644\,
            I => \N__11638\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__11641\,
            I => \N__11635\
        );

    \I__1742\ : CascadeBuf
    port map (
            O => \N__11638\,
            I => \N__11632\
        );

    \I__1741\ : CascadeBuf
    port map (
            O => \N__11635\,
            I => \N__11629\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__11632\,
            I => \N__11626\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__11629\,
            I => \N__11623\
        );

    \I__1738\ : CascadeBuf
    port map (
            O => \N__11626\,
            I => \N__11620\
        );

    \I__1737\ : CascadeBuf
    port map (
            O => \N__11623\,
            I => \N__11617\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__11620\,
            I => \N__11614\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__11617\,
            I => \N__11611\
        );

    \I__1734\ : CascadeBuf
    port map (
            O => \N__11614\,
            I => \N__11608\
        );

    \I__1733\ : CascadeBuf
    port map (
            O => \N__11611\,
            I => \N__11605\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__11608\,
            I => \N__11602\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__11605\,
            I => \N__11599\
        );

    \I__1730\ : CascadeBuf
    port map (
            O => \N__11602\,
            I => \N__11596\
        );

    \I__1729\ : CascadeBuf
    port map (
            O => \N__11599\,
            I => \N__11593\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__11596\,
            I => \N__11590\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__11593\,
            I => \N__11587\
        );

    \I__1726\ : CascadeBuf
    port map (
            O => \N__11590\,
            I => \N__11584\
        );

    \I__1725\ : CascadeBuf
    port map (
            O => \N__11587\,
            I => \N__11581\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__11584\,
            I => \N__11578\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__11581\,
            I => \N__11575\
        );

    \I__1722\ : CascadeBuf
    port map (
            O => \N__11578\,
            I => \N__11572\
        );

    \I__1721\ : CascadeBuf
    port map (
            O => \N__11575\,
            I => \N__11569\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__11572\,
            I => \N__11566\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__11569\,
            I => \N__11563\
        );

    \I__1718\ : CascadeBuf
    port map (
            O => \N__11566\,
            I => \N__11560\
        );

    \I__1717\ : CascadeBuf
    port map (
            O => \N__11563\,
            I => \N__11557\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__11560\,
            I => \N__11554\
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__11557\,
            I => \N__11551\
        );

    \I__1714\ : CascadeBuf
    port map (
            O => \N__11554\,
            I => \N__11548\
        );

    \I__1713\ : CascadeBuf
    port map (
            O => \N__11551\,
            I => \N__11545\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__11548\,
            I => \N__11542\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__11545\,
            I => \N__11539\
        );

    \I__1710\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11536\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11539\,
            I => \N__11533\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11536\,
            I => \N__11530\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__11533\,
            I => \N__11527\
        );

    \I__1706\ : Span4Mux_h
    port map (
            O => \N__11530\,
            I => \N__11524\
        );

    \I__1705\ : Span12Mux_s11_v
    port map (
            O => \N__11527\,
            I => \N__11521\
        );

    \I__1704\ : Span4Mux_h
    port map (
            O => \N__11524\,
            I => \N__11518\
        );

    \I__1703\ : Span12Mux_h
    port map (
            O => \N__11521\,
            I => \N__11513\
        );

    \I__1702\ : Sp12to4
    port map (
            O => \N__11518\,
            I => \N__11513\
        );

    \I__1701\ : Span12Mux_s11_v
    port map (
            O => \N__11513\,
            I => \N__11510\
        );

    \I__1700\ : Odrv12
    port map (
            O => \N__11510\,
            I => n27
        );

    \I__1699\ : IoInMux
    port map (
            O => \N__11507\,
            I => \N__11503\
        );

    \I__1698\ : IoInMux
    port map (
            O => \N__11506\,
            I => \N__11500\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__11503\,
            I => \N__11497\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__11500\,
            I => \N__11493\
        );

    \I__1695\ : IoSpan4Mux
    port map (
            O => \N__11497\,
            I => \N__11490\
        );

    \I__1694\ : IoInMux
    port map (
            O => \N__11496\,
            I => \N__11487\
        );

    \I__1693\ : IoSpan4Mux
    port map (
            O => \N__11493\,
            I => \N__11484\
        );

    \I__1692\ : IoSpan4Mux
    port map (
            O => \N__11490\,
            I => \N__11479\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__11487\,
            I => \N__11479\
        );

    \I__1690\ : Span4Mux_s0_h
    port map (
            O => \N__11484\,
            I => \N__11476\
        );

    \I__1689\ : IoSpan4Mux
    port map (
            O => \N__11479\,
            I => \N__11473\
        );

    \I__1688\ : Sp12to4
    port map (
            O => \N__11476\,
            I => \N__11470\
        );

    \I__1687\ : Span4Mux_s2_v
    port map (
            O => \N__11473\,
            I => \N__11467\
        );

    \I__1686\ : Span12Mux_v
    port map (
            O => \N__11470\,
            I => \N__11464\
        );

    \I__1685\ : Sp12to4
    port map (
            O => \N__11467\,
            I => \N__11461\
        );

    \I__1684\ : Span12Mux_h
    port map (
            O => \N__11464\,
            I => \N__11456\
        );

    \I__1683\ : Span12Mux_s8_v
    port map (
            O => \N__11461\,
            I => \N__11456\
        );

    \I__1682\ : Odrv12
    port map (
            O => \N__11456\,
            I => n1850
        );

    \I__1681\ : IoInMux
    port map (
            O => \N__11453\,
            I => \N__11450\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__11450\,
            I => \N__11445\
        );

    \I__1679\ : IoInMux
    port map (
            O => \N__11449\,
            I => \N__11442\
        );

    \I__1678\ : IoInMux
    port map (
            O => \N__11448\,
            I => \N__11439\
        );

    \I__1677\ : IoSpan4Mux
    port map (
            O => \N__11445\,
            I => \N__11436\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__11442\,
            I => \N__11433\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__11439\,
            I => \N__11430\
        );

    \I__1674\ : IoSpan4Mux
    port map (
            O => \N__11436\,
            I => \N__11427\
        );

    \I__1673\ : Span4Mux_s3_h
    port map (
            O => \N__11433\,
            I => \N__11424\
        );

    \I__1672\ : Span4Mux_s3_v
    port map (
            O => \N__11430\,
            I => \N__11421\
        );

    \I__1671\ : Span4Mux_s3_v
    port map (
            O => \N__11427\,
            I => \N__11418\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__11424\,
            I => \N__11415\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__11421\,
            I => \N__11412\
        );

    \I__1668\ : Sp12to4
    port map (
            O => \N__11418\,
            I => \N__11407\
        );

    \I__1667\ : Sp12to4
    port map (
            O => \N__11415\,
            I => \N__11407\
        );

    \I__1666\ : Sp12to4
    port map (
            O => \N__11412\,
            I => \N__11404\
        );

    \I__1665\ : Span12Mux_v
    port map (
            O => \N__11407\,
            I => \N__11401\
        );

    \I__1664\ : Span12Mux_h
    port map (
            O => \N__11404\,
            I => \N__11398\
        );

    \I__1663\ : Odrv12
    port map (
            O => \N__11401\,
            I => n1849
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__11398\,
            I => n1849
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__11393\,
            I => \transmit_module.video_signal_controller.n3023_cascade_\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__11390\,
            I => \transmit_module.video_signal_controller.n3697_cascade_\
        );

    \I__1659\ : InMux
    port map (
            O => \N__11387\,
            I => \N__11384\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__11384\,
            I => \transmit_module.video_signal_controller.n8\
        );

    \I__1657\ : InMux
    port map (
            O => \N__11381\,
            I => \N__11378\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__11378\,
            I => \transmit_module.video_signal_controller.n3577\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__11375\,
            I => \transmit_module.video_signal_controller.n6_adj_568_cascade_\
        );

    \I__1654\ : InMux
    port map (
            O => \N__11372\,
            I => \N__11369\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__11369\,
            I => \transmit_module.video_signal_controller.n3603\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__11366\,
            I => \transmit_module.video_signal_controller.n6_cascade_\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11359\
        );

    \I__1650\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11356\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__11359\,
            I => \transmit_module.video_signal_controller.n3575\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__11356\,
            I => \transmit_module.video_signal_controller.n3575\
        );

    \I__1647\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11347\
        );

    \I__1646\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11344\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__11347\,
            I => \transmit_module.video_signal_controller.n2015\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__11344\,
            I => \transmit_module.video_signal_controller.n2015\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11339\,
            I => \receive_module.rx_counter.n3390\
        );

    \I__1642\ : InMux
    port map (
            O => \N__11336\,
            I => \receive_module.rx_counter.n3391\
        );

    \I__1641\ : IoInMux
    port map (
            O => \N__11333\,
            I => \N__11330\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__11330\,
            I => \N__11327\
        );

    \I__1639\ : IoSpan4Mux
    port map (
            O => \N__11327\,
            I => \N__11324\
        );

    \I__1638\ : IoSpan4Mux
    port map (
            O => \N__11324\,
            I => \N__11321\
        );

    \I__1637\ : Sp12to4
    port map (
            O => \N__11321\,
            I => \N__11305\
        );

    \I__1636\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11287\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11319\,
            I => \N__11287\
        );

    \I__1634\ : InMux
    port map (
            O => \N__11318\,
            I => \N__11287\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11317\,
            I => \N__11287\
        );

    \I__1632\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11287\
        );

    \I__1631\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11270\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11270\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11313\,
            I => \N__11270\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11312\,
            I => \N__11270\
        );

    \I__1627\ : InMux
    port map (
            O => \N__11311\,
            I => \N__11270\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11310\,
            I => \N__11270\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11309\,
            I => \N__11270\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11308\,
            I => \N__11270\
        );

    \I__1623\ : Span12Mux_h
    port map (
            O => \N__11305\,
            I => \N__11267\
        );

    \I__1622\ : InMux
    port map (
            O => \N__11304\,
            I => \N__11264\
        );

    \I__1621\ : InMux
    port map (
            O => \N__11303\,
            I => \N__11259\
        );

    \I__1620\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11259\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11250\
        );

    \I__1618\ : InMux
    port map (
            O => \N__11300\,
            I => \N__11250\
        );

    \I__1617\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11250\
        );

    \I__1616\ : InMux
    port map (
            O => \N__11298\,
            I => \N__11250\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__11287\,
            I => \N__11245\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__11270\,
            I => \N__11245\
        );

    \I__1613\ : Odrv12
    port map (
            O => \N__11267\,
            I => \DEBUG_c_5\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__11264\,
            I => \DEBUG_c_5\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__11259\,
            I => \DEBUG_c_5\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__11250\,
            I => \DEBUG_c_5\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__11245\,
            I => \DEBUG_c_5\
        );

    \I__1608\ : InMux
    port map (
            O => \N__11234\,
            I => \N__11231\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__11231\,
            I => \N__11227\
        );

    \I__1606\ : InMux
    port map (
            O => \N__11230\,
            I => \N__11222\
        );

    \I__1605\ : Span4Mux_h
    port map (
            O => \N__11227\,
            I => \N__11219\
        );

    \I__1604\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11216\
        );

    \I__1603\ : InMux
    port map (
            O => \N__11225\,
            I => \N__11213\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__11222\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__11219\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__11216\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__11213\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1598\ : InMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__11201\,
            I => \N__11196\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__11200\,
            I => \N__11193\
        );

    \I__1595\ : InMux
    port map (
            O => \N__11199\,
            I => \N__11190\
        );

    \I__1594\ : Span4Mux_h
    port map (
            O => \N__11196\,
            I => \N__11187\
        );

    \I__1593\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11184\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11190\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__11187\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__11184\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1589\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11174\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__11174\,
            I => \N__11169\
        );

    \I__1587\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11165\
        );

    \I__1586\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11162\
        );

    \I__1585\ : Span4Mux_h
    port map (
            O => \N__11169\,
            I => \N__11159\
        );

    \I__1584\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11156\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__11165\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__11162\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__11159\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__11156\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1579\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11144\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__11144\,
            I => \N__11141\
        );

    \I__1577\ : Span4Mux_v
    port map (
            O => \N__11141\,
            I => \N__11138\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__11138\,
            I => \transmit_module.video_signal_controller.n21\
        );

    \I__1575\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11131\
        );

    \I__1574\ : InMux
    port map (
            O => \N__11134\,
            I => \N__11126\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__11131\,
            I => \N__11123\
        );

    \I__1572\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11118\
        );

    \I__1571\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11118\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__11126\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__1569\ : Odrv4
    port map (
            O => \N__11123\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__11118\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__1567\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__11108\,
            I => \receive_module.rx_counter.n4\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__11105\,
            I => \N__11101\
        );

    \I__1564\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11097\
        );

    \I__1563\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11094\
        );

    \I__1562\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11090\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__11097\,
            I => \N__11085\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__11094\,
            I => \N__11085\
        );

    \I__1559\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11082\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__11090\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__11085\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__11082\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__1555\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11071\
        );

    \I__1554\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11066\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__11071\,
            I => \N__11063\
        );

    \I__1552\ : InMux
    port map (
            O => \N__11070\,
            I => \N__11058\
        );

    \I__1551\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11058\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__11066\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__11063\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__11058\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1547\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11048\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__11048\,
            I => \receive_module.rx_counter.n3657\
        );

    \I__1545\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__11042\,
            I => \receive_module.rx_counter.n3619\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__11039\,
            I => \receive_module.rx_counter.n3648_cascade_\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__11036\,
            I => \DEBUG_c_5_cascade_\
        );

    \I__1541\ : SRMux
    port map (
            O => \N__11033\,
            I => \N__11030\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__11030\,
            I => \N__11024\
        );

    \I__1539\ : SRMux
    port map (
            O => \N__11029\,
            I => \N__11021\
        );

    \I__1538\ : SRMux
    port map (
            O => \N__11028\,
            I => \N__11018\
        );

    \I__1537\ : SRMux
    port map (
            O => \N__11027\,
            I => \N__11015\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__11024\,
            I => \N__11012\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__11021\,
            I => \N__11007\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__11018\,
            I => \N__11007\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__11015\,
            I => \N__11004\
        );

    \I__1532\ : Sp12to4
    port map (
            O => \N__11012\,
            I => \N__10999\
        );

    \I__1531\ : Span12Mux_s6_v
    port map (
            O => \N__11007\,
            I => \N__10999\
        );

    \I__1530\ : Span4Mux_h
    port map (
            O => \N__11004\,
            I => \N__10996\
        );

    \I__1529\ : Span12Mux_v
    port map (
            O => \N__10999\,
            I => \N__10993\
        );

    \I__1528\ : Span4Mux_h
    port map (
            O => \N__10996\,
            I => \N__10990\
        );

    \I__1527\ : Span12Mux_h
    port map (
            O => \N__10993\,
            I => \N__10987\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__10990\,
            I => \N__10984\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__10987\,
            I => \line_buffer.n641\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__10984\,
            I => \line_buffer.n641\
        );

    \I__1523\ : SRMux
    port map (
            O => \N__10979\,
            I => \N__10974\
        );

    \I__1522\ : SRMux
    port map (
            O => \N__10978\,
            I => \N__10971\
        );

    \I__1521\ : SRMux
    port map (
            O => \N__10977\,
            I => \N__10967\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10962\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__10971\,
            I => \N__10962\
        );

    \I__1518\ : SRMux
    port map (
            O => \N__10970\,
            I => \N__10959\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10967\,
            I => \N__10956\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__10962\,
            I => \N__10951\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__10959\,
            I => \N__10951\
        );

    \I__1514\ : Sp12to4
    port map (
            O => \N__10956\,
            I => \N__10946\
        );

    \I__1513\ : Sp12to4
    port map (
            O => \N__10951\,
            I => \N__10946\
        );

    \I__1512\ : Span12Mux_v
    port map (
            O => \N__10946\,
            I => \N__10943\
        );

    \I__1511\ : Span12Mux_h
    port map (
            O => \N__10943\,
            I => \N__10940\
        );

    \I__1510\ : Odrv12
    port map (
            O => \N__10940\,
            I => \line_buffer.n609\
        );

    \I__1509\ : InMux
    port map (
            O => \N__10937\,
            I => \bfn_13_10_0_\
        );

    \I__1508\ : InMux
    port map (
            O => \N__10934\,
            I => \receive_module.rx_counter.n3387\
        );

    \I__1507\ : InMux
    port map (
            O => \N__10931\,
            I => \receive_module.rx_counter.n3388\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10928\,
            I => \receive_module.rx_counter.n3389\
        );

    \I__1505\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__10922\,
            I => \transmit_module.n212\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10913\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10913\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__10913\,
            I => \transmit_module.n180\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__10910\,
            I => \transmit_module.n212_cascade_\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10904\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10904\,
            I => \N__10901\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__10895\,
            I => \transmit_module.X_DELTA_PATTERN_9\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10889\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__10889\,
            I => \transmit_module.X_DELTA_PATTERN_8\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10883\,
            I => \transmit_module.X_DELTA_PATTERN_7\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10877\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10877\,
            I => \transmit_module.X_DELTA_PATTERN_6\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__1486\ : Span4Mux_h
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__10865\,
            I => \line_buffer.n574\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__10859\,
            I => \line_buffer.n3785\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1481\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10850\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__10850\,
            I => \N__10847\
        );

    \I__1479\ : Sp12to4
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__1478\ : Span12Mux_v
    port map (
            O => \N__10844\,
            I => \N__10841\
        );

    \I__1477\ : Span12Mux_v
    port map (
            O => \N__10841\,
            I => \N__10838\
        );

    \I__1476\ : Span12Mux_h
    port map (
            O => \N__10838\,
            I => \N__10835\
        );

    \I__1475\ : Odrv12
    port map (
            O => \N__10835\,
            I => \line_buffer.n566\
        );

    \I__1474\ : SRMux
    port map (
            O => \N__10832\,
            I => \N__10828\
        );

    \I__1473\ : SRMux
    port map (
            O => \N__10831\,
            I => \N__10825\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10828\,
            I => \N__10821\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10825\,
            I => \N__10818\
        );

    \I__1470\ : SRMux
    port map (
            O => \N__10824\,
            I => \N__10815\
        );

    \I__1469\ : Span4Mux_h
    port map (
            O => \N__10821\,
            I => \N__10811\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__10818\,
            I => \N__10806\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10815\,
            I => \N__10806\
        );

    \I__1466\ : SRMux
    port map (
            O => \N__10814\,
            I => \N__10803\
        );

    \I__1465\ : Span4Mux_v
    port map (
            O => \N__10811\,
            I => \N__10800\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__10806\,
            I => \N__10797\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10803\,
            I => \N__10794\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__10800\,
            I => \N__10787\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__10797\,
            I => \N__10787\
        );

    \I__1460\ : Span4Mux_h
    port map (
            O => \N__10794\,
            I => \N__10787\
        );

    \I__1459\ : Span4Mux_h
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__10784\,
            I => \N__10781\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__10781\,
            I => \line_buffer.n577\
        );

    \I__1456\ : SRMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__10775\,
            I => \N__10770\
        );

    \I__1454\ : SRMux
    port map (
            O => \N__10774\,
            I => \N__10767\
        );

    \I__1453\ : SRMux
    port map (
            O => \N__10773\,
            I => \N__10763\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__10770\,
            I => \N__10758\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10767\,
            I => \N__10758\
        );

    \I__1450\ : SRMux
    port map (
            O => \N__10766\,
            I => \N__10755\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__10763\,
            I => \N__10748\
        );

    \I__1448\ : Sp12to4
    port map (
            O => \N__10758\,
            I => \N__10748\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__10755\,
            I => \N__10748\
        );

    \I__1446\ : Span12Mux_v
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__1445\ : Span12Mux_h
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__1444\ : Odrv12
    port map (
            O => \N__10742\,
            I => \line_buffer.n513\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10733\
        );

    \I__1442\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10733\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__10733\,
            I => \N__10726\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10732\,
            I => \N__10723\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10720\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10717\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10714\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__10726\,
            I => \N__10711\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__10723\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__10720\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__10717\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10714\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__10711\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10690\
        );

    \I__1429\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10690\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10698\,
            I => \N__10687\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10682\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10682\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10679\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__10690\,
            I => \N__10676\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__10687\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__10682\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__10679\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__10676\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1419\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__10664\,
            I => \transmit_module.n214\
        );

    \I__1417\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10657\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10660\,
            I => \N__10654\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__10657\,
            I => \transmit_module.n182\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__10654\,
            I => \transmit_module.n182\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__10649\,
            I => \transmit_module.n214_cascade_\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__1411\ : CascadeBuf
    port map (
            O => \N__10643\,
            I => \N__10639\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__10642\,
            I => \N__10636\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__10639\,
            I => \N__10633\
        );

    \I__1408\ : CascadeBuf
    port map (
            O => \N__10636\,
            I => \N__10630\
        );

    \I__1407\ : CascadeBuf
    port map (
            O => \N__10633\,
            I => \N__10627\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__10630\,
            I => \N__10624\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__10627\,
            I => \N__10621\
        );

    \I__1404\ : CascadeBuf
    port map (
            O => \N__10624\,
            I => \N__10618\
        );

    \I__1403\ : CascadeBuf
    port map (
            O => \N__10621\,
            I => \N__10615\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__10618\,
            I => \N__10612\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__10615\,
            I => \N__10609\
        );

    \I__1400\ : CascadeBuf
    port map (
            O => \N__10612\,
            I => \N__10606\
        );

    \I__1399\ : CascadeBuf
    port map (
            O => \N__10609\,
            I => \N__10603\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__10606\,
            I => \N__10600\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__10603\,
            I => \N__10597\
        );

    \I__1396\ : CascadeBuf
    port map (
            O => \N__10600\,
            I => \N__10594\
        );

    \I__1395\ : CascadeBuf
    port map (
            O => \N__10597\,
            I => \N__10591\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__10594\,
            I => \N__10588\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__10591\,
            I => \N__10585\
        );

    \I__1392\ : CascadeBuf
    port map (
            O => \N__10588\,
            I => \N__10582\
        );

    \I__1391\ : CascadeBuf
    port map (
            O => \N__10585\,
            I => \N__10579\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10582\,
            I => \N__10576\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__10579\,
            I => \N__10573\
        );

    \I__1388\ : CascadeBuf
    port map (
            O => \N__10576\,
            I => \N__10570\
        );

    \I__1387\ : CascadeBuf
    port map (
            O => \N__10573\,
            I => \N__10567\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__10570\,
            I => \N__10564\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__10567\,
            I => \N__10561\
        );

    \I__1384\ : CascadeBuf
    port map (
            O => \N__10564\,
            I => \N__10558\
        );

    \I__1383\ : CascadeBuf
    port map (
            O => \N__10561\,
            I => \N__10555\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__10558\,
            I => \N__10552\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__10555\,
            I => \N__10549\
        );

    \I__1380\ : CascadeBuf
    port map (
            O => \N__10552\,
            I => \N__10546\
        );

    \I__1379\ : CascadeBuf
    port map (
            O => \N__10549\,
            I => \N__10543\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__10546\,
            I => \N__10540\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__10543\,
            I => \N__10537\
        );

    \I__1376\ : CascadeBuf
    port map (
            O => \N__10540\,
            I => \N__10534\
        );

    \I__1375\ : CascadeBuf
    port map (
            O => \N__10537\,
            I => \N__10531\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__10534\,
            I => \N__10528\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__10531\,
            I => \N__10525\
        );

    \I__1372\ : CascadeBuf
    port map (
            O => \N__10528\,
            I => \N__10522\
        );

    \I__1371\ : CascadeBuf
    port map (
            O => \N__10525\,
            I => \N__10519\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__10522\,
            I => \N__10516\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__10519\,
            I => \N__10513\
        );

    \I__1368\ : CascadeBuf
    port map (
            O => \N__10516\,
            I => \N__10510\
        );

    \I__1367\ : CascadeBuf
    port map (
            O => \N__10513\,
            I => \N__10507\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__10510\,
            I => \N__10504\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__10507\,
            I => \N__10501\
        );

    \I__1364\ : CascadeBuf
    port map (
            O => \N__10504\,
            I => \N__10498\
        );

    \I__1363\ : CascadeBuf
    port map (
            O => \N__10501\,
            I => \N__10495\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__10498\,
            I => \N__10492\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__10495\,
            I => \N__10489\
        );

    \I__1360\ : CascadeBuf
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__1359\ : CascadeBuf
    port map (
            O => \N__10489\,
            I => \N__10483\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__10486\,
            I => \N__10480\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__10483\,
            I => \N__10477\
        );

    \I__1356\ : CascadeBuf
    port map (
            O => \N__10480\,
            I => \N__10474\
        );

    \I__1355\ : CascadeBuf
    port map (
            O => \N__10477\,
            I => \N__10471\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__10474\,
            I => \N__10468\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__10471\,
            I => \N__10465\
        );

    \I__1352\ : CascadeBuf
    port map (
            O => \N__10468\,
            I => \N__10462\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10459\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__10462\,
            I => \N__10456\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__1348\ : InMux
    port map (
            O => \N__10456\,
            I => \N__10450\
        );

    \I__1347\ : Span4Mux_v
    port map (
            O => \N__10453\,
            I => \N__10447\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__10450\,
            I => \N__10444\
        );

    \I__1345\ : Span4Mux_h
    port map (
            O => \N__10447\,
            I => \N__10441\
        );

    \I__1344\ : Span4Mux_h
    port map (
            O => \N__10444\,
            I => \N__10438\
        );

    \I__1343\ : Sp12to4
    port map (
            O => \N__10441\,
            I => \N__10435\
        );

    \I__1342\ : Sp12to4
    port map (
            O => \N__10438\,
            I => \N__10432\
        );

    \I__1341\ : Span12Mux_h
    port map (
            O => \N__10435\,
            I => \N__10427\
        );

    \I__1340\ : Span12Mux_s5_v
    port map (
            O => \N__10432\,
            I => \N__10427\
        );

    \I__1339\ : Odrv12
    port map (
            O => \N__10427\,
            I => n20
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__10424\,
            I => \transmit_module.n215_cascade_\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__10421\,
            I => \N__10417\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__10420\,
            I => \N__10414\
        );

    \I__1335\ : CascadeBuf
    port map (
            O => \N__10417\,
            I => \N__10411\
        );

    \I__1334\ : CascadeBuf
    port map (
            O => \N__10414\,
            I => \N__10408\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__10411\,
            I => \N__10405\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__10408\,
            I => \N__10402\
        );

    \I__1331\ : CascadeBuf
    port map (
            O => \N__10405\,
            I => \N__10399\
        );

    \I__1330\ : CascadeBuf
    port map (
            O => \N__10402\,
            I => \N__10396\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__10399\,
            I => \N__10393\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__10396\,
            I => \N__10390\
        );

    \I__1327\ : CascadeBuf
    port map (
            O => \N__10393\,
            I => \N__10387\
        );

    \I__1326\ : CascadeBuf
    port map (
            O => \N__10390\,
            I => \N__10384\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__10387\,
            I => \N__10381\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__10384\,
            I => \N__10378\
        );

    \I__1323\ : CascadeBuf
    port map (
            O => \N__10381\,
            I => \N__10375\
        );

    \I__1322\ : CascadeBuf
    port map (
            O => \N__10378\,
            I => \N__10372\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__10375\,
            I => \N__10369\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__10372\,
            I => \N__10366\
        );

    \I__1319\ : CascadeBuf
    port map (
            O => \N__10369\,
            I => \N__10363\
        );

    \I__1318\ : CascadeBuf
    port map (
            O => \N__10366\,
            I => \N__10360\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__10363\,
            I => \N__10357\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__10360\,
            I => \N__10354\
        );

    \I__1315\ : CascadeBuf
    port map (
            O => \N__10357\,
            I => \N__10351\
        );

    \I__1314\ : CascadeBuf
    port map (
            O => \N__10354\,
            I => \N__10348\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__10351\,
            I => \N__10345\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__10348\,
            I => \N__10342\
        );

    \I__1311\ : CascadeBuf
    port map (
            O => \N__10345\,
            I => \N__10339\
        );

    \I__1310\ : CascadeBuf
    port map (
            O => \N__10342\,
            I => \N__10336\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__10339\,
            I => \N__10333\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__10336\,
            I => \N__10330\
        );

    \I__1307\ : CascadeBuf
    port map (
            O => \N__10333\,
            I => \N__10327\
        );

    \I__1306\ : CascadeBuf
    port map (
            O => \N__10330\,
            I => \N__10324\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__10327\,
            I => \N__10321\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__10324\,
            I => \N__10318\
        );

    \I__1303\ : CascadeBuf
    port map (
            O => \N__10321\,
            I => \N__10315\
        );

    \I__1302\ : CascadeBuf
    port map (
            O => \N__10318\,
            I => \N__10312\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__10315\,
            I => \N__10309\
        );

    \I__1300\ : CascadeMux
    port map (
            O => \N__10312\,
            I => \N__10306\
        );

    \I__1299\ : CascadeBuf
    port map (
            O => \N__10309\,
            I => \N__10303\
        );

    \I__1298\ : CascadeBuf
    port map (
            O => \N__10306\,
            I => \N__10300\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__10303\,
            I => \N__10297\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__10300\,
            I => \N__10294\
        );

    \I__1295\ : CascadeBuf
    port map (
            O => \N__10297\,
            I => \N__10291\
        );

    \I__1294\ : CascadeBuf
    port map (
            O => \N__10294\,
            I => \N__10288\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__10291\,
            I => \N__10285\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__10288\,
            I => \N__10282\
        );

    \I__1291\ : CascadeBuf
    port map (
            O => \N__10285\,
            I => \N__10279\
        );

    \I__1290\ : CascadeBuf
    port map (
            O => \N__10282\,
            I => \N__10276\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__10279\,
            I => \N__10273\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__10276\,
            I => \N__10270\
        );

    \I__1287\ : CascadeBuf
    port map (
            O => \N__10273\,
            I => \N__10267\
        );

    \I__1286\ : CascadeBuf
    port map (
            O => \N__10270\,
            I => \N__10264\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__10267\,
            I => \N__10261\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__10264\,
            I => \N__10258\
        );

    \I__1283\ : CascadeBuf
    port map (
            O => \N__10261\,
            I => \N__10255\
        );

    \I__1282\ : CascadeBuf
    port map (
            O => \N__10258\,
            I => \N__10252\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__10255\,
            I => \N__10249\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__10252\,
            I => \N__10246\
        );

    \I__1279\ : CascadeBuf
    port map (
            O => \N__10249\,
            I => \N__10243\
        );

    \I__1278\ : CascadeBuf
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__10243\,
            I => \N__10237\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__10240\,
            I => \N__10234\
        );

    \I__1275\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10231\
        );

    \I__1274\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10228\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10222\
        );

    \I__1271\ : Span12Mux_h
    port map (
            O => \N__10225\,
            I => \N__10219\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__10222\,
            I => \N__10216\
        );

    \I__1269\ : Span12Mux_v
    port map (
            O => \N__10219\,
            I => \N__10213\
        );

    \I__1268\ : Sp12to4
    port map (
            O => \N__10216\,
            I => \N__10210\
        );

    \I__1267\ : Odrv12
    port map (
            O => \N__10213\,
            I => n23
        );

    \I__1266\ : Odrv12
    port map (
            O => \N__10210\,
            I => n23
        );

    \I__1265\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10199\
        );

    \I__1264\ : InMux
    port map (
            O => \N__10204\,
            I => \N__10199\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__10199\,
            I => \N__10196\
        );

    \I__1262\ : Odrv12
    port map (
            O => \N__10196\,
            I => \transmit_module.n183\
        );

    \I__1261\ : InMux
    port map (
            O => \N__10193\,
            I => \N__10190\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__10190\,
            I => \transmit_module.n215\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__10187\,
            I => \transmit_module.n3859_cascade_\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10184\,
            I => \N__10179\
        );

    \I__1257\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10176\
        );

    \I__1256\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10173\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__10179\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__10176\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__10173\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__10166\,
            I => \transmit_module.video_signal_controller.n4_cascade_\
        );

    \I__1251\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10158\
        );

    \I__1250\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10155\
        );

    \I__1249\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10152\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__10158\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__10155\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__10152\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__10145\,
            I => \transmit_module.video_signal_controller.n23_cascade_\
        );

    \I__1244\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__10139\,
            I => \transmit_module.Y_DELTA_PATTERN_98\
        );

    \I__1242\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__10133\,
            I => \transmit_module.Y_DELTA_PATTERN_97\
        );

    \I__1240\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__10127\,
            I => \transmit_module.Y_DELTA_PATTERN_96\
        );

    \I__1238\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10120\
        );

    \I__1237\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10117\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__10120\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__10117\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10108\
        );

    \I__1233\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10105\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__10108\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__10105\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__1230\ : InMux
    port map (
            O => \N__10100\,
            I => \N__10096\
        );

    \I__1229\ : InMux
    port map (
            O => \N__10099\,
            I => \N__10093\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__10096\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__10093\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__10088\,
            I => \transmit_module.video_signal_controller.n8_adj_569_cascade_\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__10085\,
            I => \transmit_module.video_signal_controller.n3029_cascade_\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__10082\,
            I => \transmit_module.video_signal_controller.n3857_cascade_\
        );

    \I__1223\ : CEMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10071\
        );

    \I__1221\ : CEMux
    port map (
            O => \N__10075\,
            I => \N__10068\
        );

    \I__1220\ : CEMux
    port map (
            O => \N__10074\,
            I => \N__10064\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__10071\,
            I => \N__10061\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__10068\,
            I => \N__10058\
        );

    \I__1217\ : CEMux
    port map (
            O => \N__10067\,
            I => \N__10055\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__10064\,
            I => \N__10052\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__10061\,
            I => \transmit_module.n2125\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__10058\,
            I => \transmit_module.n2125\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__10055\,
            I => \transmit_module.n2125\
        );

    \I__1212\ : Odrv12
    port map (
            O => \N__10052\,
            I => \transmit_module.n2125\
        );

    \I__1211\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10040\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__10040\,
            I => \transmit_module.Y_DELTA_PATTERN_99\
        );

    \I__1209\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10034\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__10034\,
            I => \transmit_module.Y_DELTA_PATTERN_90\
        );

    \I__1207\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10028\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__10028\,
            I => \transmit_module.Y_DELTA_PATTERN_87\
        );

    \I__1205\ : InMux
    port map (
            O => \N__10025\,
            I => \N__10022\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__10022\,
            I => \transmit_module.Y_DELTA_PATTERN_89\
        );

    \I__1203\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10016\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__10016\,
            I => \transmit_module.Y_DELTA_PATTERN_88\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__10013\,
            I => \receive_module.rx_counter.n14_cascade_\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__10010\,
            I => \N__10006\
        );

    \I__1199\ : InMux
    port map (
            O => \N__10009\,
            I => \N__10002\
        );

    \I__1198\ : InMux
    port map (
            O => \N__10006\,
            I => \N__9997\
        );

    \I__1197\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9997\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__10002\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9997\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9987\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9991\,
            I => \N__9982\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9990\,
            I => \N__9982\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__9987\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__9982\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__9977\,
            I => \receive_module.rx_counter.n15_cascade_\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9971\,
            I => \receive_module.rx_counter.n3861\
        );

    \I__1186\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9962\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9957\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9957\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9954\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__9962\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__9957\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__9954\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__9944\,
            I => \receive_module.rx_counter.n10_adj_570\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9935\
        );

    \I__1176\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9932\
        );

    \I__1175\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9929\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9926\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__9935\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__9932\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__9929\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__9926\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1169\ : SRMux
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__9908\,
            I => \N__9903\
        );

    \I__1165\ : SRMux
    port map (
            O => \N__9907\,
            I => \N__9900\
        );

    \I__1164\ : SRMux
    port map (
            O => \N__9906\,
            I => \N__9897\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__9903\,
            I => \N__9893\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__9900\,
            I => \N__9890\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9887\
        );

    \I__1160\ : SRMux
    port map (
            O => \N__9896\,
            I => \N__9884\
        );

    \I__1159\ : Span4Mux_v
    port map (
            O => \N__9893\,
            I => \N__9875\
        );

    \I__1158\ : Span4Mux_v
    port map (
            O => \N__9890\,
            I => \N__9875\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__9887\,
            I => \N__9875\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__9884\,
            I => \N__9875\
        );

    \I__1155\ : Span4Mux_h
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__9872\,
            I => \line_buffer.n610\
        );

    \I__1153\ : SRMux
    port map (
            O => \N__9869\,
            I => \N__9865\
        );

    \I__1152\ : SRMux
    port map (
            O => \N__9868\,
            I => \N__9862\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9865\,
            I => \N__9856\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9862\,
            I => \N__9856\
        );

    \I__1149\ : SRMux
    port map (
            O => \N__9861\,
            I => \N__9853\
        );

    \I__1148\ : Span4Mux_s3_v
    port map (
            O => \N__9856\,
            I => \N__9847\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__9853\,
            I => \N__9847\
        );

    \I__1146\ : SRMux
    port map (
            O => \N__9852\,
            I => \N__9844\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__9847\,
            I => \N__9841\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__9844\,
            I => \N__9838\
        );

    \I__1143\ : Span4Mux_h
    port map (
            O => \N__9841\,
            I => \N__9835\
        );

    \I__1142\ : Span4Mux_v
    port map (
            O => \N__9838\,
            I => \N__9832\
        );

    \I__1141\ : Span4Mux_v
    port map (
            O => \N__9835\,
            I => \N__9829\
        );

    \I__1140\ : Span4Mux_h
    port map (
            O => \N__9832\,
            I => \N__9826\
        );

    \I__1139\ : Span4Mux_v
    port map (
            O => \N__9829\,
            I => \N__9823\
        );

    \I__1138\ : Span4Mux_h
    port map (
            O => \N__9826\,
            I => \N__9820\
        );

    \I__1137\ : Span4Mux_v
    port map (
            O => \N__9823\,
            I => \N__9815\
        );

    \I__1136\ : Span4Mux_h
    port map (
            O => \N__9820\,
            I => \N__9815\
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__9815\,
            I => \line_buffer.n512\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__9812\,
            I => \N__9808\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__9811\,
            I => \N__9805\
        );

    \I__1132\ : CascadeBuf
    port map (
            O => \N__9808\,
            I => \N__9802\
        );

    \I__1131\ : CascadeBuf
    port map (
            O => \N__9805\,
            I => \N__9799\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__9802\,
            I => \N__9796\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__9799\,
            I => \N__9793\
        );

    \I__1128\ : CascadeBuf
    port map (
            O => \N__9796\,
            I => \N__9790\
        );

    \I__1127\ : CascadeBuf
    port map (
            O => \N__9793\,
            I => \N__9787\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__9790\,
            I => \N__9784\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__9787\,
            I => \N__9781\
        );

    \I__1124\ : CascadeBuf
    port map (
            O => \N__9784\,
            I => \N__9778\
        );

    \I__1123\ : CascadeBuf
    port map (
            O => \N__9781\,
            I => \N__9775\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__9778\,
            I => \N__9772\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__9775\,
            I => \N__9769\
        );

    \I__1120\ : CascadeBuf
    port map (
            O => \N__9772\,
            I => \N__9766\
        );

    \I__1119\ : CascadeBuf
    port map (
            O => \N__9769\,
            I => \N__9763\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__9766\,
            I => \N__9760\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__9763\,
            I => \N__9757\
        );

    \I__1116\ : CascadeBuf
    port map (
            O => \N__9760\,
            I => \N__9754\
        );

    \I__1115\ : CascadeBuf
    port map (
            O => \N__9757\,
            I => \N__9751\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__9754\,
            I => \N__9748\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__9751\,
            I => \N__9745\
        );

    \I__1112\ : CascadeBuf
    port map (
            O => \N__9748\,
            I => \N__9742\
        );

    \I__1111\ : CascadeBuf
    port map (
            O => \N__9745\,
            I => \N__9739\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__9742\,
            I => \N__9736\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__9739\,
            I => \N__9733\
        );

    \I__1108\ : CascadeBuf
    port map (
            O => \N__9736\,
            I => \N__9730\
        );

    \I__1107\ : CascadeBuf
    port map (
            O => \N__9733\,
            I => \N__9727\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__9730\,
            I => \N__9724\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__9727\,
            I => \N__9721\
        );

    \I__1104\ : CascadeBuf
    port map (
            O => \N__9724\,
            I => \N__9718\
        );

    \I__1103\ : CascadeBuf
    port map (
            O => \N__9721\,
            I => \N__9715\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__9718\,
            I => \N__9712\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__9715\,
            I => \N__9709\
        );

    \I__1100\ : CascadeBuf
    port map (
            O => \N__9712\,
            I => \N__9706\
        );

    \I__1099\ : CascadeBuf
    port map (
            O => \N__9709\,
            I => \N__9703\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__9706\,
            I => \N__9700\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__9703\,
            I => \N__9697\
        );

    \I__1096\ : CascadeBuf
    port map (
            O => \N__9700\,
            I => \N__9694\
        );

    \I__1095\ : CascadeBuf
    port map (
            O => \N__9697\,
            I => \N__9691\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__9694\,
            I => \N__9688\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__9691\,
            I => \N__9685\
        );

    \I__1092\ : CascadeBuf
    port map (
            O => \N__9688\,
            I => \N__9682\
        );

    \I__1091\ : CascadeBuf
    port map (
            O => \N__9685\,
            I => \N__9679\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__9682\,
            I => \N__9676\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__9679\,
            I => \N__9673\
        );

    \I__1088\ : CascadeBuf
    port map (
            O => \N__9676\,
            I => \N__9670\
        );

    \I__1087\ : CascadeBuf
    port map (
            O => \N__9673\,
            I => \N__9667\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__9670\,
            I => \N__9664\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__1084\ : CascadeBuf
    port map (
            O => \N__9664\,
            I => \N__9658\
        );

    \I__1083\ : CascadeBuf
    port map (
            O => \N__9661\,
            I => \N__9655\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__9658\,
            I => \N__9652\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__9655\,
            I => \N__9649\
        );

    \I__1080\ : CascadeBuf
    port map (
            O => \N__9652\,
            I => \N__9646\
        );

    \I__1079\ : CascadeBuf
    port map (
            O => \N__9649\,
            I => \N__9643\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__9646\,
            I => \N__9640\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__9643\,
            I => \N__9637\
        );

    \I__1076\ : CascadeBuf
    port map (
            O => \N__9640\,
            I => \N__9634\
        );

    \I__1075\ : CascadeBuf
    port map (
            O => \N__9637\,
            I => \N__9631\
        );

    \I__1074\ : CascadeMux
    port map (
            O => \N__9634\,
            I => \N__9628\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__9631\,
            I => \N__9625\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9622\
        );

    \I__1071\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9619\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__9622\,
            I => \N__9616\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__9619\,
            I => \N__9613\
        );

    \I__1068\ : Span12Mux_h
    port map (
            O => \N__9616\,
            I => \N__9610\
        );

    \I__1067\ : Span12Mux_h
    port map (
            O => \N__9613\,
            I => \N__9607\
        );

    \I__1066\ : Span12Mux_v
    port map (
            O => \N__9610\,
            I => \N__9602\
        );

    \I__1065\ : Span12Mux_v
    port map (
            O => \N__9607\,
            I => \N__9602\
        );

    \I__1064\ : Odrv12
    port map (
            O => \N__9602\,
            I => n22
        );

    \I__1063\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__9596\,
            I => \transmit_module.X_DELTA_PATTERN_15\
        );

    \I__1061\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__9590\,
            I => \transmit_module.X_DELTA_PATTERN_14\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9584\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__9584\,
            I => \N__9581\
        );

    \I__1057\ : Span4Mux_v
    port map (
            O => \N__9581\,
            I => \N__9578\
        );

    \I__1056\ : Span4Mux_h
    port map (
            O => \N__9578\,
            I => \N__9575\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__9575\,
            I => \line_buffer.n630\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__9572\,
            I => \N__9569\
        );

    \I__1053\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9566\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__9566\,
            I => \N__9563\
        );

    \I__1051\ : Span4Mux_h
    port map (
            O => \N__9563\,
            I => \N__9560\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__9557\,
            I => \line_buffer.n638\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9549\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9544\
        );

    \I__1046\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9544\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9549\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9544\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1043\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9534\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9538\,
            I => \N__9531\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9528\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__9534\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__9531\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9528\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__9521\,
            I => \receive_module.rx_counter.n3619_cascade_\
        );

    \I__1036\ : SRMux
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__9515\,
            I => \N__9511\
        );

    \I__1034\ : SRMux
    port map (
            O => \N__9514\,
            I => \N__9508\
        );

    \I__1033\ : Span4Mux_v
    port map (
            O => \N__9511\,
            I => \N__9502\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__9508\,
            I => \N__9502\
        );

    \I__1031\ : SRMux
    port map (
            O => \N__9507\,
            I => \N__9499\
        );

    \I__1030\ : Span4Mux_v
    port map (
            O => \N__9502\,
            I => \N__9493\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9493\
        );

    \I__1028\ : SRMux
    port map (
            O => \N__9498\,
            I => \N__9490\
        );

    \I__1027\ : Span4Mux_v
    port map (
            O => \N__9493\,
            I => \N__9485\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__9490\,
            I => \N__9485\
        );

    \I__1025\ : Span4Mux_h
    port map (
            O => \N__9485\,
            I => \N__9482\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__9482\,
            I => \N__9479\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__9479\,
            I => \line_buffer.n642\
        );

    \I__1022\ : SRMux
    port map (
            O => \N__9476\,
            I => \N__9472\
        );

    \I__1021\ : SRMux
    port map (
            O => \N__9475\,
            I => \N__9469\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__9472\,
            I => \N__9465\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__9469\,
            I => \N__9462\
        );

    \I__1018\ : SRMux
    port map (
            O => \N__9468\,
            I => \N__9459\
        );

    \I__1017\ : Span4Mux_v
    port map (
            O => \N__9465\,
            I => \N__9455\
        );

    \I__1016\ : Span4Mux_s3_v
    port map (
            O => \N__9462\,
            I => \N__9450\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__9459\,
            I => \N__9450\
        );

    \I__1014\ : SRMux
    port map (
            O => \N__9458\,
            I => \N__9447\
        );

    \I__1013\ : Span4Mux_h
    port map (
            O => \N__9455\,
            I => \N__9444\
        );

    \I__1012\ : Span4Mux_h
    port map (
            O => \N__9450\,
            I => \N__9439\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9447\,
            I => \N__9439\
        );

    \I__1010\ : Span4Mux_v
    port map (
            O => \N__9444\,
            I => \N__9436\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__9439\,
            I => \N__9433\
        );

    \I__1008\ : Span4Mux_v
    port map (
            O => \N__9436\,
            I => \N__9428\
        );

    \I__1007\ : Span4Mux_h
    port map (
            O => \N__9433\,
            I => \N__9428\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__9428\,
            I => \line_buffer.n578\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9425\,
            I => \bfn_11_16_0_\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9422\,
            I => \transmit_module.video_signal_controller.n3385\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9419\,
            I => \transmit_module.video_signal_controller.n3386\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9413\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__9413\,
            I => \N__9410\
        );

    \I__1000\ : Odrv12
    port map (
            O => \N__9410\,
            I => \transmit_module.Y_DELTA_PATTERN_28\
        );

    \I__999\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__9404\,
            I => \transmit_module.Y_DELTA_PATTERN_29\
        );

    \I__997\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9398\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9398\,
            I => \transmit_module.Y_DELTA_PATTERN_30\
        );

    \I__995\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__9392\,
            I => \transmit_module.Y_DELTA_PATTERN_31\
        );

    \I__993\ : InMux
    port map (
            O => \N__9389\,
            I => \N__9386\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__9386\,
            I => \transmit_module.Y_DELTA_PATTERN_73\
        );

    \I__991\ : InMux
    port map (
            O => \N__9383\,
            I => \N__9380\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__989\ : Span4Mux_h
    port map (
            O => \N__9377\,
            I => \N__9374\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__9374\,
            I => \transmit_module.Y_DELTA_PATTERN_72\
        );

    \I__987\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9368\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__9368\,
            I => \transmit_module.Y_DELTA_PATTERN_92\
        );

    \I__985\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9362\,
            I => \transmit_module.Y_DELTA_PATTERN_91\
        );

    \I__983\ : InMux
    port map (
            O => \N__9359\,
            I => \bfn_11_15_0_\
        );

    \I__982\ : InMux
    port map (
            O => \N__9356\,
            I => \transmit_module.video_signal_controller.n3377\
        );

    \I__981\ : InMux
    port map (
            O => \N__9353\,
            I => \transmit_module.video_signal_controller.n3378\
        );

    \I__980\ : InMux
    port map (
            O => \N__9350\,
            I => \transmit_module.video_signal_controller.n3379\
        );

    \I__979\ : InMux
    port map (
            O => \N__9347\,
            I => \transmit_module.video_signal_controller.n3380\
        );

    \I__978\ : InMux
    port map (
            O => \N__9344\,
            I => \transmit_module.video_signal_controller.n3381\
        );

    \I__977\ : InMux
    port map (
            O => \N__9341\,
            I => \transmit_module.video_signal_controller.n3382\
        );

    \I__976\ : InMux
    port map (
            O => \N__9338\,
            I => \transmit_module.video_signal_controller.n3383\
        );

    \I__975\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9332\,
            I => \transmit_module.Y_DELTA_PATTERN_12\
        );

    \I__973\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9326\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__9326\,
            I => \transmit_module.Y_DELTA_PATTERN_11\
        );

    \I__971\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9320\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__969\ : Span4Mux_h
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__9314\,
            I => \transmit_module.Y_DELTA_PATTERN_83\
        );

    \I__967\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9308\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9308\,
            I => \transmit_module.Y_DELTA_PATTERN_84\
        );

    \I__965\ : InMux
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__9302\,
            I => \transmit_module.Y_DELTA_PATTERN_95\
        );

    \I__963\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9296\,
            I => \transmit_module.Y_DELTA_PATTERN_94\
        );

    \I__961\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9290\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__9290\,
            I => \transmit_module.Y_DELTA_PATTERN_93\
        );

    \I__959\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9284\,
            I => \transmit_module.Y_DELTA_PATTERN_85\
        );

    \I__957\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__9278\,
            I => \transmit_module.Y_DELTA_PATTERN_86\
        );

    \I__955\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9272\,
            I => \transmit_module.Y_DELTA_PATTERN_26\
        );

    \I__953\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9266\,
            I => \transmit_module.Y_DELTA_PATTERN_25\
        );

    \I__951\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__9260\,
            I => \transmit_module.Y_DELTA_PATTERN_7\
        );

    \I__949\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__9254\,
            I => \transmit_module.Y_DELTA_PATTERN_27\
        );

    \I__947\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__9248\,
            I => \transmit_module.Y_DELTA_PATTERN_10\
        );

    \I__945\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__943\ : Span4Mux_h
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__9236\,
            I => \transmit_module.Y_DELTA_PATTERN_13\
        );

    \I__941\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__9230\,
            I => \transmit_module.Y_DELTA_PATTERN_9\
        );

    \I__939\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__9224\,
            I => \transmit_module.Y_DELTA_PATTERN_8\
        );

    \I__937\ : InMux
    port map (
            O => \N__9221\,
            I => \bfn_11_9_0_\
        );

    \I__936\ : InMux
    port map (
            O => \N__9218\,
            I => \receive_module.rx_counter.n3349\
        );

    \I__935\ : InMux
    port map (
            O => \N__9215\,
            I => \receive_module.rx_counter.n3350\
        );

    \I__934\ : InMux
    port map (
            O => \N__9212\,
            I => \receive_module.rx_counter.n3351\
        );

    \I__933\ : InMux
    port map (
            O => \N__9209\,
            I => \receive_module.rx_counter.n3352\
        );

    \I__932\ : InMux
    port map (
            O => \N__9206\,
            I => \receive_module.rx_counter.n3353\
        );

    \I__931\ : InMux
    port map (
            O => \N__9203\,
            I => \receive_module.rx_counter.n3354\
        );

    \I__930\ : InMux
    port map (
            O => \N__9200\,
            I => \receive_module.rx_counter.n3355\
        );

    \I__929\ : InMux
    port map (
            O => \N__9197\,
            I => \bfn_11_10_0_\
        );

    \I__928\ : CEMux
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__9191\,
            I => \N__9187\
        );

    \I__926\ : CEMux
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__925\ : Sp12to4
    port map (
            O => \N__9187\,
            I => \N__9179\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__9184\,
            I => \N__9179\
        );

    \I__923\ : Odrv12
    port map (
            O => \N__9179\,
            I => n2057
        );

    \I__922\ : InMux
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__9170\,
            I => \transmit_module.Y_DELTA_PATTERN_51\
        );

    \I__919\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__9161\,
            I => \transmit_module.Y_DELTA_PATTERN_63\
        );

    \I__916\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__9155\,
            I => \transmit_module.Y_DELTA_PATTERN_62\
        );

    \I__914\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__9149\,
            I => \transmit_module.Y_DELTA_PATTERN_74\
        );

    \I__912\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9143\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__9143\,
            I => \transmit_module.Y_DELTA_PATTERN_50\
        );

    \I__910\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__9137\,
            I => \transmit_module.Y_DELTA_PATTERN_49\
        );

    \I__908\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__9131\,
            I => \transmit_module.Y_DELTA_PATTERN_65\
        );

    \I__906\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__9122\,
            I => \transmit_module.Y_DELTA_PATTERN_64\
        );

    \I__903\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__9116\,
            I => \transmit_module.X_DELTA_PATTERN_12\
        );

    \I__901\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__9110\,
            I => \transmit_module.X_DELTA_PATTERN_13\
        );

    \I__899\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__9104\,
            I => \old_HS\
        );

    \I__897\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__9098\,
            I => \transmit_module.Y_DELTA_PATTERN_79\
        );

    \I__895\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__9089\,
            I => \transmit_module.Y_DELTA_PATTERN_48\
        );

    \I__892\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__9083\,
            I => \transmit_module.Y_DELTA_PATTERN_47\
        );

    \I__890\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__9077\,
            I => \transmit_module.Y_DELTA_PATTERN_67\
        );

    \I__888\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__9071\,
            I => \transmit_module.Y_DELTA_PATTERN_82\
        );

    \I__886\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__9065\,
            I => \transmit_module.Y_DELTA_PATTERN_44\
        );

    \I__884\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__9059\,
            I => \transmit_module.Y_DELTA_PATTERN_43\
        );

    \I__882\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__9053\,
            I => \transmit_module.Y_DELTA_PATTERN_81\
        );

    \I__880\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__9047\,
            I => \transmit_module.Y_DELTA_PATTERN_80\
        );

    \I__878\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__9041\,
            I => \transmit_module.Y_DELTA_PATTERN_66\
        );

    \I__876\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__9032\,
            I => \transmit_module.Y_DELTA_PATTERN_76\
        );

    \I__873\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__9026\,
            I => \transmit_module.Y_DELTA_PATTERN_75\
        );

    \I__871\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9020\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__9020\,
            I => \transmit_module.Y_DELTA_PATTERN_45\
        );

    \I__869\ : InMux
    port map (
            O => \N__9017\,
            I => \N__9014\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__9014\,
            I => \transmit_module.Y_DELTA_PATTERN_77\
        );

    \I__867\ : InMux
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__9008\,
            I => \transmit_module.Y_DELTA_PATTERN_3\
        );

    \I__865\ : InMux
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__9002\,
            I => \transmit_module.Y_DELTA_PATTERN_2\
        );

    \I__863\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__8996\,
            I => \transmit_module.Y_DELTA_PATTERN_46\
        );

    \I__861\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8990\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__8990\,
            I => \transmit_module.Y_DELTA_PATTERN_78\
        );

    \I__859\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8984\,
            I => \transmit_module.Y_DELTA_PATTERN_68\
        );

    \I__857\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__8978\,
            I => \transmit_module.Y_DELTA_PATTERN_6\
        );

    \I__855\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__8972\,
            I => \transmit_module.Y_DELTA_PATTERN_20\
        );

    \I__853\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8966\,
            I => \transmit_module.Y_DELTA_PATTERN_21\
        );

    \I__851\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8960\,
            I => \N__8957\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__8957\,
            I => \transmit_module.Y_DELTA_PATTERN_23\
        );

    \I__848\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8951\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__8951\,
            I => \transmit_module.Y_DELTA_PATTERN_22\
        );

    \I__846\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__8942\,
            I => \transmit_module.Y_DELTA_PATTERN_5\
        );

    \I__843\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__8936\,
            I => \transmit_module.Y_DELTA_PATTERN_1\
        );

    \I__841\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__8930\,
            I => \transmit_module.Y_DELTA_PATTERN_4\
        );

    \I__839\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__8924\,
            I => \transmit_module.Y_DELTA_PATTERN_69\
        );

    \I__837\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8918\,
            I => \N__8915\
        );

    \I__835\ : Span4Mux_h
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__8912\,
            I => \transmit_module.Y_DELTA_PATTERN_56\
        );

    \I__833\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8906\,
            I => \transmit_module.Y_DELTA_PATTERN_58\
        );

    \I__831\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8900\,
            I => \transmit_module.Y_DELTA_PATTERN_57\
        );

    \I__829\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__8894\,
            I => \transmit_module.Y_DELTA_PATTERN_61\
        );

    \I__827\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8888\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__8888\,
            I => \N__8885\
        );

    \I__825\ : Span4Mux_v
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__824\ : Odrv4
    port map (
            O => \N__8882\,
            I => \line_buffer.n639\
        );

    \I__823\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8876\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__821\ : Odrv4
    port map (
            O => \N__8873\,
            I => \line_buffer.n631\
        );

    \I__820\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8867\,
            I => \transmit_module.X_DELTA_PATTERN_11\
        );

    \I__818\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8861\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__8861\,
            I => \N__8858\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__8858\,
            I => \transmit_module.X_DELTA_PATTERN_10\
        );

    \I__815\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8852\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8852\,
            I => \transmit_module.Y_DELTA_PATTERN_24\
        );

    \I__813\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__8846\,
            I => \transmit_module.Y_DELTA_PATTERN_71\
        );

    \I__811\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__8840\,
            I => \transmit_module.Y_DELTA_PATTERN_70\
        );

    \I__809\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__8834\,
            I => \transmit_module.Y_DELTA_PATTERN_60\
        );

    \I__807\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8828\,
            I => \transmit_module.Y_DELTA_PATTERN_59\
        );

    \I__805\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8822\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8822\,
            I => \transmit_module.Y_DELTA_PATTERN_42\
        );

    \I__803\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8816\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__8816\,
            I => \transmit_module.Y_DELTA_PATTERN_41\
        );

    \I__801\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__8810\,
            I => \transmit_module.Y_DELTA_PATTERN_14\
        );

    \I__799\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__8804\,
            I => \transmit_module.Y_DELTA_PATTERN_15\
        );

    \I__797\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8798\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__8798\,
            I => \transmit_module.Y_DELTA_PATTERN_16\
        );

    \I__795\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__8792\,
            I => \transmit_module.Y_DELTA_PATTERN_17\
        );

    \I__793\ : InMux
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__8786\,
            I => \transmit_module.Y_DELTA_PATTERN_19\
        );

    \I__791\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__8780\,
            I => \transmit_module.Y_DELTA_PATTERN_18\
        );

    \I__789\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__787\ : Span4Mux_s2_v
    port map (
            O => \N__8771\,
            I => \N__8767\
        );

    \I__786\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8764\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__8767\,
            I => \N__8759\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__8764\,
            I => \N__8759\
        );

    \I__783\ : Span4Mux_v
    port map (
            O => \N__8759\,
            I => \N__8755\
        );

    \I__782\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8752\
        );

    \I__781\ : Span4Mux_v
    port map (
            O => \N__8755\,
            I => \N__8746\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__8752\,
            I => \N__8746\
        );

    \I__779\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8743\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__8746\,
            I => \N__8738\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__8743\,
            I => \N__8738\
        );

    \I__776\ : Span4Mux_v
    port map (
            O => \N__8738\,
            I => \N__8733\
        );

    \I__775\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8730\
        );

    \I__774\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8727\
        );

    \I__773\ : Span4Mux_v
    port map (
            O => \N__8733\,
            I => \N__8722\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8730\,
            I => \N__8722\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__8727\,
            I => \N__8719\
        );

    \I__770\ : Span4Mux_h
    port map (
            O => \N__8722\,
            I => \N__8715\
        );

    \I__769\ : Span4Mux_h
    port map (
            O => \N__8719\,
            I => \N__8712\
        );

    \I__768\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8709\
        );

    \I__767\ : Span4Mux_h
    port map (
            O => \N__8715\,
            I => \N__8706\
        );

    \I__766\ : Span4Mux_v
    port map (
            O => \N__8712\,
            I => \N__8702\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__8709\,
            I => \N__8699\
        );

    \I__764\ : Span4Mux_h
    port map (
            O => \N__8706\,
            I => \N__8696\
        );

    \I__763\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8693\
        );

    \I__762\ : Span4Mux_v
    port map (
            O => \N__8702\,
            I => \N__8688\
        );

    \I__761\ : Span4Mux_h
    port map (
            O => \N__8699\,
            I => \N__8688\
        );

    \I__760\ : Span4Mux_h
    port map (
            O => \N__8696\,
            I => \N__8683\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__8693\,
            I => \N__8683\
        );

    \I__758\ : Span4Mux_v
    port map (
            O => \N__8688\,
            I => \N__8680\
        );

    \I__757\ : Span4Mux_h
    port map (
            O => \N__8683\,
            I => \N__8677\
        );

    \I__756\ : Span4Mux_v
    port map (
            O => \N__8680\,
            I => \N__8674\
        );

    \I__755\ : Span4Mux_v
    port map (
            O => \N__8677\,
            I => \N__8671\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__8674\,
            I => \TVP_VIDEO_c_2\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__8671\,
            I => \TVP_VIDEO_c_2\
        );

    \I__752\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8663\,
            I => \transmit_module.Y_DELTA_PATTERN_55\
        );

    \I__750\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__8657\,
            I => \transmit_module.Y_DELTA_PATTERN_54\
        );

    \I__748\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__8651\,
            I => \transmit_module.Y_DELTA_PATTERN_53\
        );

    \I__746\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8645\,
            I => \transmit_module.Y_DELTA_PATTERN_52\
        );

    \I__744\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__8639\,
            I => \N__8633\
        );

    \I__742\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8630\
        );

    \I__741\ : InMux
    port map (
            O => \N__8637\,
            I => \N__8627\
        );

    \I__740\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8623\
        );

    \I__739\ : Span4Mux_v
    port map (
            O => \N__8633\,
            I => \N__8616\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__8630\,
            I => \N__8616\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8616\
        );

    \I__736\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8613\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__8623\,
            I => \N__8609\
        );

    \I__734\ : Span4Mux_v
    port map (
            O => \N__8616\,
            I => \N__8604\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8613\,
            I => \N__8604\
        );

    \I__732\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8601\
        );

    \I__731\ : Span4Mux_v
    port map (
            O => \N__8609\,
            I => \N__8596\
        );

    \I__730\ : Span4Mux_v
    port map (
            O => \N__8604\,
            I => \N__8591\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__8601\,
            I => \N__8591\
        );

    \I__728\ : InMux
    port map (
            O => \N__8600\,
            I => \N__8588\
        );

    \I__727\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8585\
        );

    \I__726\ : Span4Mux_v
    port map (
            O => \N__8596\,
            I => \N__8582\
        );

    \I__725\ : Span4Mux_v
    port map (
            O => \N__8591\,
            I => \N__8579\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__8588\,
            I => \N__8576\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__8585\,
            I => \N__8573\
        );

    \I__722\ : Sp12to4
    port map (
            O => \N__8582\,
            I => \N__8570\
        );

    \I__721\ : Span4Mux_v
    port map (
            O => \N__8579\,
            I => \N__8567\
        );

    \I__720\ : Span4Mux_h
    port map (
            O => \N__8576\,
            I => \N__8564\
        );

    \I__719\ : Span4Mux_h
    port map (
            O => \N__8573\,
            I => \N__8561\
        );

    \I__718\ : Span12Mux_h
    port map (
            O => \N__8570\,
            I => \N__8558\
        );

    \I__717\ : Sp12to4
    port map (
            O => \N__8567\,
            I => \N__8555\
        );

    \I__716\ : IoSpan4Mux
    port map (
            O => \N__8564\,
            I => \N__8552\
        );

    \I__715\ : Span4Mux_h
    port map (
            O => \N__8561\,
            I => \N__8549\
        );

    \I__714\ : Span12Mux_v
    port map (
            O => \N__8558\,
            I => \N__8546\
        );

    \I__713\ : Span12Mux_h
    port map (
            O => \N__8555\,
            I => \N__8543\
        );

    \I__712\ : IoSpan4Mux
    port map (
            O => \N__8552\,
            I => \N__8540\
        );

    \I__711\ : Span4Mux_h
    port map (
            O => \N__8549\,
            I => \N__8537\
        );

    \I__710\ : Odrv12
    port map (
            O => \N__8546\,
            I => \TVP_VIDEO_c_8\
        );

    \I__709\ : Odrv12
    port map (
            O => \N__8543\,
            I => \TVP_VIDEO_c_8\
        );

    \I__708\ : Odrv4
    port map (
            O => \N__8540\,
            I => \TVP_VIDEO_c_8\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__8537\,
            I => \TVP_VIDEO_c_8\
        );

    \I__706\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8524\
        );

    \I__705\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8521\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__8524\,
            I => \N__8515\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8515\
        );

    \I__702\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8512\
        );

    \I__701\ : Span4Mux_v
    port map (
            O => \N__8515\,
            I => \N__8507\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__8512\,
            I => \N__8507\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__8507\,
            I => \N__8503\
        );

    \I__698\ : InMux
    port map (
            O => \N__8506\,
            I => \N__8500\
        );

    \I__697\ : Span4Mux_v
    port map (
            O => \N__8503\,
            I => \N__8494\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__8500\,
            I => \N__8494\
        );

    \I__695\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8490\
        );

    \I__694\ : Span4Mux_h
    port map (
            O => \N__8494\,
            I => \N__8487\
        );

    \I__693\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8484\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__8490\,
            I => \N__8481\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__8487\,
            I => \N__8478\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8475\
        );

    \I__689\ : Span12Mux_s11_h
    port map (
            O => \N__8481\,
            I => \N__8471\
        );

    \I__688\ : Sp12to4
    port map (
            O => \N__8478\,
            I => \N__8468\
        );

    \I__687\ : Span12Mux_s8_h
    port map (
            O => \N__8475\,
            I => \N__8465\
        );

    \I__686\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8462\
        );

    \I__685\ : Span12Mux_v
    port map (
            O => \N__8471\,
            I => \N__8459\
        );

    \I__684\ : Span12Mux_v
    port map (
            O => \N__8468\,
            I => \N__8456\
        );

    \I__683\ : Span12Mux_v
    port map (
            O => \N__8465\,
            I => \N__8453\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8450\
        );

    \I__681\ : Span12Mux_h
    port map (
            O => \N__8459\,
            I => \N__8446\
        );

    \I__680\ : Span12Mux_h
    port map (
            O => \N__8456\,
            I => \N__8441\
        );

    \I__679\ : Span12Mux_v
    port map (
            O => \N__8453\,
            I => \N__8441\
        );

    \I__678\ : Span4Mux_h
    port map (
            O => \N__8450\,
            I => \N__8438\
        );

    \I__677\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8435\
        );

    \I__676\ : Odrv12
    port map (
            O => \N__8446\,
            I => \TVP_VIDEO_c_9\
        );

    \I__675\ : Odrv12
    port map (
            O => \N__8441\,
            I => \TVP_VIDEO_c_9\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__8438\,
            I => \TVP_VIDEO_c_9\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__8435\,
            I => \TVP_VIDEO_c_9\
        );

    \I__672\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8423\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__8423\,
            I => \N__8417\
        );

    \I__670\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8414\
        );

    \I__669\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8411\
        );

    \I__668\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8408\
        );

    \I__667\ : Span4Mux_h
    port map (
            O => \N__8417\,
            I => \N__8405\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8401\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8398\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8394\
        );

    \I__663\ : Span4Mux_h
    port map (
            O => \N__8405\,
            I => \N__8391\
        );

    \I__662\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8388\
        );

    \I__661\ : Span4Mux_h
    port map (
            O => \N__8401\,
            I => \N__8385\
        );

    \I__660\ : Span4Mux_v
    port map (
            O => \N__8398\,
            I => \N__8382\
        );

    \I__659\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8377\
        );

    \I__658\ : Span12Mux_h
    port map (
            O => \N__8394\,
            I => \N__8374\
        );

    \I__657\ : Sp12to4
    port map (
            O => \N__8391\,
            I => \N__8371\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__8388\,
            I => \N__8368\
        );

    \I__655\ : Span4Mux_h
    port map (
            O => \N__8385\,
            I => \N__8365\
        );

    \I__654\ : Span4Mux_v
    port map (
            O => \N__8382\,
            I => \N__8362\
        );

    \I__653\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8359\
        );

    \I__652\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8356\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__8377\,
            I => \N__8353\
        );

    \I__650\ : Span12Mux_v
    port map (
            O => \N__8374\,
            I => \N__8350\
        );

    \I__649\ : Span12Mux_v
    port map (
            O => \N__8371\,
            I => \N__8343\
        );

    \I__648\ : Span12Mux_h
    port map (
            O => \N__8368\,
            I => \N__8343\
        );

    \I__647\ : Sp12to4
    port map (
            O => \N__8365\,
            I => \N__8343\
        );

    \I__646\ : Sp12to4
    port map (
            O => \N__8362\,
            I => \N__8338\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8338\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__8356\,
            I => \N__8335\
        );

    \I__643\ : Span4Mux_h
    port map (
            O => \N__8353\,
            I => \N__8332\
        );

    \I__642\ : Span12Mux_v
    port map (
            O => \N__8350\,
            I => \N__8329\
        );

    \I__641\ : Span12Mux_v
    port map (
            O => \N__8343\,
            I => \N__8322\
        );

    \I__640\ : Span12Mux_h
    port map (
            O => \N__8338\,
            I => \N__8322\
        );

    \I__639\ : Span12Mux_h
    port map (
            O => \N__8335\,
            I => \N__8322\
        );

    \I__638\ : Span4Mux_h
    port map (
            O => \N__8332\,
            I => \N__8319\
        );

    \I__637\ : Odrv12
    port map (
            O => \N__8329\,
            I => \TVP_VIDEO_c_7\
        );

    \I__636\ : Odrv12
    port map (
            O => \N__8322\,
            I => \TVP_VIDEO_c_7\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__8319\,
            I => \TVP_VIDEO_c_7\
        );

    \I__634\ : InMux
    port map (
            O => \N__8312\,
            I => \N__8308\
        );

    \I__633\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8305\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__8308\,
            I => \N__8302\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__8305\,
            I => \N__8298\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__8302\,
            I => \N__8295\
        );

    \I__629\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8292\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__8298\,
            I => \N__8288\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__8295\,
            I => \N__8283\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__8292\,
            I => \N__8283\
        );

    \I__625\ : InMux
    port map (
            O => \N__8291\,
            I => \N__8280\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__8288\,
            I => \N__8277\
        );

    \I__623\ : Span4Mux_v
    port map (
            O => \N__8283\,
            I => \N__8271\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__8280\,
            I => \N__8271\
        );

    \I__621\ : Span4Mux_v
    port map (
            O => \N__8277\,
            I => \N__8267\
        );

    \I__620\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8264\
        );

    \I__619\ : Span4Mux_v
    port map (
            O => \N__8271\,
            I => \N__8260\
        );

    \I__618\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8257\
        );

    \I__617\ : Span4Mux_v
    port map (
            O => \N__8267\,
            I => \N__8252\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__8264\,
            I => \N__8252\
        );

    \I__615\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8249\
        );

    \I__614\ : Span4Mux_v
    port map (
            O => \N__8260\,
            I => \N__8244\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__8257\,
            I => \N__8244\
        );

    \I__612\ : Span4Mux_v
    port map (
            O => \N__8252\,
            I => \N__8239\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__8249\,
            I => \N__8239\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__8244\,
            I => \N__8235\
        );

    \I__609\ : Span4Mux_v
    port map (
            O => \N__8239\,
            I => \N__8232\
        );

    \I__608\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8229\
        );

    \I__607\ : Sp12to4
    port map (
            O => \N__8235\,
            I => \N__8226\
        );

    \I__606\ : Span4Mux_v
    port map (
            O => \N__8232\,
            I => \N__8221\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__8229\,
            I => \N__8221\
        );

    \I__604\ : Span12Mux_h
    port map (
            O => \N__8226\,
            I => \N__8218\
        );

    \I__603\ : Span4Mux_h
    port map (
            O => \N__8221\,
            I => \N__8215\
        );

    \I__602\ : Odrv12
    port map (
            O => \N__8218\,
            I => \TVP_VIDEO_c_6\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__8215\,
            I => \TVP_VIDEO_c_6\
        );

    \I__600\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8206\
        );

    \I__599\ : InMux
    port map (
            O => \N__8209\,
            I => \N__8203\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__8206\,
            I => \N__8200\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__8203\,
            I => \N__8196\
        );

    \I__596\ : Span4Mux_v
    port map (
            O => \N__8200\,
            I => \N__8193\
        );

    \I__595\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8190\
        );

    \I__594\ : Span4Mux_v
    port map (
            O => \N__8196\,
            I => \N__8187\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__8193\,
            I => \N__8181\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__8190\,
            I => \N__8181\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__8187\,
            I => \N__8177\
        );

    \I__590\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8174\
        );

    \I__589\ : Span4Mux_v
    port map (
            O => \N__8181\,
            I => \N__8171\
        );

    \I__588\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8168\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__8177\,
            I => \N__8162\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__8174\,
            I => \N__8162\
        );

    \I__585\ : Span4Mux_v
    port map (
            O => \N__8171\,
            I => \N__8156\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__8168\,
            I => \N__8156\
        );

    \I__583\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8153\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__8162\,
            I => \N__8150\
        );

    \I__581\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8147\
        );

    \I__580\ : Span4Mux_v
    port map (
            O => \N__8156\,
            I => \N__8142\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__8153\,
            I => \N__8142\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__8150\,
            I => \N__8137\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__8147\,
            I => \N__8137\
        );

    \I__576\ : Span4Mux_v
    port map (
            O => \N__8142\,
            I => \N__8133\
        );

    \I__575\ : Span4Mux_v
    port map (
            O => \N__8137\,
            I => \N__8130\
        );

    \I__574\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8127\
        );

    \I__573\ : Sp12to4
    port map (
            O => \N__8133\,
            I => \N__8124\
        );

    \I__572\ : Span4Mux_v
    port map (
            O => \N__8130\,
            I => \N__8119\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__8127\,
            I => \N__8119\
        );

    \I__570\ : Span12Mux_h
    port map (
            O => \N__8124\,
            I => \N__8116\
        );

    \I__569\ : Span4Mux_h
    port map (
            O => \N__8119\,
            I => \N__8113\
        );

    \I__568\ : Odrv12
    port map (
            O => \N__8116\,
            I => \TVP_VIDEO_c_5\
        );

    \I__567\ : Odrv4
    port map (
            O => \N__8113\,
            I => \TVP_VIDEO_c_5\
        );

    \I__566\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__564\ : Span4Mux_v
    port map (
            O => \N__8102\,
            I => \N__8096\
        );

    \I__563\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8093\
        );

    \I__562\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8089\
        );

    \I__561\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8085\
        );

    \I__560\ : Span4Mux_v
    port map (
            O => \N__8096\,
            I => \N__8080\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8080\
        );

    \I__558\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8077\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__8089\,
            I => \N__8074\
        );

    \I__556\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8071\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8068\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__8080\,
            I => \N__8063\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__8077\,
            I => \N__8063\
        );

    \I__552\ : Span4Mux_h
    port map (
            O => \N__8074\,
            I => \N__8060\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__8071\,
            I => \N__8057\
        );

    \I__550\ : Span4Mux_s1_v
    port map (
            O => \N__8068\,
            I => \N__8053\
        );

    \I__549\ : Span4Mux_v
    port map (
            O => \N__8063\,
            I => \N__8050\
        );

    \I__548\ : Span4Mux_h
    port map (
            O => \N__8060\,
            I => \N__8047\
        );

    \I__547\ : Span4Mux_h
    port map (
            O => \N__8057\,
            I => \N__8044\
        );

    \I__546\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8041\
        );

    \I__545\ : Sp12to4
    port map (
            O => \N__8053\,
            I => \N__8038\
        );

    \I__544\ : Span4Mux_h
    port map (
            O => \N__8050\,
            I => \N__8035\
        );

    \I__543\ : Span4Mux_h
    port map (
            O => \N__8047\,
            I => \N__8032\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__8044\,
            I => \N__8029\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__8041\,
            I => \N__8026\
        );

    \I__540\ : Span12Mux_s10_h
    port map (
            O => \N__8038\,
            I => \N__8022\
        );

    \I__539\ : Sp12to4
    port map (
            O => \N__8035\,
            I => \N__8019\
        );

    \I__538\ : Span4Mux_h
    port map (
            O => \N__8032\,
            I => \N__8012\
        );

    \I__537\ : Span4Mux_v
    port map (
            O => \N__8029\,
            I => \N__8012\
        );

    \I__536\ : Span4Mux_h
    port map (
            O => \N__8026\,
            I => \N__8012\
        );

    \I__535\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8009\
        );

    \I__534\ : Span12Mux_v
    port map (
            O => \N__8022\,
            I => \N__8006\
        );

    \I__533\ : Span12Mux_h
    port map (
            O => \N__8019\,
            I => \N__8003\
        );

    \I__532\ : Span4Mux_v
    port map (
            O => \N__8012\,
            I => \N__8000\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__8009\,
            I => \N__7997\
        );

    \I__530\ : Span12Mux_v
    port map (
            O => \N__8006\,
            I => \N__7994\
        );

    \I__529\ : Span12Mux_v
    port map (
            O => \N__8003\,
            I => \N__7991\
        );

    \I__528\ : Span4Mux_v
    port map (
            O => \N__8000\,
            I => \N__7988\
        );

    \I__527\ : Span4Mux_h
    port map (
            O => \N__7997\,
            I => \N__7985\
        );

    \I__526\ : Odrv12
    port map (
            O => \N__7994\,
            I => \TVP_VIDEO_c_4\
        );

    \I__525\ : Odrv12
    port map (
            O => \N__7991\,
            I => \TVP_VIDEO_c_4\
        );

    \I__524\ : Odrv4
    port map (
            O => \N__7988\,
            I => \TVP_VIDEO_c_4\
        );

    \I__523\ : Odrv4
    port map (
            O => \N__7985\,
            I => \TVP_VIDEO_c_4\
        );

    \I__522\ : InMux
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__520\ : Span4Mux_v
    port map (
            O => \N__7970\,
            I => \N__7966\
        );

    \I__519\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7963\
        );

    \I__518\ : Span4Mux_v
    port map (
            O => \N__7966\,
            I => \N__7957\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__7963\,
            I => \N__7957\
        );

    \I__516\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7954\
        );

    \I__515\ : Span4Mux_v
    port map (
            O => \N__7957\,
            I => \N__7951\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__7954\,
            I => \N__7948\
        );

    \I__513\ : Span4Mux_v
    port map (
            O => \N__7951\,
            I => \N__7942\
        );

    \I__512\ : Span4Mux_v
    port map (
            O => \N__7948\,
            I => \N__7942\
        );

    \I__511\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7939\
        );

    \I__510\ : Span4Mux_v
    port map (
            O => \N__7942\,
            I => \N__7933\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__7939\,
            I => \N__7933\
        );

    \I__508\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7930\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__7933\,
            I => \N__7924\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__7930\,
            I => \N__7924\
        );

    \I__505\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7921\
        );

    \I__504\ : Span4Mux_v
    port map (
            O => \N__7924\,
            I => \N__7916\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__7921\,
            I => \N__7913\
        );

    \I__502\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7910\
        );

    \I__501\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7907\
        );

    \I__500\ : Sp12to4
    port map (
            O => \N__7916\,
            I => \N__7904\
        );

    \I__499\ : Span4Mux_h
    port map (
            O => \N__7913\,
            I => \N__7901\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__7910\,
            I => \N__7898\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7895\
        );

    \I__496\ : Span12Mux_h
    port map (
            O => \N__7904\,
            I => \N__7892\
        );

    \I__495\ : Sp12to4
    port map (
            O => \N__7901\,
            I => \N__7889\
        );

    \I__494\ : Span4Mux_h
    port map (
            O => \N__7898\,
            I => \N__7886\
        );

    \I__493\ : Span12Mux_h
    port map (
            O => \N__7895\,
            I => \N__7883\
        );

    \I__492\ : Span12Mux_h
    port map (
            O => \N__7892\,
            I => \N__7876\
        );

    \I__491\ : Span12Mux_v
    port map (
            O => \N__7889\,
            I => \N__7876\
        );

    \I__490\ : Sp12to4
    port map (
            O => \N__7886\,
            I => \N__7876\
        );

    \I__489\ : Odrv12
    port map (
            O => \N__7883\,
            I => \TVP_VIDEO_c_3\
        );

    \I__488\ : Odrv12
    port map (
            O => \N__7876\,
            I => \TVP_VIDEO_c_3\
        );

    \INVADV_R__i1C\ : INV
    port map (
            O => \INVADV_R__i1C_net\,
            I => \N__22090\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3373\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3384\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.n3343\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3356\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3364\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.n3330\,
            carryinitout => \bfn_14_12_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i53_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8660\,
            lcout => \transmit_module.Y_DELTA_PATTERN_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22149\,
            ce => \N__17981\,
            sr => \N__20660\
        );

    \transmit_module.Y_DELTA_PATTERN_i55_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8921\,
            lcout => \transmit_module.Y_DELTA_PATTERN_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22149\,
            ce => \N__17981\,
            sr => \N__20660\
        );

    \transmit_module.Y_DELTA_PATTERN_i54_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8666\,
            lcout => \transmit_module.Y_DELTA_PATTERN_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22149\,
            ce => \N__17981\,
            sr => \N__20660\
        );

    \transmit_module.Y_DELTA_PATTERN_i52_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8654\,
            lcout => \transmit_module.Y_DELTA_PATTERN_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22149\,
            ce => \N__17981\,
            sr => \N__20660\
        );

    \transmit_module.Y_DELTA_PATTERN_i51_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8648\,
            lcout => \transmit_module.Y_DELTA_PATTERN_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22149\,
            ce => \N__17981\,
            sr => \N__20660\
        );

    \transmit_module.Y_DELTA_PATTERN_i63_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9128\,
            lcout => \transmit_module.Y_DELTA_PATTERN_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22070\,
            ce => \N__17980\,
            sr => \N__20690\
        );

    \transmit_module.X_DELTA_PATTERN_i9_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8864\,
            lcout => \transmit_module.X_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22087\,
            ce => \N__12880\,
            sr => \N__18724\
        );

    \transmit_module.Y_DELTA_PATTERN_i19_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8975\,
            lcout => \transmit_module.Y_DELTA_PATTERN_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21816\,
            ce => \N__18713\,
            sr => \N__20568\
        );

    \transmit_module.Y_DELTA_PATTERN_i13_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8813\,
            lcout => \transmit_module.Y_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21816\,
            ce => \N__18713\,
            sr => \N__20568\
        );

    \transmit_module.Y_DELTA_PATTERN_i14_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8807\,
            lcout => \transmit_module.Y_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21816\,
            ce => \N__18713\,
            sr => \N__20568\
        );

    \transmit_module.Y_DELTA_PATTERN_i15_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8801\,
            lcout => \transmit_module.Y_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21816\,
            ce => \N__18713\,
            sr => \N__20568\
        );

    \transmit_module.Y_DELTA_PATTERN_i16_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8795\,
            lcout => \transmit_module.Y_DELTA_PATTERN_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21816\,
            ce => \N__18713\,
            sr => \N__20568\
        );

    \transmit_module.Y_DELTA_PATTERN_i17_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8783\,
            lcout => \transmit_module.Y_DELTA_PATTERN_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21816\,
            ce => \N__18713\,
            sr => \N__20568\
        );

    \transmit_module.Y_DELTA_PATTERN_i18_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8789\,
            lcout => \transmit_module.Y_DELTA_PATTERN_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21816\,
            ce => \N__18713\,
            sr => \N__20568\
        );

    \transmit_module.Y_DELTA_PATTERN_i70_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8849\,
            lcout => \transmit_module.Y_DELTA_PATTERN_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22139\,
            ce => \N__17939\,
            sr => \N__20717\
        );

    \transmit_module.Y_DELTA_PATTERN_i71_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9383\,
            lcout => \transmit_module.Y_DELTA_PATTERN_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22139\,
            ce => \N__17939\,
            sr => \N__20717\
        );

    \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9062\,
            lcout => \transmit_module.Y_DELTA_PATTERN_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22139\,
            ce => \N__17939\,
            sr => \N__20717\
        );

    \transmit_module.Y_DELTA_PATTERN_i69_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8843\,
            lcout => \transmit_module.Y_DELTA_PATTERN_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22139\,
            ce => \N__17939\,
            sr => \N__20717\
        );

    \transmit_module.Y_DELTA_PATTERN_i59_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8837\,
            lcout => \transmit_module.Y_DELTA_PATTERN_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22086\,
            ce => \N__17984\,
            sr => \N__20713\
        );

    \transmit_module.Y_DELTA_PATTERN_i60_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8897\,
            lcout => \transmit_module.Y_DELTA_PATTERN_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22086\,
            ce => \N__17984\,
            sr => \N__20713\
        );

    \transmit_module.Y_DELTA_PATTERN_i58_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8831\,
            lcout => \transmit_module.Y_DELTA_PATTERN_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22086\,
            ce => \N__17984\,
            sr => \N__20713\
        );

    \transmit_module.Y_DELTA_PATTERN_i40_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8819\,
            lcout => \transmit_module.Y_DELTA_PATTERN_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22086\,
            ce => \N__17984\,
            sr => \N__20713\
        );

    \transmit_module.Y_DELTA_PATTERN_i41_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8825\,
            lcout => \transmit_module.Y_DELTA_PATTERN_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22086\,
            ce => \N__17984\,
            sr => \N__20713\
        );

    \transmit_module.Y_DELTA_PATTERN_i68_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8927\,
            lcout => \transmit_module.Y_DELTA_PATTERN_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22086\,
            ce => \N__17984\,
            sr => \N__20713\
        );

    \transmit_module.Y_DELTA_PATTERN_i56_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8903\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22088\,
            ce => \N__17983\,
            sr => \N__20691\
        );

    \transmit_module.Y_DELTA_PATTERN_i57_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8909\,
            lcout => \transmit_module.Y_DELTA_PATTERN_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22088\,
            ce => \N__17983\,
            sr => \N__20691\
        );

    \transmit_module.Y_DELTA_PATTERN_i61_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9158\,
            lcout => \transmit_module.Y_DELTA_PATTERN_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22088\,
            ce => \N__17983\,
            sr => \N__20691\
        );

    \transmit_module.Y_DELTA_PATTERN_i48_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9140\,
            lcout => \transmit_module.Y_DELTA_PATTERN_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22088\,
            ce => \N__17983\,
            sr => \N__20691\
        );

    \line_buffer.i2341_3_lut_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8891\,
            in1 => \N__8879\,
            in2 => \_gnd_net_\,
            in3 => \N__23108\,
            lcout => \line_buffer.n3703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i11_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9119\,
            lcout => \transmit_module.X_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => \N__12878\,
            sr => \N__18703\
        );

    \transmit_module.X_DELTA_PATTERN_i10_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8870\,
            lcout => \transmit_module.X_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => \N__12878\,
            sr => \N__18703\
        );

    \transmit_module.Y_DELTA_PATTERN_i23_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8855\,
            lcout => \transmit_module.Y_DELTA_PATTERN_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22145\,
            ce => \N__18730\,
            sr => \N__20698\
        );

    \transmit_module.Y_DELTA_PATTERN_i24_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9269\,
            lcout => \transmit_module.Y_DELTA_PATTERN_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22145\,
            ce => \N__18730\,
            sr => \N__20698\
        );

    \transmit_module.Y_DELTA_PATTERN_i6_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9263\,
            lcout => \transmit_module.Y_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22143\,
            ce => \N__18731\,
            sr => \N__20694\
        );

    \transmit_module.Y_DELTA_PATTERN_i5_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8981\,
            lcout => \transmit_module.Y_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22143\,
            ce => \N__18731\,
            sr => \N__20694\
        );

    \transmit_module.Y_DELTA_PATTERN_i20_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8969\,
            lcout => \transmit_module.Y_DELTA_PATTERN_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22104\,
            ce => \N__18726\,
            sr => \N__20697\
        );

    \transmit_module.Y_DELTA_PATTERN_i21_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8954\,
            lcout => \transmit_module.Y_DELTA_PATTERN_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22104\,
            ce => \N__18726\,
            sr => \N__20697\
        );

    \transmit_module.Y_DELTA_PATTERN_i22_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8963\,
            lcout => \transmit_module.Y_DELTA_PATTERN_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22104\,
            ce => \N__18726\,
            sr => \N__20697\
        );

    \transmit_module.Y_DELTA_PATTERN_i4_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8948\,
            lcout => \transmit_module.Y_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22142\,
            ce => \N__18725\,
            sr => \N__20695\
        );

    \transmit_module.Y_DELTA_PATTERN_i0_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8939\,
            lcout => \transmit_module.Y_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22142\,
            ce => \N__18725\,
            sr => \N__20695\
        );

    \transmit_module.Y_DELTA_PATTERN_i1_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22142\,
            ce => \N__18725\,
            sr => \N__20695\
        );

    \transmit_module.Y_DELTA_PATTERN_i3_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8933\,
            lcout => \transmit_module.Y_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22142\,
            ce => \N__18725\,
            sr => \N__20695\
        );

    \transmit_module.Y_DELTA_PATTERN_i44_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9023\,
            lcout => \transmit_module.Y_DELTA_PATTERN_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22103\,
            ce => \N__17962\,
            sr => \N__20517\
        );

    \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9017\,
            lcout => \transmit_module.Y_DELTA_PATTERN_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22103\,
            ce => \N__17962\,
            sr => \N__20517\
        );

    \transmit_module.Y_DELTA_PATTERN_i45_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8999\,
            lcout => \transmit_module.Y_DELTA_PATTERN_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22103\,
            ce => \N__17962\,
            sr => \N__20517\
        );

    \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8993\,
            lcout => \transmit_module.Y_DELTA_PATTERN_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22103\,
            ce => \N__17962\,
            sr => \N__20517\
        );

    \transmit_module.Y_DELTA_PATTERN_i2_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9011\,
            lcout => \transmit_module.Y_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22103\,
            ce => \N__17962\,
            sr => \N__20517\
        );

    \transmit_module.Y_DELTA_PATTERN_i46_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9086\,
            lcout => \transmit_module.Y_DELTA_PATTERN_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22103\,
            ce => \N__17962\,
            sr => \N__20517\
        );

    \transmit_module.Y_DELTA_PATTERN_i78_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9101\,
            lcout => \transmit_module.Y_DELTA_PATTERN_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22103\,
            ce => \N__17962\,
            sr => \N__20517\
        );

    \transmit_module.Y_DELTA_PATTERN_i67_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8987\,
            lcout => \transmit_module.Y_DELTA_PATTERN_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22138\,
            ce => \N__17970\,
            sr => \N__20649\
        );

    \transmit_module.Y_DELTA_PATTERN_i81_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9074\,
            lcout => \transmit_module.Y_DELTA_PATTERN_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22138\,
            ce => \N__17970\,
            sr => \N__20649\
        );

    \transmit_module.Y_DELTA_PATTERN_i79_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9050\,
            lcout => \transmit_module.Y_DELTA_PATTERN_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22138\,
            ce => \N__17970\,
            sr => \N__20649\
        );

    \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9095\,
            lcout => \transmit_module.Y_DELTA_PATTERN_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22138\,
            ce => \N__17970\,
            sr => \N__20649\
        );

    \transmit_module.Y_DELTA_PATTERN_i66_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9080\,
            lcout => \transmit_module.Y_DELTA_PATTERN_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22138\,
            ce => \N__17970\,
            sr => \N__20649\
        );

    \transmit_module.Y_DELTA_PATTERN_i82_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9323\,
            lcout => \transmit_module.Y_DELTA_PATTERN_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22138\,
            ce => \N__17970\,
            sr => \N__20649\
        );

    \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9068\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22138\,
            ce => \N__17970\,
            sr => \N__20649\
        );

    \transmit_module.Y_DELTA_PATTERN_i80_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9056\,
            lcout => \transmit_module.Y_DELTA_PATTERN_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22138\,
            ce => \N__17970\,
            sr => \N__20649\
        );

    \transmit_module.Y_DELTA_PATTERN_i74_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9029\,
            lcout => \transmit_module.Y_DELTA_PATTERN_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22099\,
            ce => \N__17969\,
            sr => \N__20518\
        );

    \transmit_module.Y_DELTA_PATTERN_i65_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9044\,
            lcout => \transmit_module.Y_DELTA_PATTERN_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22099\,
            ce => \N__17969\,
            sr => \N__20518\
        );

    \transmit_module.Y_DELTA_PATTERN_i75_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9038\,
            lcout => \transmit_module.Y_DELTA_PATTERN_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22099\,
            ce => \N__17969\,
            sr => \N__20518\
        );

    \transmit_module.Y_DELTA_PATTERN_i50_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9176\,
            lcout => \transmit_module.Y_DELTA_PATTERN_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22118\,
            ce => \N__17982\,
            sr => \N__20656\
        );

    \transmit_module.Y_DELTA_PATTERN_i62_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9167\,
            lcout => \transmit_module.Y_DELTA_PATTERN_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22118\,
            ce => \N__17982\,
            sr => \N__20656\
        );

    \transmit_module.Y_DELTA_PATTERN_i73_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9152\,
            lcout => \transmit_module.Y_DELTA_PATTERN_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22118\,
            ce => \N__17982\,
            sr => \N__20656\
        );

    \transmit_module.Y_DELTA_PATTERN_i49_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9146\,
            lcout => \transmit_module.Y_DELTA_PATTERN_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22118\,
            ce => \N__17982\,
            sr => \N__20656\
        );

    \transmit_module.Y_DELTA_PATTERN_i64_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9134\,
            lcout => \transmit_module.Y_DELTA_PATTERN_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22118\,
            ce => \N__17982\,
            sr => \N__20656\
        );

    \transmit_module.X_DELTA_PATTERN_i12_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9113\,
            lcout => \transmit_module.X_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21983\,
            ce => \N__12881\,
            sr => \N__18701\
        );

    \transmit_module.X_DELTA_PATTERN_i13_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9593\,
            lcout => \transmit_module.X_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21983\,
            ce => \N__12881\,
            sr => \N__18701\
        );

    \receive_module.rx_counter.old_HS_50_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19913\,
            lcout => \old_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i272_3_lut_3_lut_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__19912\,
            in1 => \N__9107\,
            in2 => \_gnd_net_\,
            in3 => \N__17770\,
            lcout => n2057,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.Y__i0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9968\,
            in2 => \_gnd_net_\,
            in3 => \N__9221\,
            lcout => \receive_module.rx_counter.Y_0\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \receive_module.rx_counter.n3349\,
            clk => \N__21012\,
            ce => \N__9190\,
            sr => \N__17697\
        );

    \receive_module.rx_counter.Y__i1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11074\,
            in2 => \_gnd_net_\,
            in3 => \N__9218\,
            lcout => \receive_module.rx_counter.Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3349\,
            carryout => \receive_module.rx_counter.n3350\,
            clk => \N__21012\,
            ce => \N__9190\,
            sr => \N__17697\
        );

    \receive_module.rx_counter.Y__i2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9940\,
            in2 => \_gnd_net_\,
            in3 => \N__9215\,
            lcout => \receive_module.rx_counter.Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3350\,
            carryout => \receive_module.rx_counter.n3351\,
            clk => \N__21012\,
            ce => \N__9190\,
            sr => \N__17697\
        );

    \receive_module.rx_counter.Y__i3_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11104\,
            in2 => \_gnd_net_\,
            in3 => \N__9212\,
            lcout => \receive_module.rx_counter.Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3351\,
            carryout => \receive_module.rx_counter.n3352\,
            clk => \N__21012\,
            ce => \N__9190\,
            sr => \N__17697\
        );

    \receive_module.rx_counter.Y__i4_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11134\,
            in2 => \_gnd_net_\,
            in3 => \N__9209\,
            lcout => \receive_module.rx_counter.Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3352\,
            carryout => \receive_module.rx_counter.n3353\,
            clk => \N__21012\,
            ce => \N__9190\,
            sr => \N__17697\
        );

    \receive_module.rx_counter.Y__i5_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9539\,
            in2 => \_gnd_net_\,
            in3 => \N__9206\,
            lcout => \receive_module.rx_counter.Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3353\,
            carryout => \receive_module.rx_counter.n3354\,
            clk => \N__21012\,
            ce => \N__9190\,
            sr => \N__17697\
        );

    \receive_module.rx_counter.Y__i6_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9554\,
            in2 => \_gnd_net_\,
            in3 => \N__9203\,
            lcout => \receive_module.rx_counter.Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3354\,
            carryout => \receive_module.rx_counter.n3355\,
            clk => \N__21012\,
            ce => \N__9190\,
            sr => \N__17697\
        );

    \receive_module.rx_counter.Y__i7_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9992\,
            in2 => \_gnd_net_\,
            in3 => \N__9200\,
            lcout => \receive_module.rx_counter.Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3355\,
            carryout => \receive_module.rx_counter.n3356\,
            clk => \N__21012\,
            ce => \N__9190\,
            sr => \N__17697\
        );

    \receive_module.rx_counter.Y__i8_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10009\,
            in2 => \_gnd_net_\,
            in3 => \N__9197\,
            lcout => \receive_module.rx_counter.Y_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21017\,
            ce => \N__9194\,
            sr => \N__17675\
        );

    \transmit_module.Y_DELTA_PATTERN_i26_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9257\,
            lcout => \transmit_module.Y_DELTA_PATTERN_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22117\,
            ce => \N__18712\,
            sr => \N__20692\
        );

    \transmit_module.Y_DELTA_PATTERN_i25_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9275\,
            lcout => \transmit_module.Y_DELTA_PATTERN_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22117\,
            ce => \N__18712\,
            sr => \N__20692\
        );

    \transmit_module.Y_DELTA_PATTERN_i7_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9227\,
            lcout => \transmit_module.Y_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22117\,
            ce => \N__18712\,
            sr => \N__20692\
        );

    \transmit_module.Y_DELTA_PATTERN_i10_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9329\,
            lcout => \transmit_module.Y_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22072\,
            ce => \N__18720\,
            sr => \N__20696\
        );

    \transmit_module.Y_DELTA_PATTERN_i27_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9416\,
            lcout => \transmit_module.Y_DELTA_PATTERN_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22072\,
            ce => \N__18720\,
            sr => \N__20696\
        );

    \transmit_module.Y_DELTA_PATTERN_i99_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19188\,
            lcout => \transmit_module.Y_DELTA_PATTERN_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22072\,
            ce => \N__18720\,
            sr => \N__20696\
        );

    \transmit_module.Y_DELTA_PATTERN_i9_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9251\,
            lcout => \transmit_module.Y_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22072\,
            ce => \N__18720\,
            sr => \N__20696\
        );

    \transmit_module.Y_DELTA_PATTERN_i12_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9245\,
            lcout => \transmit_module.Y_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22072\,
            ce => \N__18720\,
            sr => \N__20696\
        );

    \transmit_module.Y_DELTA_PATTERN_i8_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9233\,
            lcout => \transmit_module.Y_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22072\,
            ce => \N__18720\,
            sr => \N__20696\
        );

    \transmit_module.Y_DELTA_PATTERN_i11_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9335\,
            lcout => \transmit_module.Y_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22072\,
            ce => \N__18720\,
            sr => \N__20696\
        );

    \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10130\,
            lcout => \transmit_module.Y_DELTA_PATTERN_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22141\,
            ce => \N__10079\,
            sr => \N__20693\
        );

    \transmit_module.Y_DELTA_PATTERN_i83_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9311\,
            lcout => \transmit_module.Y_DELTA_PATTERN_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22141\,
            ce => \N__10079\,
            sr => \N__20693\
        );

    \transmit_module.Y_DELTA_PATTERN_i84_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9287\,
            lcout => \transmit_module.Y_DELTA_PATTERN_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22141\,
            ce => \N__10079\,
            sr => \N__20693\
        );

    \transmit_module.Y_DELTA_PATTERN_i93_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9299\,
            lcout => \transmit_module.Y_DELTA_PATTERN_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22141\,
            ce => \N__10079\,
            sr => \N__20693\
        );

    \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9305\,
            lcout => \transmit_module.Y_DELTA_PATTERN_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22141\,
            ce => \N__10079\,
            sr => \N__20693\
        );

    \transmit_module.Y_DELTA_PATTERN_i92_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9293\,
            lcout => \transmit_module.Y_DELTA_PATTERN_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22071\,
            ce => \N__10067\,
            sr => \N__20516\
        );

    \transmit_module.Y_DELTA_PATTERN_i90_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9365\,
            lcout => \transmit_module.Y_DELTA_PATTERN_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22071\,
            ce => \N__10067\,
            sr => \N__20516\
        );

    \transmit_module.Y_DELTA_PATTERN_i85_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9281\,
            lcout => \transmit_module.Y_DELTA_PATTERN_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22071\,
            ce => \N__10067\,
            sr => \N__20516\
        );

    \transmit_module.Y_DELTA_PATTERN_i86_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10031\,
            lcout => \transmit_module.Y_DELTA_PATTERN_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22071\,
            ce => \N__10067\,
            sr => \N__20516\
        );

    \transmit_module.Y_DELTA_PATTERN_i91_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9371\,
            lcout => \transmit_module.Y_DELTA_PATTERN_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22071\,
            ce => \N__10067\,
            sr => \N__20516\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i1_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10100\,
            in2 => \_gnd_net_\,
            in3 => \N__9359\,
            lcout => \transmit_module.video_signal_controller.VGA_X_0\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \transmit_module.video_signal_controller.n3377\,
            clk => \N__22095\,
            ce => 'H',
            sr => \N__17644\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i2_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10124\,
            in2 => \_gnd_net_\,
            in3 => \N__9356\,
            lcout => \transmit_module.video_signal_controller.VGA_X_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3377\,
            carryout => \transmit_module.video_signal_controller.n3378\,
            clk => \N__22095\,
            ce => 'H',
            sr => \N__17644\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i3_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10112\,
            in2 => \_gnd_net_\,
            in3 => \N__9353\,
            lcout => \transmit_module.video_signal_controller.VGA_X_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3378\,
            carryout => \transmit_module.video_signal_controller.n3379\,
            clk => \N__22095\,
            ce => 'H',
            sr => \N__17644\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i4_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11199\,
            in2 => \_gnd_net_\,
            in3 => \N__9350\,
            lcout => \transmit_module.video_signal_controller.VGA_X_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3379\,
            carryout => \transmit_module.video_signal_controller.n3380\,
            clk => \N__22095\,
            ce => 'H',
            sr => \N__17644\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i5_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11230\,
            in2 => \_gnd_net_\,
            in3 => \N__9347\,
            lcout => \transmit_module.video_signal_controller.VGA_X_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3380\,
            carryout => \transmit_module.video_signal_controller.n3381\,
            clk => \N__22095\,
            ce => 'H',
            sr => \N__17644\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i6_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11173\,
            in2 => \_gnd_net_\,
            in3 => \N__9344\,
            lcout => \transmit_module.video_signal_controller.VGA_X_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3381\,
            carryout => \transmit_module.video_signal_controller.n3382\,
            clk => \N__22095\,
            ce => 'H',
            sr => \N__17644\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i7_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10162\,
            in2 => \_gnd_net_\,
            in3 => \N__9341\,
            lcout => \transmit_module.video_signal_controller.VGA_X_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3382\,
            carryout => \transmit_module.video_signal_controller.n3383\,
            clk => \N__22095\,
            ce => 'H',
            sr => \N__17644\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i8_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10183\,
            in2 => \_gnd_net_\,
            in3 => \N__9338\,
            lcout => \transmit_module.video_signal_controller.VGA_X_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3383\,
            carryout => \transmit_module.video_signal_controller.n3384\,
            clk => \N__22095\,
            ce => 'H',
            sr => \N__17644\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i9_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12016\,
            in2 => \_gnd_net_\,
            in3 => \N__9425\,
            lcout => \transmit_module.video_signal_controller.VGA_X_8\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \transmit_module.video_signal_controller.n3385\,
            clk => \N__21949\,
            ce => 'H',
            sr => \N__17645\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i10_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10698\,
            in2 => \_gnd_net_\,
            in3 => \N__9422\,
            lcout => \transmit_module.video_signal_controller.VGA_X_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3385\,
            carryout => \transmit_module.video_signal_controller.n3386\,
            clk => \N__21949\,
            ce => 'H',
            sr => \N__17645\
        );

    \transmit_module.video_signal_controller.VGA_X_266_267__i11_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10732\,
            in2 => \_gnd_net_\,
            in3 => \N__9419\,
            lcout => \transmit_module.video_signal_controller.VGA_X_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21949\,
            ce => 'H',
            sr => \N__17645\
        );

    \transmit_module.Y_DELTA_PATTERN_i28_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9407\,
            lcout => \transmit_module.Y_DELTA_PATTERN_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__18707\,
            sr => \N__20630\
        );

    \transmit_module.Y_DELTA_PATTERN_i29_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9401\,
            lcout => \transmit_module.Y_DELTA_PATTERN_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__18707\,
            sr => \N__20630\
        );

    \transmit_module.Y_DELTA_PATTERN_i30_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9395\,
            lcout => \transmit_module.Y_DELTA_PATTERN_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__18707\,
            sr => \N__20630\
        );

    \transmit_module.Y_DELTA_PATTERN_i31_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18743\,
            lcout => \transmit_module.Y_DELTA_PATTERN_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__18707\,
            sr => \N__20630\
        );

    \transmit_module.Y_DELTA_PATTERN_i72_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9389\,
            lcout => \transmit_module.Y_DELTA_PATTERN_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21946\,
            ce => \N__18707\,
            sr => \N__20630\
        );

    \transmit_module.i2_4_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__16575\,
            in1 => \N__19708\,
            in2 => \N__20684\,
            in3 => \N__19605\,
            lcout => \transmit_module.n2099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1681_4_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__10660\,
            in1 => \N__10667\,
            in2 => \N__20712\,
            in3 => \N__20252\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i15_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12931\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22042\,
            ce => \N__12867\,
            sr => \N__18694\
        );

    \transmit_module.X_DELTA_PATTERN_i14_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9599\,
            lcout => \transmit_module.X_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22042\,
            ce => \N__12867\,
            sr => \N__18694\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2435_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__9587\,
            in1 => \N__22929\,
            in2 => \N__9572\,
            in3 => \N__23132\,
            lcout => \line_buffer.n3785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_rep_25_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9537\,
            in2 => \_gnd_net_\,
            in3 => \N__9552\,
            lcout => \receive_module.rx_counter.n3861\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_4_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9553\,
            in1 => \N__9991\,
            in2 => \N__10010\,
            in3 => \N__9538\,
            lcout => \receive_module.rx_counter.n3619\,
            ltout => \receive_module.rx_counter.n3619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i4_4_lut_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__11070\,
            in1 => \N__11100\,
            in2 => \N__9521\,
            in3 => \N__11130\,
            lcout => \receive_module.rx_counter.n10_adj_570\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15912\,
            in1 => \N__15752\,
            in2 => \N__15860\,
            in3 => \N__11302\,
            lcout => \line_buffer.n642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_9_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__11303\,
            in1 => \N__15913\,
            in2 => \N__15765\,
            in3 => \N__15859\,
            lcout => \line_buffer.n578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9965\,
            in2 => \_gnd_net_\,
            in3 => \N__11069\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_4_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__11093\,
            in1 => \N__11129\,
            in2 => \N__10013\,
            in3 => \N__9939\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__10005\,
            in1 => \N__9990\,
            in2 => \N__9977\,
            in3 => \N__9974\,
            lcout => \receive_module.rx_counter.n3657\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_16_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9938\,
            in2 => \_gnd_net_\,
            in3 => \N__9966\,
            lcout => \receive_module.rx_counter.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.SYNC_45_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9967\,
            in1 => \N__9947\,
            in2 => \_gnd_net_\,
            in3 => \N__9941\,
            lcout => \DEBUG_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__15853\,
            in1 => \N__15911\,
            in2 => \N__15760\,
            in3 => \N__11304\,
            lcout => \line_buffer.n610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2390_2_lut_3_lut_4_lut_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__15847\,
            in1 => \N__15910\,
            in2 => \N__15759\,
            in3 => \N__11308\,
            lcout => \line_buffer.n512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i13_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__11310\,
            in1 => \N__15739\,
            in2 => \N__17838\,
            in3 => \N__15689\,
            lcout => \DEBUG_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21018\,
            ce => 'H',
            sr => \N__17690\
        );

    \receive_module.BRAM_ADDR__i3_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__15089\,
            in1 => \N__15113\,
            in2 => \N__17836\,
            in3 => \N__11314\,
            lcout => \RX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21018\,
            ce => 'H',
            sr => \N__17690\
        );

    \receive_module.BRAM_ADDR__i2_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__11311\,
            in1 => \N__15353\,
            in2 => \N__17840\,
            in3 => \N__15377\,
            lcout => \RX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21018\,
            ce => 'H',
            sr => \N__17690\
        );

    \receive_module.BRAM_ADDR__i1_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__17813\,
            in1 => \N__12980\,
            in2 => \N__13035\,
            in3 => \N__11313\,
            lcout => \RX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21018\,
            ce => 'H',
            sr => \N__17690\
        );

    \receive_module.BRAM_ADDR__i10_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__11309\,
            in1 => \N__15956\,
            in2 => \N__17837\,
            in3 => \N__15932\,
            lcout => \RX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21018\,
            ce => 'H',
            sr => \N__17690\
        );

    \receive_module.BRAM_ADDR__i9_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__13619\,
            in1 => \N__13598\,
            in2 => \N__17835\,
            in3 => \N__11315\,
            lcout => \RX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21018\,
            ce => 'H',
            sr => \N__17690\
        );

    \receive_module.BRAM_ADDR__i8_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__11312\,
            in1 => \N__13880\,
            in2 => \N__17839\,
            in3 => \N__13853\,
            lcout => \RX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21018\,
            ce => 'H',
            sr => \N__17690\
        );

    \transmit_module.Y_DELTA_PATTERN_i98_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10043\,
            lcout => \transmit_module.Y_DELTA_PATTERN_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22085\,
            ce => \N__10075\,
            sr => \N__20367\
        );

    \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10037\,
            lcout => \transmit_module.Y_DELTA_PATTERN_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22140\,
            ce => \N__10074\,
            sr => \N__20368\
        );

    \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10019\,
            lcout => \transmit_module.Y_DELTA_PATTERN_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22140\,
            ce => \N__10074\,
            sr => \N__20368\
        );

    \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10025\,
            lcout => \transmit_module.Y_DELTA_PATTERN_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22140\,
            ce => \N__10074\,
            sr => \N__20368\
        );

    \transmit_module.Y_DELTA_PATTERN_i97_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10142\,
            lcout => \transmit_module.Y_DELTA_PATTERN_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22140\,
            ce => \N__10074\,
            sr => \N__20368\
        );

    \transmit_module.Y_DELTA_PATTERN_i96_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10136\,
            lcout => \transmit_module.Y_DELTA_PATTERN_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22140\,
            ce => \N__10074\,
            sr => \N__20368\
        );

    \transmit_module.video_signal_controller.i3_3_lut_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__10123\,
            in1 => \_gnd_net_\,
            in2 => \N__11200\,
            in3 => \N__10111\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n8_adj_569_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1759_4_lut_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__11225\,
            in1 => \N__10099\,
            in2 => \N__10088\,
            in3 => \N__12045\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3029_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1777_4_lut_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__10739\,
            in1 => \N__10700\,
            in2 => \N__10085\,
            in3 => \N__12019\,
            lcout => \transmit_module.video_signal_controller.n2030\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_rep_21_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__10182\,
            in1 => \N__11168\,
            in2 => \_gnd_net_\,
            in3 => \N__10161\,
            lcout => \transmit_module.video_signal_controller.n3857\,
            ltout => \transmit_module.video_signal_controller.n3857_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2242_3_lut_4_lut_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__10738\,
            in1 => \N__10699\,
            in2 => \N__10082\,
            in3 => \N__12018\,
            lcout => \transmit_module.video_signal_controller.n3603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__rep_1_i0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__16568\,
            in1 => \N__12755\,
            in2 => \N__16511\,
            in3 => \N__19545\,
            lcout => \TX_ADDR_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__17497\,
            sr => \N__20609\
        );

    \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__19544\,
            in1 => \N__16261\,
            in2 => \N__20572\,
            in3 => \N__16213\,
            lcout => \transmit_module.n2125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_28_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__16260\,
            in1 => \N__20452\,
            in2 => \N__16221\,
            in3 => \N__19543\,
            lcout => \transmit_module.n3864\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1133_1_lut_2_lut_3_lut_4_lut_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111111111"
        )
    port map (
            in0 => \N__12044\,
            in1 => \N__12011\,
            in2 => \N__11974\,
            in3 => \N__19542\,
            lcout => n2404,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16259\,
            in2 => \_gnd_net_\,
            in3 => \N__16208\,
            lcout => \transmit_module.n3859\,
            ltout => \transmit_module.n3859_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1076_3_lut_4_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__16481\,
            in1 => \N__12965\,
            in2 => \N__10187\,
            in3 => \N__19589\,
            lcout => \transmit_module.BRAM_ADDR_13_N_256_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_20_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10730\,
            in2 => \_gnd_net_\,
            in3 => \N__10696\,
            lcout => \transmit_module.video_signal_controller.n3856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.old_VGA_HS_39_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16209\,
            lcout => \transmit_module.old_VGA_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_adj_14_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11226\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11172\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i37_4_lut_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100101110"
        )
    port map (
            in0 => \N__11147\,
            in1 => \N__10184\,
            in2 => \N__10166\,
            in3 => \N__10163\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_HS_54_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__10731\,
            in1 => \N__12017\,
            in2 => \N__10145\,
            in3 => \N__10697\,
            lcout => \ADV_HSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21948\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i6_3_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19249\,
            in1 => \N__16406\,
            in2 => \_gnd_net_\,
            in3 => \N__16435\,
            lcout => \transmit_module.n183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_19_3_lut_4_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__10729\,
            in1 => \N__10695\,
            in2 => \N__12053\,
            in3 => \N__12012\,
            lcout => \transmit_module.n3855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i7_3_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19253\,
            in1 => \N__16682\,
            in2 => \_gnd_net_\,
            in3 => \N__16701\,
            lcout => \transmit_module.n182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i7_3_lut_4_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__16702\,
            in1 => \N__12785\,
            in2 => \N__19727\,
            in3 => \N__19607\,
            lcout => \transmit_module.n214\,
            ltout => \transmit_module.n214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i6_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__20573\,
            in1 => \N__10661\,
            in2 => \N__10649\,
            in3 => \N__20206\,
            lcout => \transmit_module.TX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1683_4_lut_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__10918\,
            in1 => \N__10925\,
            in2 => \N__20681\,
            in3 => \N__20234\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i9_3_lut_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19257\,
            in1 => \N__12938\,
            in2 => \_gnd_net_\,
            in3 => \N__12955\,
            lcout => \transmit_module.n180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i6_3_lut_4_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__19616\,
            in1 => \N__12794\,
            in2 => \N__19737\,
            in3 => \N__16431\,
            lcout => \transmit_module.n215\,
            ltout => \transmit_module.n215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1680_4_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__20233\,
            in1 => \N__20605\,
            in2 => \N__10424\,
            in3 => \N__10204\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i5_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__10205\,
            in1 => \N__10193\,
            in2 => \N__20682\,
            in3 => \N__20235\,
            lcout => \transmit_module.TX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i9_3_lut_4_lut_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__19723\,
            in1 => \N__12956\,
            in2 => \N__12773\,
            in3 => \N__19615\,
            lcout => \transmit_module.n212\,
            ltout => \transmit_module.n212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i8_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__10919\,
            in1 => \N__20508\,
            in2 => \N__10910\,
            in3 => \N__20236\,
            lcout => \transmit_module.TX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i8_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10907\,
            lcout => \transmit_module.X_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21786\,
            ce => \N__12879\,
            sr => \N__18693\
        );

    \transmit_module.X_DELTA_PATTERN_i7_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10892\,
            lcout => \transmit_module.X_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21786\,
            ce => \N__12879\,
            sr => \N__18693\
        );

    \transmit_module.X_DELTA_PATTERN_i6_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10886\,
            lcout => \transmit_module.X_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21786\,
            ce => \N__12879\,
            sr => \N__18693\
        );

    \transmit_module.X_DELTA_PATTERN_i5_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10880\,
            lcout => \transmit_module.X_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21786\,
            ce => \N__12879\,
            sr => \N__18693\
        );

    \line_buffer.n3785_bdd_4_lut_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__10874\,
            in1 => \N__10862\,
            in2 => \N__10856\,
            in3 => \N__22930\,
            lcout => \line_buffer.n3788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__15917\,
            in1 => \N__15751\,
            in2 => \N__15855\,
            in3 => \N__11300\,
            lcout => \line_buffer.n577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_10_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__11298\,
            in1 => \N__15840\,
            in2 => \N__15764\,
            in3 => \N__15915\,
            lcout => \line_buffer.n513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i2393_2_lut_rep_18_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__17758\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11301\,
            lcout => \receive_module.n3854\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_adj_17_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__11135\,
            in1 => \N__11111\,
            in2 => \N__11105\,
            in3 => \N__11075\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3648_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2397_4_lut_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__11051\,
            in1 => \N__11045\,
            in2 => \N__11039\,
            in3 => \N__18845\,
            lcout => \DEBUG_c_5\,
            ltout => \DEBUG_c_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_7_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15746\,
            in1 => \N__15839\,
            in2 => \N__11036\,
            in3 => \N__15916\,
            lcout => \line_buffer.n641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_8_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15914\,
            in1 => \N__15747\,
            in2 => \N__15854\,
            in3 => \N__11299\,
            lcout => \line_buffer.n609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.FRAME_COUNTER_264__i0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13535\,
            in2 => \_gnd_net_\,
            in3 => \N__10937\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_0\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \receive_module.rx_counter.n3387\,
            clk => \N__21010\,
            ce => \N__16720\,
            sr => \N__13487\
        );

    \receive_module.rx_counter.FRAME_COUNTER_264__i1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13547\,
            in2 => \_gnd_net_\,
            in3 => \N__10934\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3387\,
            carryout => \receive_module.rx_counter.n3388\,
            clk => \N__21010\,
            ce => \N__16720\,
            sr => \N__13487\
        );

    \receive_module.rx_counter.FRAME_COUNTER_264__i2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13571\,
            in2 => \_gnd_net_\,
            in3 => \N__10931\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3388\,
            carryout => \receive_module.rx_counter.n3389\,
            clk => \N__21010\,
            ce => \N__16720\,
            sr => \N__13487\
        );

    \receive_module.rx_counter.FRAME_COUNTER_264__i3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13523\,
            in2 => \_gnd_net_\,
            in3 => \N__10928\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3389\,
            carryout => \receive_module.rx_counter.n3390\,
            clk => \N__21010\,
            ce => \N__16720\,
            sr => \N__13487\
        );

    \receive_module.rx_counter.FRAME_COUNTER_264__i4_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13583\,
            in2 => \_gnd_net_\,
            in3 => \N__11339\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3390\,
            carryout => \receive_module.rx_counter.n3391\,
            clk => \N__21010\,
            ce => \N__16720\,
            sr => \N__13487\
        );

    \receive_module.rx_counter.FRAME_COUNTER_264__i5_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13559\,
            in2 => \_gnd_net_\,
            in3 => \N__11336\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21010\,
            ce => \N__16720\,
            sr => \N__13487\
        );

    \receive_module.BRAM_ADDR__i7_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__14129\,
            in1 => \N__14105\,
            in2 => \N__17833\,
            in3 => \N__11320\,
            lcout => \RX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21014\,
            ce => 'H',
            sr => \N__17702\
        );

    \receive_module.BRAM_ADDR__i6_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__11317\,
            in1 => \N__17812\,
            in2 => \N__14357\,
            in3 => \N__14381\,
            lcout => \RX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21014\,
            ce => 'H',
            sr => \N__17702\
        );

    \receive_module.BRAM_ADDR__i5_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__14591\,
            in1 => \N__14611\,
            in2 => \N__17834\,
            in3 => \N__11319\,
            lcout => \RX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21014\,
            ce => 'H',
            sr => \N__17702\
        );

    \receive_module.BRAM_ADDR__i4_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__11316\,
            in1 => \N__17811\,
            in2 => \N__14846\,
            in3 => \N__14870\,
            lcout => \RX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21014\,
            ce => 'H',
            sr => \N__17702\
        );

    \receive_module.BRAM_ADDR__i0_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__13241\,
            in1 => \N__13268\,
            in2 => \N__17832\,
            in3 => \N__11318\,
            lcout => \RX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21014\,
            ce => 'H',
            sr => \N__17702\
        );

    \transmit_module.video_signal_controller.i1_3_lut_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__11234\,
            in1 => \N__11204\,
            in2 => \_gnd_net_\,
            in3 => \N__11177\,
            lcout => \transmit_module.video_signal_controller.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1753_4_lut_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__15660\,
            in1 => \N__16388\,
            in2 => \N__15620\,
            in3 => \N__15639\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3023_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__16366\,
            in1 => \N__16345\,
            in2 => \N__11393\,
            in3 => \N__11363\,
            lcout => \transmit_module.video_signal_controller.n3577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16324\,
            in2 => \_gnd_net_\,
            in3 => \N__16309\,
            lcout => \transmit_module.video_signal_controller.n3575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i487_3_lut_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__15638\,
            in1 => \N__15614\,
            in2 => \_gnd_net_\,
            in3 => \N__15659\,
            lcout => \transmit_module.video_signal_controller.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2335_3_lut_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__15618\,
            in1 => \N__16389\,
            in2 => \_gnd_net_\,
            in3 => \N__11351\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3697_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VS_55_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__15640\,
            in1 => \N__15677\,
            in2 => \N__11390\,
            in3 => \N__15661\,
            lcout => \ADV_VSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21667\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__17330\,
            in1 => \N__11387\,
            in2 => \N__16397\,
            in3 => \N__11350\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n6_adj_568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i3_4_lut_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__16294\,
            in1 => \N__11381\,
            in2 => \N__11375\,
            in3 => \N__11372\,
            lcout => \transmit_module.n3549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__17369\,
            in1 => \N__17347\,
            in2 => \_gnd_net_\,
            in3 => \N__16344\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i4_4_lut_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16293\,
            in1 => \N__16365\,
            in2 => \N__11366\,
            in3 => \N__11362\,
            lcout => \transmit_module.video_signal_controller.n2015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i12_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__12740\,
            in1 => \N__16577\,
            in2 => \N__16496\,
            in3 => \N__19590\,
            lcout => \TX_ADDR_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22084\,
            ce => \N__17498\,
            sr => \N__20366\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_16_3_lut_4_lut_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__12049\,
            in1 => \N__12023\,
            in2 => \N__11975\,
            in3 => \N__19549\,
            lcout => n3852,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i1_3_lut_4_lut_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__19548\,
            in1 => \N__19722\,
            in2 => \N__12686\,
            in3 => \N__16472\,
            lcout => \transmit_module.n220\,
            ltout => \transmit_module.n220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1670_4_lut_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__20384\,
            in1 => \N__16588\,
            in2 => \N__11957\,
            in3 => \N__20178\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i13_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21214\,
            in1 => \N__11735\,
            in2 => \_gnd_net_\,
            in3 => \N__17490\,
            lcout => \DEBUG_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22077\,
            ce => 'H',
            sr => \N__20613\
        );

    \transmit_module.video_signal_controller.mux_15_i2_3_lut_4_lut_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__19547\,
            in1 => \N__19721\,
            in2 => \N__12674\,
            in3 => \N__16544\,
            lcout => \transmit_module.n219\,
            ltout => \transmit_module.n219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1676_4_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__20383\,
            in1 => \N__12728\,
            in2 => \N__11729\,
            in3 => \N__20179\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_17_3_lut_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19546\,
            in1 => \N__16258\,
            in2 => \_gnd_net_\,
            in3 => \N__16220\,
            lcout => \transmit_module.n3853\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADV_R__i1_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22169\,
            lcout => n1850,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \ADV_R__i2_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17381\,
            lcout => n1849,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \ADV_R__i3_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18143\,
            lcout => n1848,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \ADV_R__i4_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18236\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n1847,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \ADV_R__i5_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20759\,
            lcout => n1846,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \ADV_R__i6_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18761\,
            lcout => n1845,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \ADV_R__i7_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12809\,
            lcout => n1844,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \ADV_R__i8_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18047\,
            lcout => \ADV_B_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \transmit_module.BRAM_ADDR__i0_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__16595\,
            in1 => \N__12278\,
            in2 => \N__20601\,
            in3 => \N__20194\,
            lcout => \transmit_module.TX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i3_3_lut_4_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__19707\,
            in1 => \N__16669\,
            in2 => \N__12656\,
            in3 => \N__19606\,
            lcout => \transmit_module.n218\,
            ltout => \transmit_module.n218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1677_4_lut_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__20490\,
            in1 => \N__12694\,
            in2 => \N__12269\,
            in3 => \N__20193\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i2_3_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19226\,
            in1 => \N__16517\,
            in2 => \_gnd_net_\,
            in3 => \N__16539\,
            lcout => \transmit_module.n187\,
            ltout => \transmit_module.n187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i1_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__12716\,
            in1 => \N__20512\,
            in2 => \N__12707\,
            in3 => \N__20195\,
            lcout => \transmit_module.TX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i2_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20196\,
            in1 => \N__20491\,
            in2 => \N__12698\,
            in3 => \N__12704\,
            lcout => \transmit_module.TX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i3_3_lut_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19227\,
            in1 => \N__16649\,
            in2 => \_gnd_net_\,
            in3 => \N__16668\,
            lcout => \transmit_module.n186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_2_lut_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16463\,
            in2 => \N__12932\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n204\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \transmit_module.n3336\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_3_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16538\,
            in2 => \_gnd_net_\,
            in3 => \N__12659\,
            lcout => \transmit_module.n203\,
            ltout => OPEN,
            carryin => \transmit_module.n3336\,
            carryout => \transmit_module.n3337\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_4_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16667\,
            in2 => \_gnd_net_\,
            in3 => \N__12644\,
            lcout => \transmit_module.n202\,
            ltout => OPEN,
            carryin => \transmit_module.n3337\,
            carryout => \transmit_module.n3338\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_5_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19768\,
            in2 => \_gnd_net_\,
            in3 => \N__12641\,
            lcout => \transmit_module.n201\,
            ltout => OPEN,
            carryin => \transmit_module.n3338\,
            carryout => \transmit_module.n3339\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_6_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16619\,
            in2 => \_gnd_net_\,
            in3 => \N__12797\,
            lcout => \transmit_module.n200\,
            ltout => OPEN,
            carryin => \transmit_module.n3339\,
            carryout => \transmit_module.n3340\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_7_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16427\,
            in2 => \_gnd_net_\,
            in3 => \N__12788\,
            lcout => \transmit_module.n199\,
            ltout => OPEN,
            carryin => \transmit_module.n3340\,
            carryout => \transmit_module.n3341\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_8_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16700\,
            in2 => \_gnd_net_\,
            in3 => \N__12779\,
            lcout => \transmit_module.n198\,
            ltout => OPEN,
            carryin => \transmit_module.n3341\,
            carryout => \transmit_module.n3342\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_9_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17315\,
            in2 => \_gnd_net_\,
            in3 => \N__12776\,
            lcout => \transmit_module.n197\,
            ltout => OPEN,
            carryin => \transmit_module.n3342\,
            carryout => \transmit_module.n3343\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_10_lut_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12953\,
            in2 => \_gnd_net_\,
            in3 => \N__12764\,
            lcout => \transmit_module.n196\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \transmit_module.n3344\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_11_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19634\,
            in2 => \_gnd_net_\,
            in3 => \N__12761\,
            lcout => \transmit_module.n195\,
            ltout => OPEN,
            carryin => \transmit_module.n3344\,
            carryout => \transmit_module.n3345\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_12_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19133\,
            in2 => \_gnd_net_\,
            in3 => \N__12758\,
            lcout => \transmit_module.n194\,
            ltout => OPEN,
            carryin => \transmit_module.n3345\,
            carryout => \transmit_module.n3346\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_13_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23133\,
            in2 => \_gnd_net_\,
            in3 => \N__12743\,
            lcout => \transmit_module.n193\,
            ltout => OPEN,
            carryin => \transmit_module.n3346\,
            carryout => \transmit_module.n3347\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_14_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22832\,
            in2 => \_gnd_net_\,
            in3 => \N__12731\,
            lcout => \transmit_module.n192\,
            ltout => OPEN,
            carryin => \transmit_module.n3347\,
            carryout => \transmit_module.n3348\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_15_lut_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21257\,
            in2 => \_gnd_net_\,
            in3 => \N__12968\,
            lcout => \transmit_module.n191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i9_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21828\,
            ce => \N__18466\,
            sr => \N__20661\
        );

    \transmit_module.ADDR_Y_COMPONENT__i8_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12954\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21828\,
            ce => \N__18466\,
            sr => \N__20661\
        );

    \transmit_module.X_DELTA_PATTERN_i0_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12911\,
            lcout => \transmit_module.X_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => \N__12874\,
            sr => \N__18702\
        );

    \transmit_module.X_DELTA_PATTERN_i1_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12905\,
            lcout => \transmit_module.X_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => \N__12874\,
            sr => \N__18702\
        );

    \transmit_module.X_DELTA_PATTERN_i2_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12887\,
            lcout => \transmit_module.X_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => \N__12874\,
            sr => \N__18702\
        );

    \transmit_module.X_DELTA_PATTERN_i4_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12899\,
            lcout => \transmit_module.X_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => \N__12874\,
            sr => \N__18702\
        );

    \transmit_module.X_DELTA_PATTERN_i3_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12893\,
            lcout => \transmit_module.X_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => \N__12874\,
            sr => \N__18702\
        );

    \line_buffer.dout_i6_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21284\,
            in1 => \N__12815\,
            in2 => \_gnd_net_\,
            in3 => \N__16790\,
            lcout => \TX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_VS_51_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17801\,
            lcout => \receive_module.rx_counter.PULSE_1HZ_N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_18_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13582\,
            in2 => \_gnd_net_\,
            in3 => \N__13570\,
            lcout => \receive_module.rx_counter.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i140_2_lut_rep_26_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__13499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17773\,
            lcout => \receive_module.rx_counter.n3862\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2331_2_lut_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13558\,
            in2 => \_gnd_net_\,
            in3 => \N__13546\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_4_lut_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__13534\,
            in1 => \N__13522\,
            in2 => \N__13511\,
            in3 => \N__13508\,
            lcout => \receive_module.rx_counter.n11\,
            ltout => \receive_module.rx_counter.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1294_2_lut_3_lut_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__17772\,
            in1 => \_gnd_net_\,
            in2 => \N__13502\,
            in3 => \N__13498\,
            lcout => \receive_module.rx_counter.n2562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_2_lut_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13269\,
            in2 => \_gnd_net_\,
            in3 => \N__13235\,
            lcout => \receive_module.n136\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \receive_module.n3323\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_3_lut_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13010\,
            in2 => \_gnd_net_\,
            in3 => \N__12971\,
            lcout => \receive_module.n135\,
            ltout => OPEN,
            carryin => \receive_module.n3323\,
            carryout => \receive_module.n3324\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_4_lut_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15387\,
            in2 => \_gnd_net_\,
            in3 => \N__15341\,
            lcout => \receive_module.n134\,
            ltout => OPEN,
            carryin => \receive_module.n3324\,
            carryout => \receive_module.n3325\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_5_lut_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15120\,
            in2 => \_gnd_net_\,
            in3 => \N__15080\,
            lcout => \receive_module.n133\,
            ltout => OPEN,
            carryin => \receive_module.n3325\,
            carryout => \receive_module.n3326\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_6_lut_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14871\,
            in2 => \_gnd_net_\,
            in3 => \N__14837\,
            lcout => \receive_module.n132\,
            ltout => OPEN,
            carryin => \receive_module.n3326\,
            carryout => \receive_module.n3327\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_7_lut_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14610\,
            in2 => \_gnd_net_\,
            in3 => \N__14585\,
            lcout => \receive_module.n131\,
            ltout => OPEN,
            carryin => \receive_module.n3327\,
            carryout => \receive_module.n3328\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_8_lut_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14382\,
            in2 => \_gnd_net_\,
            in3 => \N__14348\,
            lcout => \receive_module.n130\,
            ltout => OPEN,
            carryin => \receive_module.n3328\,
            carryout => \receive_module.n3329\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_9_lut_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14130\,
            in2 => \_gnd_net_\,
            in3 => \N__14099\,
            lcout => \receive_module.n129\,
            ltout => OPEN,
            carryin => \receive_module.n3329\,
            carryout => \receive_module.n3330\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_10_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13899\,
            in2 => \_gnd_net_\,
            in3 => \N__13841\,
            lcout => \receive_module.n128\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \receive_module.n3331\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_11_lut_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13638\,
            in2 => \_gnd_net_\,
            in3 => \N__13586\,
            lcout => \receive_module.n127\,
            ltout => OPEN,
            carryin => \receive_module.n3331\,
            carryout => \receive_module.n3332\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_12_lut_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15975\,
            in2 => \_gnd_net_\,
            in3 => \N__15920\,
            lcout => \receive_module.n126\,
            ltout => OPEN,
            carryin => \receive_module.n3332\,
            carryout => \receive_module.n3333\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i11_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15909\,
            in2 => \_gnd_net_\,
            in3 => \N__15863\,
            lcout => \RX_ADDR_11\,
            ltout => OPEN,
            carryin => \receive_module.n3333\,
            carryout => \receive_module.n3334\,
            clk => \N__21015\,
            ce => \N__15785\,
            sr => \N__17698\
        );

    \receive_module.BRAM_ADDR__i12_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15829\,
            in2 => \_gnd_net_\,
            in3 => \N__15788\,
            lcout => \RX_ADDR_12\,
            ltout => OPEN,
            carryin => \receive_module.n3334\,
            carryout => \receive_module.n3335\,
            clk => \N__21015\,
            ce => \N__15785\,
            sr => \N__17698\
        );

    \receive_module.add_12_15_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15766\,
            in2 => \_gnd_net_\,
            in3 => \N__15692\,
            lcout => \receive_module.n123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i0_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15676\,
            in2 => \_gnd_net_\,
            in3 => \N__15665\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_0\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \transmit_module.video_signal_controller.n3366\,
            clk => \N__22037\,
            ce => \N__17643\,
            sr => \N__17594\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15662\,
            in2 => \_gnd_net_\,
            in3 => \N__15644\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3366\,
            carryout => \transmit_module.video_signal_controller.n3367\,
            clk => \N__22037\,
            ce => \N__17643\,
            sr => \N__17594\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i2_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15641\,
            in2 => \_gnd_net_\,
            in3 => \N__15623\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3367\,
            carryout => \transmit_module.video_signal_controller.n3368\,
            clk => \N__22037\,
            ce => \N__17643\,
            sr => \N__17594\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i3_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15619\,
            in2 => \_gnd_net_\,
            in3 => \N__15599\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3368\,
            carryout => \transmit_module.video_signal_controller.n3369\,
            clk => \N__22037\,
            ce => \N__17643\,
            sr => \N__17594\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i4_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16393\,
            in2 => \_gnd_net_\,
            in3 => \N__16370\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3369\,
            carryout => \transmit_module.video_signal_controller.n3370\,
            clk => \N__22037\,
            ce => \N__17643\,
            sr => \N__17594\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i5_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16367\,
            in2 => \_gnd_net_\,
            in3 => \N__16349\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3370\,
            carryout => \transmit_module.video_signal_controller.n3371\,
            clk => \N__22037\,
            ce => \N__17643\,
            sr => \N__17594\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i6_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16346\,
            in2 => \_gnd_net_\,
            in3 => \N__16328\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3371\,
            carryout => \transmit_module.video_signal_controller.n3372\,
            clk => \N__22037\,
            ce => \N__17643\,
            sr => \N__17594\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i7_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16325\,
            in2 => \_gnd_net_\,
            in3 => \N__16313\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3372\,
            carryout => \transmit_module.video_signal_controller.n3373\,
            clk => \N__22037\,
            ce => \N__17643\,
            sr => \N__17594\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i8_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16310\,
            in2 => \_gnd_net_\,
            in3 => \N__16298\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_8\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \transmit_module.video_signal_controller.n3374\,
            clk => \N__22041\,
            ce => \N__17638\,
            sr => \N__17593\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i9_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16295\,
            in2 => \_gnd_net_\,
            in3 => \N__16280\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3374\,
            carryout => \transmit_module.video_signal_controller.n3375\,
            clk => \N__22041\,
            ce => \N__17638\,
            sr => \N__17593\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i10_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17348\,
            in2 => \_gnd_net_\,
            in3 => \N__16277\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3375\,
            carryout => \transmit_module.video_signal_controller.n3376\,
            clk => \N__22041\,
            ce => \N__17638\,
            sr => \N__17593\
        );

    \transmit_module.video_signal_controller.VGA_Y_265__i11_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17368\,
            in2 => \_gnd_net_\,
            in3 => \N__16274\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22041\,
            ce => \N__17638\,
            sr => \N__17593\
        );

    \transmit_module.video_signal_controller.i271_2_lut_3_lut_4_lut_rep_29_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__19568\,
            in1 => \N__20489\,
            in2 => \N__16271\,
            in3 => \N__16228\,
            lcout => \transmit_module.n3865\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i1_3_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19221\,
            in1 => \N__16445\,
            in2 => \_gnd_net_\,
            in3 => \N__16471\,
            lcout => \transmit_module.n188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__19222\,
            in1 => \N__16576\,
            in2 => \N__20600\,
            in3 => \N__19567\,
            lcout => \transmit_module.n2321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16543\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__18458\,
            sr => \N__20686\
        );

    \transmit_module.ADDR_Y_COMPONENT__i11_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23094\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__18458\,
            sr => \N__20686\
        );

    \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22926\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__18458\,
            sr => \N__20686\
        );

    \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21253\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__18458\,
            sr => \N__20686\
        );

    \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16470\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__18458\,
            sr => \N__20686\
        );

    \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16622\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => \N__18459\,
            sr => \N__20711\
        );

    \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16439\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => \N__18459\,
            sr => \N__20711\
        );

    \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16709\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => \N__18459\,
            sr => \N__20711\
        );

    \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17318\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => \N__18459\,
            sr => \N__20711\
        );

    \transmit_module.ADDR_Y_COMPONENT__i3_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19772\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => \N__18459\,
            sr => \N__20711\
        );

    \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16670\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => \N__18459\,
            sr => \N__20711\
        );

    \transmit_module.mux_12_i8_3_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16643\,
            in1 => \N__19251\,
            in2 => \_gnd_net_\,
            in3 => \N__17316\,
            lcout => \transmit_module.n181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i5_3_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19250\,
            in1 => \N__16637\,
            in2 => \_gnd_net_\,
            in3 => \N__16620\,
            lcout => \transmit_module.n184\,
            ltout => \transmit_module.n184_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i4_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20249\,
            in1 => \N__20619\,
            in2 => \N__16631\,
            in3 => \N__17291\,
            lcout => \transmit_module.TX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i5_3_lut_4_lut_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__16628\,
            in1 => \N__16621\,
            in2 => \N__19739\,
            in3 => \N__19609\,
            lcout => \transmit_module.n216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i8_3_lut_4_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__17317\,
            in1 => \N__16601\,
            in2 => \N__19738\,
            in3 => \N__19608\,
            lcout => \transmit_module.n213\,
            ltout => \transmit_module.n213_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i7_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__20250\,
            in1 => \N__20620\,
            in2 => \N__17321\,
            in3 => \N__17060\,
            lcout => \transmit_module.TX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i9_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__20746\,
            in1 => \N__20732\,
            in2 => \N__20685\,
            in3 => \N__20251\,
            lcout => \transmit_module.TX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1679_4_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__17297\,
            in1 => \N__17290\,
            in2 => \N__20701\,
            in3 => \N__20239\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i10_3_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19252\,
            in1 => \N__17066\,
            in2 => \_gnd_net_\,
            in3 => \N__19636\,
            lcout => \transmit_module.n179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1682_4_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__17059\,
            in1 => \N__17048\,
            in2 => \N__20700\,
            in3 => \N__20240\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3767_bdd_4_lut_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__16832\,
            in1 => \N__18338\,
            in2 => \N__16811\,
            in3 => \N__22907\,
            lcout => \line_buffer.n3770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2343_3_lut_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16784\,
            in1 => \N__16766\,
            in2 => \_gnd_net_\,
            in3 => \N__23125\,
            lcout => \line_buffer.n3705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16732\,
            in2 => \_gnd_net_\,
            in3 => \N__16754\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21006\,
            ce => \N__16721\,
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i23_1_lut_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17771\,
            lcout => \receive_module.BRAM_ADDR_13__N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1289_2_lut_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17534\,
            in2 => \_gnd_net_\,
            in3 => \N__17639\,
            lcout => \transmit_module.video_signal_controller.n2551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.SYNC_BUFF1_51_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17560\,
            lcout => \transmit_module.video_signal_controller.SYNC_BUFF1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.SYNC_BUFF2_52_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17540\,
            lcout => \transmit_module.video_signal_controller.SYNC_BUFF2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1716_4_lut_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110100"
        )
    port map (
            in0 => \N__19258\,
            in1 => \N__20232\,
            in2 => \N__20617\,
            in3 => \N__17518\,
            lcout => \transmit_module.n2039\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2353_3_lut_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17459\,
            in1 => \N__17441\,
            in2 => \_gnd_net_\,
            in3 => \N__23107\,
            lcout => \line_buffer.n3715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3827_bdd_4_lut_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__17426\,
            in1 => \N__18389\,
            in2 => \N__17405\,
            in3 => \N__22872\,
            lcout => OPEN,
            ltout => \line_buffer.n3830_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i1_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21277\,
            in2 => \N__17384\,
            in3 => \N__22703\,
            lcout => \TX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17364\,
            in2 => \_gnd_net_\,
            in3 => \N__17346\,
            lcout => \transmit_module.video_signal_controller.n3858\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i38_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17996\,
            lcout => \transmit_module.Y_DELTA_PATTERN_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => \N__17913\,
            sr => \N__20683\
        );

    \transmit_module.Y_DELTA_PATTERN_i37_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18035\,
            lcout => \transmit_module.Y_DELTA_PATTERN_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => \N__17913\,
            sr => \N__20683\
        );

    \transmit_module.Y_DELTA_PATTERN_i35_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18017\,
            lcout => \transmit_module.Y_DELTA_PATTERN_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => \N__17913\,
            sr => \N__20683\
        );

    \transmit_module.Y_DELTA_PATTERN_i34_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18029\,
            lcout => \transmit_module.Y_DELTA_PATTERN_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => \N__17913\,
            sr => \N__20683\
        );

    \transmit_module.Y_DELTA_PATTERN_i36_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18023\,
            lcout => \transmit_module.Y_DELTA_PATTERN_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => \N__17913\,
            sr => \N__20683\
        );

    \transmit_module.Y_DELTA_PATTERN_i39_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18011\,
            lcout => \transmit_module.Y_DELTA_PATTERN_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => \N__17913\,
            sr => \N__20683\
        );

    \transmit_module.Y_DELTA_PATTERN_i33_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17990\,
            lcout => \transmit_module.Y_DELTA_PATTERN_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => \N__17913\,
            sr => \N__20683\
        );

    \line_buffer.n3779_bdd_4_lut_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__22921\,
            in1 => \N__17885\,
            in2 => \N__17870\,
            in3 => \N__18065\,
            lcout => \line_buffer.n3782\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2425_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__18110\,
            in1 => \N__17849\,
            in2 => \N__21289\,
            in3 => \N__22919\,
            lcout => OPEN,
            ltout => \line_buffer.n3773_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i3_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__18299\,
            in1 => \N__18248\,
            in2 => \N__18239\,
            in3 => \N__21272\,
            lcout => \TX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2440_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18227\,
            in1 => \N__22918\,
            in2 => \N__18215\,
            in3 => \N__23093\,
            lcout => OPEN,
            ltout => \line_buffer.n3803_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3803_bdd_4_lut_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__22920\,
            in1 => \N__18194\,
            in2 => \N__18173\,
            in3 => \N__18170\,
            lcout => OPEN,
            ltout => \line_buffer.n3806_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i2_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__21271\,
            in1 => \_gnd_net_\,
            in2 => \N__18152\,
            in3 => \N__18149\,
            lcout => \TX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2344_3_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18134\,
            in1 => \N__18125\,
            in2 => \_gnd_net_\,
            in3 => \N__23091\,
            lcout => \line_buffer.n3706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2420_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18104\,
            in1 => \N__22908\,
            in2 => \N__18083\,
            in3 => \N__23090\,
            lcout => \line_buffer.n3779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2430_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__18059\,
            in1 => \N__18479\,
            in2 => \N__21290\,
            in3 => \N__22925\,
            lcout => OPEN,
            ltout => \line_buffer.n3791_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i7_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__18533\,
            in1 => \N__21276\,
            in2 => \N__18050\,
            in3 => \N__18260\,
            lcout => \TX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2340_3_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18515\,
            in1 => \N__18500\,
            in2 => \_gnd_net_\,
            in3 => \N__23092\,
            lcout => \line_buffer.n3702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i4_3_lut_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19259\,
            in1 => \N__18473\,
            in2 => \_gnd_net_\,
            in3 => \N__19763\,
            lcout => \transmit_module.n185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i10_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19128\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21827\,
            ce => \N__18467\,
            sr => \N__20618\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2460_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18428\,
            in1 => \N__22934\,
            in2 => \N__18407\,
            in3 => \N__23130\,
            lcout => \line_buffer.n3827\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2415_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18377\,
            in1 => \N__22928\,
            in2 => \N__18356\,
            in3 => \N__23131\,
            lcout => \line_buffer.n3767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2352_3_lut_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18332\,
            in1 => \N__18317\,
            in2 => \_gnd_net_\,
            in3 => \N__23129\,
            lcout => \line_buffer.n3714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2355_3_lut_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18287\,
            in1 => \N__18275\,
            in2 => \_gnd_net_\,
            in3 => \N__23143\,
            lcout => \line_buffer.n3717\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__19852\,
            in1 => \N__19822\,
            in2 => \_gnd_net_\,
            in3 => \N__19837\,
            lcout => \receive_module.rx_counter.n3547\,
            ltout => \receive_module.rx_counter.n3547_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2251_3_lut_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__19807\,
            in1 => \_gnd_net_\,
            in2 => \N__18863\,
            in3 => \N__21097\,
            lcout => \receive_module.rx_counter.n3613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_adj_15_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21096\,
            in1 => \N__19806\,
            in2 => \_gnd_net_\,
            in3 => \N__18860\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i35_4_lut_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010111001"
        )
    port map (
            in0 => \N__21061\,
            in1 => \N__21079\,
            in2 => \N__18854\,
            in3 => \N__18851\,
            lcout => \receive_module.rx_counter.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2406_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18836\,
            in1 => \N__22896\,
            in2 => \N__18818\,
            in3 => \N__23118\,
            lcout => OPEN,
            ltout => \line_buffer.n3761_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3761_bdd_4_lut_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__22897\,
            in1 => \N__18806\,
            in2 => \N__18788\,
            in3 => \N__18785\,
            lcout => \line_buffer.n3764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i5_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21261\,
            in1 => \N__18767\,
            in2 => \_gnd_net_\,
            in3 => \N__20774\,
            lcout => \TX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i32_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18749\,
            lcout => \transmit_module.Y_DELTA_PATTERN_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21479\,
            ce => \N__18708\,
            sr => \N__20577\
        );

    \line_buffer.i2356_3_lut_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18569\,
            in1 => \N__18551\,
            in2 => \_gnd_net_\,
            in3 => \N__23117\,
            lcout => \line_buffer.n3718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i11_3_lut_4_lut_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__19730\,
            in1 => \N__18527\,
            in2 => \N__19132\,
            in3 => \N__19593\,
            lcout => \transmit_module.n210\,
            ltout => \transmit_module.n210_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i10_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__19100\,
            in1 => \N__20598\,
            in2 => \N__19790\,
            in3 => \N__20237\,
            lcout => \transmit_module.TX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i4_3_lut_4_lut_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__19728\,
            in1 => \N__19764\,
            in2 => \N__19787\,
            in3 => \N__19591\,
            lcout => \transmit_module.n217\,
            ltout => \transmit_module.n217_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i3_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__19490\,
            in1 => \N__20599\,
            in2 => \N__19775\,
            in3 => \N__20238\,
            lcout => \transmit_module.TX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_15_i10_3_lut_4_lut_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__19729\,
            in1 => \N__19658\,
            in2 => \N__19646\,
            in3 => \N__19592\,
            lcout => \transmit_module.n211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1678_4_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__19496\,
            in1 => \N__19489\,
            in2 => \N__20666\,
            in3 => \N__20253\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i11_3_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19245\,
            in1 => \N__19139\,
            in2 => \_gnd_net_\,
            in3 => \N__19127\,
            lcout => \transmit_module.n178\,
            ltout => \transmit_module.n178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1685_4_lut_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__20587\,
            in1 => \N__19094\,
            in2 => \N__19088\,
            in3 => \N__20254\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_TVP_CLK_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i26_1_lut_rep_24_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19906\,
            lcout => n3860,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.X_263__i0_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19880\,
            in2 => \_gnd_net_\,
            in3 => \N__19874\,
            lcout => \receive_module.rx_counter.n10\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \receive_module.rx_counter.n3357\,
            clk => \N__21000\,
            ce => 'H',
            sr => \N__20899\
        );

    \receive_module.rx_counter.X_263__i1_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19871\,
            in2 => \_gnd_net_\,
            in3 => \N__19865\,
            lcout => \receive_module.rx_counter.n9\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3357\,
            carryout => \receive_module.rx_counter.n3358\,
            clk => \N__21000\,
            ce => 'H',
            sr => \N__20899\
        );

    \receive_module.rx_counter.X_263__i2_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19862\,
            in2 => \_gnd_net_\,
            in3 => \N__19856\,
            lcout => \receive_module.rx_counter.n8\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3358\,
            carryout => \receive_module.rx_counter.n3359\,
            clk => \N__21000\,
            ce => 'H',
            sr => \N__20899\
        );

    \receive_module.rx_counter.X_263__i3_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19853\,
            in2 => \_gnd_net_\,
            in3 => \N__19841\,
            lcout => \receive_module.rx_counter.X_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3359\,
            carryout => \receive_module.rx_counter.n3360\,
            clk => \N__21000\,
            ce => 'H',
            sr => \N__20899\
        );

    \receive_module.rx_counter.X_263__i4_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19838\,
            in2 => \_gnd_net_\,
            in3 => \N__19826\,
            lcout => \receive_module.rx_counter.X_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3360\,
            carryout => \receive_module.rx_counter.n3361\,
            clk => \N__21000\,
            ce => 'H',
            sr => \N__20899\
        );

    \receive_module.rx_counter.X_263__i5_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19823\,
            in2 => \_gnd_net_\,
            in3 => \N__19811\,
            lcout => \receive_module.rx_counter.X_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3361\,
            carryout => \receive_module.rx_counter.n3362\,
            clk => \N__21000\,
            ce => 'H',
            sr => \N__20899\
        );

    \receive_module.rx_counter.X_263__i6_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19808\,
            in2 => \_gnd_net_\,
            in3 => \N__19793\,
            lcout => \receive_module.rx_counter.X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3362\,
            carryout => \receive_module.rx_counter.n3363\,
            clk => \N__21000\,
            ce => 'H',
            sr => \N__20899\
        );

    \receive_module.rx_counter.X_263__i7_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21098\,
            in2 => \_gnd_net_\,
            in3 => \N__21083\,
            lcout => \receive_module.rx_counter.X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3363\,
            carryout => \receive_module.rx_counter.n3364\,
            clk => \N__21000\,
            ce => 'H',
            sr => \N__20899\
        );

    \receive_module.rx_counter.X_263__i8_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21080\,
            in2 => \_gnd_net_\,
            in3 => \N__21068\,
            lcout => \receive_module.rx_counter.X_8\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \receive_module.rx_counter.n3365\,
            clk => \N__21002\,
            ce => 'H',
            sr => \N__20903\
        );

    \receive_module.rx_counter.X_263__i9_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21062\,
            in2 => \_gnd_net_\,
            in3 => \N__21065\,
            lcout => \receive_module.rx_counter.X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21002\,
            ce => 'H',
            sr => \N__20903\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__20882\,
            in1 => \N__22892\,
            in2 => \N__20873\,
            in3 => \N__23136\,
            lcout => \line_buffer.n3833\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2359_3_lut_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20852\,
            in1 => \N__20834\,
            in2 => \_gnd_net_\,
            in3 => \N__23137\,
            lcout => \line_buffer.n3721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3833_bdd_4_lut_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__20822\,
            in1 => \N__20804\,
            in2 => \N__20798\,
            in3 => \N__22866\,
            lcout => \line_buffer.n3836\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i4_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__20768\,
            in1 => \N__21288\,
            in2 => \N__22340\,
            in3 => \N__21155\,
            lcout => \TX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1684_4_lut_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__20747\,
            in1 => \N__20728\,
            in2 => \N__20665\,
            in3 => \N__20255\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2358_3_lut_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22367\,
            in1 => \N__22358\,
            in2 => \_gnd_net_\,
            in3 => \N__23144\,
            lcout => \line_buffer.n3720\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2450_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__22328\,
            in1 => \N__22927\,
            in2 => \N__22313\,
            in3 => \N__23106\,
            lcout => \line_buffer.n3815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2337_3_lut_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22292\,
            in1 => \N__22277\,
            in2 => \_gnd_net_\,
            in3 => \N__23141\,
            lcout => \line_buffer.n3699\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3815_bdd_4_lut_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__22262\,
            in1 => \N__22241\,
            in2 => \N__22235\,
            in3 => \N__22932\,
            lcout => \line_buffer.n3818\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3821_bdd_4_lut_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__22211\,
            in1 => \N__23183\,
            in2 => \N__22196\,
            in3 => \N__22933\,
            lcout => OPEN,
            ltout => \line_buffer.n3824_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i0_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21291\,
            in2 => \N__22178\,
            in3 => \N__22175\,
            lcout => \TX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21924\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__21107\,
            in1 => \N__21308\,
            in2 => \N__21295\,
            in3 => \N__22931\,
            lcout => \line_buffer.n3797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2338_3_lut_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21146\,
            in1 => \N__21128\,
            in2 => \_gnd_net_\,
            in3 => \N__23134\,
            lcout => \line_buffer.n3700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2455_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__23135\,
            in1 => \N__23222\,
            in2 => \N__23201\,
            in3 => \N__22891\,
            lcout => \line_buffer.n3821\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2445_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23174\,
            in1 => \N__22864\,
            in2 => \N__23159\,
            in3 => \N__23142\,
            lcout => OPEN,
            ltout => \line_buffer.n3809_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3809_bdd_4_lut_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__22865\,
            in1 => \N__22742\,
            in2 => \N__22724\,
            in3 => \N__22721\,
            lcout => \line_buffer.n3812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_24_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
