// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Sun Sep 23 23:04:52 2018
//
// Verilog Description of module main
//

module main (DEBUG, TVP_CLK, TVP_HSYNC, TVP_VSYNC, TVP_VIDEO, LED, 
            ADV_HSYNC, ADV_VSYNC, ADV_R, ADV_G, ADV_B, ADV_CLK, 
            ADV_SYNC_N, ADV_BLANK_N) /* synthesis syn_module_defined=1 */ ;   // ../main.v(1[8:12])
    output [7:0]DEBUG;   // ../main.v(2[19:24])
    input TVP_CLK;   // ../main.v(3[13:20])
    input TVP_HSYNC;   // ../main.v(4[13:22])
    input TVP_VSYNC;   // ../main.v(5[13:22])
    input [9:0]TVP_VIDEO;   // ../main.v(6[19:28])
    output LED;   // ../main.v(7[14:17])
    output ADV_HSYNC;   // ../main.v(8[14:23])
    output ADV_VSYNC;   // ../main.v(9[14:23])
    output [7:0]ADV_R;   // ../main.v(10[19:24])
    output [7:0]ADV_G;   // ../main.v(11[19:24])
    output [7:0]ADV_B;   // ../main.v(12[19:24])
    output ADV_CLK;   // ../main.v(13[14:21])
    output ADV_SYNC_N;   // ../main.v(14[14:24])
    output ADV_BLANK_N;   // ../main.v(15[14:25])
    
    wire DEBUG_c_1_c /* synthesis SET_AS_NETWORK=DEBUG_c_1_c, is_clock=1 */ ;   // ../main.v(2[19:24])
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    
    wire GND_net, VCC_net, DEBUG_c_6, DEBUG_c_5, DEBUG_c_3, DEBUG_c_2, 
        DEBUG_c_0, TVP_HSYNC_c, TVP_VSYNC_c, TVP_VIDEO_c_9, TVP_VIDEO_c_8, 
        TVP_VIDEO_c_7, TVP_VIDEO_c_6, TVP_VIDEO_c_5, TVP_VIDEO_c_4, 
        TVP_VIDEO_c_3, TVP_VIDEO_c_2, LED_c, ADV_HSYNC_c, ADV_VSYNC_c, 
        ADV_B_c, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
        n28;
    wire [13:0]RX_ADDR;   // ../main.v(53[14:21])
    wire [13:0]TX_ADDR;   // ../main.v(72[14:21])
    wire [7:0]TX_DATA;   // ../main.v(73[13:20])
    
    wire n4214, n20, n2587, old_HS, n26, n25, n24, n23, n19, 
        n22, n21, n27, n2283, n4210, n691, n690, n659, n658, 
        n18;
    
    VCC i2 (.Y(VCC_net));
    RX receive_module (.GND_net(GND_net), .DEBUG_c_3(DEBUG_c_3), .\RX_ADDR[12] (RX_ADDR[12]), 
       .\RX_ADDR[11] (RX_ADDR[11]), .\RX_ADDR[10] (RX_ADDR[10]), .\RX_ADDR[9] (RX_ADDR[9]), 
       .\RX_ADDR[8] (RX_ADDR[8]), .\RX_ADDR[7] (RX_ADDR[7]), .\RX_ADDR[6] (RX_ADDR[6]), 
       .VCC_net(VCC_net), .\RX_ADDR[5] (RX_ADDR[5]), .TVP_HSYNC_c(TVP_HSYNC_c), 
       .old_HS(old_HS), .DEBUG_c_1_c(DEBUG_c_1_c), .TVP_VSYNC_c(TVP_VSYNC_c), 
       .DEBUG_c_6(DEBUG_c_6), .\RX_ADDR[0] (RX_ADDR[0]), .n4214(n4214), 
       .LED_c(LED_c), .n2283(n2283), .DEBUG_c_5(DEBUG_c_5), .n691(n691), 
       .\RX_ADDR[2] (RX_ADDR[2]), .\RX_ADDR[4] (RX_ADDR[4]), .\RX_ADDR[3] (RX_ADDR[3]), 
       .\RX_ADDR[1] (RX_ADDR[1]), .n659(n659), .n690(n690), .n658(n658)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(58[5] 69[29])
    TX transmit_module (.GND_net(GND_net), .ADV_CLK_c(ADV_CLK_c), .ADV_VSYNC_c(ADV_VSYNC_c), 
       .n28(n28), .ADV_HSYNC_c(ADV_HSYNC_c), .DEBUG_c_2(DEBUG_c_2), .n18(n18), 
       .n19(n19), .n4210(n4210), .n20(n20), .n21(n21), .n22(n22), 
       .n23(n23), .n24(n24), .n25(n25), .n26(n26), .n27(n27), .\TX_ADDR[12] (TX_ADDR[12]), 
       .\TX_ADDR[11] (TX_ADDR[11]), .DEBUG_c_6(DEBUG_c_6), .VCC_net(VCC_net), 
       .n2587(n2587)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(78[5] 91[26])
    SB_IO ADV_G_pad_4 (.PACKAGE_PIN(ADV_G[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1992));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_4.PULLUP = 1'b0;
    defparam ADV_G_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_5 (.PACKAGE_PIN(ADV_G[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1991));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_5.PULLUP = 1'b0;
    defparam ADV_G_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_6 (.PACKAGE_PIN(ADV_G[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1990));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_6.PULLUP = 1'b0;
    defparam ADV_G_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_3 (.PACKAGE_PIN(ADV_G[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1993));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_3.PULLUP = 1'b0;
    defparam ADV_G_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_7 (.PACKAGE_PIN(ADV_G[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_7.PULLUP = 1'b0;
    defparam ADV_G_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_0 (.PACKAGE_PIN(ADV_R[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1996));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_0.PULLUP = 1'b0;
    defparam ADV_R_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_1 (.PACKAGE_PIN(ADV_R[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1995));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_1.PULLUP = 1'b0;
    defparam ADV_R_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_2 (.PACKAGE_PIN(ADV_R[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1994));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_2.PULLUP = 1'b0;
    defparam ADV_R_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_3 (.PACKAGE_PIN(ADV_R[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1993));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_3.PULLUP = 1'b0;
    defparam ADV_R_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_4 (.PACKAGE_PIN(ADV_R[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1992));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_4.PULLUP = 1'b0;
    defparam ADV_R_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_5 (.PACKAGE_PIN(ADV_R[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1991));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_5.PULLUP = 1'b0;
    defparam ADV_R_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_6 (.PACKAGE_PIN(ADV_R[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1990));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_6.PULLUP = 1'b0;
    defparam ADV_R_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_7 (.PACKAGE_PIN(ADV_R[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_7.PULLUP = 1'b0;
    defparam ADV_R_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_VSYNC_pad (.PACKAGE_PIN(ADV_VSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_VSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_VSYNC_pad.PIN_TYPE = 6'b011001;
    defparam ADV_VSYNC_pad.PULLUP = 1'b0;
    defparam ADV_VSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_VSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_6 (.PACKAGE_PIN(DEBUG[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_6));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_6.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_6.PULLUP = 1'b0;
    defparam DEBUG_pad_6.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_HSYNC_pad (.PACKAGE_PIN(ADV_HSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_HSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_HSYNC_pad.PIN_TYPE = 6'b011001;
    defparam ADV_HSYNC_pad.PULLUP = 1'b0;
    defparam ADV_HSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_HSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_0 (.PACKAGE_PIN(DEBUG[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_0));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_0.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_0.PULLUP = 1'b0;
    defparam DEBUG_pad_0.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_1 (.PACKAGE_PIN(DEBUG[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_1_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_1.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_1.PULLUP = 1'b0;
    defparam DEBUG_pad_1.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_2 (.PACKAGE_PIN(DEBUG[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_2));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_2.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_2.PULLUP = 1'b0;
    defparam DEBUG_pad_2.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_3 (.PACKAGE_PIN(DEBUG[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_3));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_3.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_3.PULLUP = 1'b0;
    defparam DEBUG_pad_3.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_4 (.PACKAGE_PIN(DEBUG[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n4210));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_4.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_4.PULLUP = 1'b0;
    defparam DEBUG_pad_4.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_7 (.PACKAGE_PIN(DEBUG[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_7.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_7.PULLUP = 1'b0;
    defparam DEBUG_pad_7.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_5 (.PACKAGE_PIN(DEBUG[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_5));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_5.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_5.PULLUP = 1'b0;
    defparam DEBUG_pad_5.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_2 (.PACKAGE_PIN(TVP_VIDEO[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_2));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_2.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_2.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_2.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_3 (.PACKAGE_PIN(TVP_VIDEO[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_3));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_3.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_3.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_3.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_4 (.PACKAGE_PIN(TVP_VIDEO[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_4));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_4.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_4.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_4.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_5 (.PACKAGE_PIN(TVP_VIDEO[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_5));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_5.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_5.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_5.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_6 (.PACKAGE_PIN(TVP_VIDEO[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_6));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_6.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_6.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_6.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_7 (.PACKAGE_PIN(TVP_VIDEO[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_7));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_7.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_7.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_7.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_8 (.PACKAGE_PIN(TVP_VIDEO[8]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_8));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_8.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_8.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_8.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_8.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_9 (.PACKAGE_PIN(TVP_VIDEO[9]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_9));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_9.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_9.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_9.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_9.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VSYNC_pad (.PACKAGE_PIN(TVP_VSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VSYNC_pad.PIN_TYPE = 6'b000001;
    defparam TVP_VSYNC_pad.PULLUP = 1'b0;
    defparam TVP_VSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_VSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_HSYNC_pad (.PACKAGE_PIN(TVP_HSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_HSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_HSYNC_pad.PIN_TYPE = 6'b000001;
    defparam TVP_HSYNC_pad.PULLUP = 1'b0;
    defparam TVP_HSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_HSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO DEBUG_c_1_pad (.PACKAGE_PIN(TVP_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(DEBUG_c_1_c));   // ../main.v(3[13:20])
    defparam DEBUG_c_1_pad.PIN_TYPE = 6'b000001;
    defparam DEBUG_c_1_pad.PULLUP = 1'b0;
    defparam DEBUG_c_1_pad.NEG_TRIGGER = 1'b0;
    defparam DEBUG_c_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_BLANK_N_pad (.PACKAGE_PIN(ADV_BLANK_N), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_BLANK_N_pad.PIN_TYPE = 6'b011001;
    defparam ADV_BLANK_N_pad.PULLUP = 1'b0;
    defparam ADV_BLANK_N_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_BLANK_N_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_SYNC_N_pad (.PACKAGE_PIN(ADV_SYNC_N), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_SYNC_N_pad.PIN_TYPE = 6'b011001;
    defparam ADV_SYNC_N_pad.PULLUP = 1'b0;
    defparam ADV_SYNC_N_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_SYNC_N_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_CLK_pad (.PACKAGE_PIN(ADV_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(ADV_CLK_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_CLK_pad.PIN_TYPE = 6'b011001;
    defparam ADV_CLK_pad.PULLUP = 1'b0;
    defparam ADV_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_0 (.PACKAGE_PIN(ADV_B[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1996));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_0.PULLUP = 1'b0;
    defparam ADV_B_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_1 (.PACKAGE_PIN(ADV_B[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1995));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_1.PULLUP = 1'b0;
    defparam ADV_B_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_2 (.PACKAGE_PIN(ADV_B[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1994));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_2.PULLUP = 1'b0;
    defparam ADV_B_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_3 (.PACKAGE_PIN(ADV_B[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1993));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_3.PULLUP = 1'b0;
    defparam ADV_B_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_4 (.PACKAGE_PIN(ADV_B[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1992));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_4.PULLUP = 1'b0;
    defparam ADV_B_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_5 (.PACKAGE_PIN(ADV_B[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1991));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_5.PULLUP = 1'b0;
    defparam ADV_B_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_6 (.PACKAGE_PIN(ADV_B[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1990));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_6.PULLUP = 1'b0;
    defparam ADV_B_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_7 (.PACKAGE_PIN(ADV_B[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_7.PULLUP = 1'b0;
    defparam ADV_B_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_0 (.PACKAGE_PIN(ADV_G[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1996));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_0.PULLUP = 1'b0;
    defparam ADV_G_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_1 (.PACKAGE_PIN(ADV_G[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1995));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_1.PULLUP = 1'b0;
    defparam ADV_G_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_2 (.PACKAGE_PIN(ADV_G[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1994));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_2.PULLUP = 1'b0;
    defparam ADV_G_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_DFFNSR ADV_R__i2 (.Q(n1995), .C(ADV_CLK_c), .D(TX_DATA[1]), .R(n2587));   // ../main.v(96[9] 100[5])
    SB_DFFNSR ADV_R__i3 (.Q(n1994), .C(ADV_CLK_c), .D(TX_DATA[2]), .R(n2587));   // ../main.v(96[9] 100[5])
    SB_DFFNSR ADV_R__i4 (.Q(n1993), .C(ADV_CLK_c), .D(TX_DATA[3]), .R(n2587));   // ../main.v(96[9] 100[5])
    SB_DFFNSR ADV_R__i5 (.Q(n1992), .C(ADV_CLK_c), .D(TX_DATA[4]), .R(n2587));   // ../main.v(96[9] 100[5])
    SB_DFFNSR ADV_R__i6 (.Q(n1991), .C(ADV_CLK_c), .D(TX_DATA[5]), .R(n2587));   // ../main.v(96[9] 100[5])
    SB_DFFNSR ADV_R__i7 (.Q(n1990), .C(ADV_CLK_c), .D(TX_DATA[6]), .R(n2587));   // ../main.v(96[9] 100[5])
    SB_DFFNSR ADV_R__i8 (.Q(ADV_B_c), .C(ADV_CLK_c), .D(TX_DATA[7]), .R(n2587));   // ../main.v(96[9] 100[5])
    SB_DFFNSR ADV_R__i1 (.Q(n1996), .C(ADV_CLK_c), .D(TX_DATA[0]), .R(n2587));   // ../main.v(96[9] 100[5])
    GND i1 (.Y(GND_net));
    SB_LUT4 i284_3_lut_3_lut (.I0(TVP_HSYNC_c), .I1(TVP_VSYNC_c), .I2(old_HS), 
            .I3(GND_net), .O(n2283));   // ../main.v(4[13:22])
    defparam i284_3_lut_3_lut.LUT_INIT = 16'h7373;
    SB_LUT4 i28_1_lut_rep_23 (.I0(TVP_HSYNC_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4214));   // ../main.v(4[13:22])
    defparam i28_1_lut_rep_23.LUT_INIT = 16'h5555;
    DIV_BY_5 db5 (.DEBUG_c_1_c(DEBUG_c_1_c), .GND_net(GND_net), .DEBUG_c_0(DEBUG_c_0)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(28[11] 29[26])
    TX_PLL tx_pll (.DEBUG_c_1_c(DEBUG_c_1_c), .VCC_net(VCC_net), .GND_net(GND_net), 
           .ADV_CLK_c(ADV_CLK_c)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(21[9] 25[27])
    RAM line_buffer (.TX_DATA({TX_DATA}), .ADV_CLK_c(ADV_CLK_c), .\TX_ADDR[11] (TX_ADDR[11]), 
        .\TX_ADDR[12] (TX_ADDR[12]), .GND_net(GND_net), .DEBUG_c_2(DEBUG_c_2), 
        .\RX_ADDR[11] (RX_ADDR[11]), .\RX_ADDR[12] (RX_ADDR[12]), .DEBUG_c_5(DEBUG_c_5), 
        .DEBUG_c_3(DEBUG_c_3), .\RX_ADDR[0] (RX_ADDR[0]), .\RX_ADDR[1] (RX_ADDR[1]), 
        .\RX_ADDR[2] (RX_ADDR[2]), .\RX_ADDR[3] (RX_ADDR[3]), .\RX_ADDR[4] (RX_ADDR[4]), 
        .\RX_ADDR[5] (RX_ADDR[5]), .\RX_ADDR[6] (RX_ADDR[6]), .\RX_ADDR[7] (RX_ADDR[7]), 
        .\RX_ADDR[8] (RX_ADDR[8]), .\RX_ADDR[9] (RX_ADDR[9]), .\RX_ADDR[10] (RX_ADDR[10]), 
        .n28(n28), .n27(n27), .n26(n26), .n25(n25), .n24(n24), .n23(n23), 
        .n22(n22), .n21(n21), .n20(n20), .n19(n19), .n18(n18), .TVP_VIDEO_c_8(TVP_VIDEO_c_8), 
        .TVP_VIDEO_c_9(TVP_VIDEO_c_9), .DEBUG_c_1_c(DEBUG_c_1_c), .VCC_net(VCC_net), 
        .TVP_VIDEO_c_6(TVP_VIDEO_c_6), .TVP_VIDEO_c_7(TVP_VIDEO_c_7), .TVP_VIDEO_c_4(TVP_VIDEO_c_4), 
        .TVP_VIDEO_c_5(TVP_VIDEO_c_5), .TVP_VIDEO_c_2(TVP_VIDEO_c_2), .TVP_VIDEO_c_3(TVP_VIDEO_c_3), 
        .n658(n658), .n690(n690), .n659(n659), .n691(n691)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(103[6] 109[21])
    
endmodule
//
// Verilog Description of module RX
//

module RX (GND_net, DEBUG_c_3, \RX_ADDR[12] , \RX_ADDR[11] , \RX_ADDR[10] , 
           \RX_ADDR[9] , \RX_ADDR[8] , \RX_ADDR[7] , \RX_ADDR[6] , VCC_net, 
           \RX_ADDR[5] , TVP_HSYNC_c, old_HS, DEBUG_c_1_c, TVP_VSYNC_c, 
           DEBUG_c_6, \RX_ADDR[0] , n4214, LED_c, n2283, DEBUG_c_5, 
           n691, \RX_ADDR[2] , \RX_ADDR[4] , \RX_ADDR[3] , \RX_ADDR[1] , 
           n659, n690, n658) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output DEBUG_c_3;
    output \RX_ADDR[12] ;
    output \RX_ADDR[11] ;
    output \RX_ADDR[10] ;
    output \RX_ADDR[9] ;
    output \RX_ADDR[8] ;
    output \RX_ADDR[7] ;
    output \RX_ADDR[6] ;
    input VCC_net;
    output \RX_ADDR[5] ;
    input TVP_HSYNC_c;
    output old_HS;
    input DEBUG_c_1_c;
    input TVP_VSYNC_c;
    output DEBUG_c_6;
    output \RX_ADDR[0] ;
    input n4214;
    output LED_c;
    input n2283;
    output DEBUG_c_5;
    output n691;
    output \RX_ADDR[2] ;
    output \RX_ADDR[4] ;
    output \RX_ADDR[3] ;
    output \RX_ADDR[1] ;
    output n659;
    output n690;
    output n658;
    
    wire DEBUG_c_1_c /* synthesis SET_AS_NETWORK=DEBUG_c_1_c, is_clock=1 */ ;   // ../main.v(2[19:24])
    wire [9:0]O_X;   // ../rx.v(37[16:19])
    wire [8:0]O_Y;   // ../rx.v(38[16:19])
    
    wire n3699;
    wire [7:0]n2;
    
    wire n4212, n3705, n3704, n3703, n3702, n3701, n3700, n4213;
    
    SB_CARRY add_629_2 (.CI(GND_net), .I0(O_X[6]), .I1(O_Y[0]), .CO(n3699));
    SB_LUT4 i652_2_lut_org (.I0(O_X[9]), .I1(O_Y[0]), .I2(GND_net), .I3(GND_net), 
            .O(n2[3]));   // ../rx.v(62[30:39])
    defparam i652_2_lut_org.LUT_INIT = 16'h6666;
    SB_LUT4 i660_3_lut (.I0(O_Y[1]), .I1(O_X[9]), .I2(O_Y[0]), .I3(GND_net), 
            .O(n2[4]));   // ../rx.v(62[30:39])
    defparam i660_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i681_4_lut (.I0(O_Y[4]), .I1(O_Y[3]), .I2(O_X[9]), .I3(n4212), 
            .O(n2[7]));   // ../rx.v(62[30:39])
    defparam i681_4_lut.LUT_INIT = 16'h6aaa;
    SB_LUT4 add_629_9_lut (.I0(GND_net), .I1(n2[7]), .I2(O_Y[7]), .I3(n3705), 
            .O(DEBUG_c_3)) /* synthesis syn_instantiated=1 */ ;
    defparam add_629_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_629_8_lut (.I0(GND_net), .I1(n2[6]), .I2(O_Y[6]), .I3(n3704), 
            .O(\RX_ADDR[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_629_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_629_8 (.CI(n3704), .I0(n2[6]), .I1(O_Y[6]), .CO(n3705));
    SB_LUT4 add_629_7_lut (.I0(GND_net), .I1(n2[5]), .I2(O_Y[5]), .I3(n3703), 
            .O(\RX_ADDR[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_629_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_629_7 (.CI(n3703), .I0(n2[5]), .I1(O_Y[5]), .CO(n3704));
    SB_LUT4 add_629_6_lut (.I0(GND_net), .I1(n2[4]), .I2(O_Y[4]), .I3(n3702), 
            .O(\RX_ADDR[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_629_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_629_6 (.CI(n3702), .I0(n2[4]), .I1(O_Y[4]), .CO(n3703));
    SB_LUT4 add_629_5_lut (.I0(GND_net), .I1(n2[3]), .I2(O_Y[3]), .I3(n3701), 
            .O(\RX_ADDR[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_629_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_629_5 (.CI(n3701), .I0(n2[3]), .I1(O_Y[3]), .CO(n3702));
    SB_LUT4 add_629_4_lut (.I0(GND_net), .I1(O_X[8]), .I2(O_Y[2]), .I3(n3700), 
            .O(\RX_ADDR[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_629_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_629_4 (.CI(n3700), .I0(O_X[8]), .I1(O_Y[2]), .CO(n3701));
    SB_LUT4 add_629_3_lut (.I0(GND_net), .I1(O_X[7]), .I2(O_Y[1]), .I3(n3699), 
            .O(\RX_ADDR[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_629_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_629_3 (.CI(n3699), .I0(O_X[7]), .I1(O_Y[1]), .CO(n3700));
    SB_LUT4 add_629_2_lut (.I0(GND_net), .I1(O_X[6]), .I2(O_Y[0]), .I3(GND_net), 
            .O(\RX_ADDR[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam add_629_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i667_3_lut_4_lut (.I0(O_Y[1]), .I1(O_Y[0]), .I2(O_X[9]), .I3(O_Y[2]), 
            .O(n2[5]));   // ../rx.v(62[30:39])
    defparam i667_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i1_2_lut_rep_21_3_lut (.I0(O_Y[1]), .I1(O_Y[0]), .I2(O_Y[2]), 
            .I3(GND_net), .O(n4212));   // ../rx.v(62[30:39])
    defparam i1_2_lut_rep_21_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_rep_22 (.I0(O_Y[1]), .I1(O_Y[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4213));   // ../rx.v(62[30:39])
    defparam i1_2_lut_rep_22.LUT_INIT = 16'h8888;
    SB_LUT4 i674_3_lut_4_lut (.I0(O_Y[2]), .I1(n4213), .I2(O_X[9]), .I3(O_Y[3]), 
            .O(n2[6]));   // ../rx.v(62[30:39])
    defparam i674_3_lut_4_lut.LUT_INIT = 16'h7f80;
    O_COUNTER rx_counter (.GND_net(GND_net), .\O_Y[6] (O_Y[6]), .VCC_net(VCC_net), 
            .\RX_ADDR[5] (\RX_ADDR[5] ), .TVP_HSYNC_c(TVP_HSYNC_c), .old_HS(old_HS), 
            .DEBUG_c_1_c(DEBUG_c_1_c), .TVP_VSYNC_c(TVP_VSYNC_c), .DEBUG_c_6(DEBUG_c_6), 
            .\RX_ADDR[0] (\RX_ADDR[0] ), .n4214(n4214), .LED_c(LED_c), 
            .\O_Y[5] (O_Y[5]), .n2283(n2283), .\O_Y[4] (O_Y[4]), .\O_Y[3] (O_Y[3]), 
            .\O_Y[2] (O_Y[2]), .\O_Y[1] (O_Y[1]), .\RX_ADDR[12] (\RX_ADDR[12] ), 
            .DEBUG_c_5(DEBUG_c_5), .\RX_ADDR[11] (\RX_ADDR[11] ), .DEBUG_c_3(DEBUG_c_3), 
            .n691(n691), .\RX_ADDR[2] (\RX_ADDR[2] ), .\O_X[9] (O_X[9]), 
            .\O_Y[0] (O_Y[0]), .\RX_ADDR[4] (\RX_ADDR[4] ), .\RX_ADDR[3] (\RX_ADDR[3] ), 
            .\O_X[8] (O_X[8]), .\O_X[7] (O_X[7]), .\O_X[6] (O_X[6]), .\RX_ADDR[1] (\RX_ADDR[1] ), 
            .n659(n659), .n690(n690), .\O_Y[7] (O_Y[7]), .n658(n658)) /* synthesis syn_module_defined=1 */ ;   // ../rx.v(41[15] 49[41])
    
endmodule
//
// Verilog Description of module O_COUNTER
//

module O_COUNTER (GND_net, \O_Y[6] , VCC_net, \RX_ADDR[5] , TVP_HSYNC_c, 
            old_HS, DEBUG_c_1_c, TVP_VSYNC_c, DEBUG_c_6, \RX_ADDR[0] , 
            n4214, LED_c, \O_Y[5] , n2283, \O_Y[4] , \O_Y[3] , \O_Y[2] , 
            \O_Y[1] , \RX_ADDR[12] , DEBUG_c_5, \RX_ADDR[11] , DEBUG_c_3, 
            n691, \RX_ADDR[2] , \O_X[9] , \O_Y[0] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \O_X[8] , \O_X[7] , \O_X[6] , \RX_ADDR[1] , 
            n659, n690, \O_Y[7] , n658) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \O_Y[6] ;
    input VCC_net;
    output \RX_ADDR[5] ;
    input TVP_HSYNC_c;
    output old_HS;
    input DEBUG_c_1_c;
    input TVP_VSYNC_c;
    output DEBUG_c_6;
    output \RX_ADDR[0] ;
    input n4214;
    output LED_c;
    output \O_Y[5] ;
    input n2283;
    output \O_Y[4] ;
    output \O_Y[3] ;
    output \O_Y[2] ;
    output \O_Y[1] ;
    input \RX_ADDR[12] ;
    output DEBUG_c_5;
    input \RX_ADDR[11] ;
    input DEBUG_c_3;
    output n691;
    output \RX_ADDR[2] ;
    output \O_X[9] ;
    output \O_Y[0] ;
    output \RX_ADDR[4] ;
    output \RX_ADDR[3] ;
    output \O_X[8] ;
    output \O_X[7] ;
    output \O_X[6] ;
    output \RX_ADDR[1] ;
    output n659;
    output n690;
    output \O_Y[7] ;
    output n658;
    
    wire DEBUG_c_1_c /* synthesis SET_AS_NETWORK=DEBUG_c_1_c, is_clock=1 */ ;   // ../main.v(2[19:24])
    
    wire n3673;
    wire [8:0]Y;   // ../o_counter.v(48[19:20])
    
    wire n3674, n3716;
    wire [8:0]n303;
    
    wire n3672, n3669;
    wire [5:0]n29;
    wire [5:0]FRAME_COUNTER;   // ../o_counter.v(46[19:32])
    
    wire n3708, n3709, n3707;
    wire [9:0]X;   // ../o_counter.v(47[19:20])
    
    wire n3651, n3938, n3706, old_VS, n3717, SYNC_N_98;
    wire [9:0]n45;
    
    wire n12, n13, n4222, n2605, PULSE_1HZ_N_94, PULSE_1HZ_N_97, 
        n3671, n3715, n3652, n3714, n3670, n3713, n3712, n3676, 
        n3711, n3728, n3727, n3726, n3725, n3724, n3723, n3722, 
        n3721, n3650, n3675, n3655, n3710, n3654, n3653, n11, 
        n4, n4219, n3720, n3176, n3208, n4_adj_575, n3979, n3718, 
        O_VISIBLE_N_89, n3204, O_VISIBLE_N_86, n4_adj_576, n5;
    
    SB_CARRY add_65_7 (.CI(n3673), .I0(Y[5]), .I1(GND_net), .CO(n3674));
    SB_LUT4 sub_23_add_2_8_lut (.I0(GND_net), .I1(Y[6]), .I2(VCC_net), 
            .I3(n3716), .O(\O_Y[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_23_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_65_6_lut (.I0(GND_net), .I1(Y[4]), .I2(GND_net), .I3(n3672), 
            .O(n303[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_2 (.CI(VCC_net), .I0(Y[0]), .I1(GND_net), .CO(n3669));
    SB_LUT4 FRAME_COUNTER_278_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[3]), 
            .I3(n3708), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_278_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_278_add_4_5 (.CI(n3708), .I0(GND_net), .I1(FRAME_COUNTER[3]), 
            .CO(n3709));
    SB_LUT4 FRAME_COUNTER_278_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[2]), 
            .I3(n3707), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_278_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_29_add_2_4_lut (.I0(GND_net), .I1(X[5]), .I2(VCC_net), 
            .I3(n3651), .O(\RX_ADDR[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_29_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut (.I0(Y[5]), .I1(Y[6]), .I2(GND_net), .I3(GND_net), 
            .O(n3938));   // ../o_counter.v(53[21:30])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_65_6 (.CI(n3672), .I0(Y[4]), .I1(GND_net), .CO(n3673));
    SB_CARRY FRAME_COUNTER_278_add_4_4 (.CI(n3707), .I0(GND_net), .I1(FRAME_COUNTER[2]), 
            .CO(n3708));
    SB_DFF old_HS_50 (.Q(old_HS), .C(DEBUG_c_1_c), .D(TVP_HSYNC_c));   // ../o_counter.v(51[16] 80[12])
    SB_LUT4 FRAME_COUNTER_278_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[1]), 
            .I3(n3706), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_278_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF old_VS_51 (.Q(old_VS), .C(DEBUG_c_1_c), .D(TVP_VSYNC_c));   // ../o_counter.v(51[16] 80[12])
    SB_CARRY sub_23_add_2_8 (.CI(n3716), .I0(Y[6]), .I1(VCC_net), .CO(n3717));
    SB_DFF SYNC_45 (.Q(DEBUG_c_6), .C(DEBUG_c_1_c), .D(SYNC_N_98));   // ../o_counter.v(51[16] 80[12])
    SB_CARRY FRAME_COUNTER_278_add_4_3 (.CI(n3706), .I0(GND_net), .I1(FRAME_COUNTER[1]), 
            .CO(n3707));
    SB_DFFSR X_277__i1 (.Q(\RX_ADDR[0] ), .C(DEBUG_c_1_c), .D(n45[0]), 
            .R(n4214));   // ../o_counter.v(62[26:31])
    SB_LUT4 i4_2_lut (.I0(Y[8]), .I1(Y[3]), .I2(GND_net), .I3(GND_net), 
            .O(n12));
    defparam i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 FRAME_COUNTER_278_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[0]), 
            .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_278_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut (.I0(n3938), .I1(Y[4]), .I2(Y[7]), .I3(Y[1]), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR FRAME_COUNTER_278__i2 (.Q(FRAME_COUNTER[2]), .C(DEBUG_c_1_c), 
            .E(n4222), .D(n29[2]), .R(n2605));   // ../o_counter.v(72[46:63])
    SB_CARRY FRAME_COUNTER_278_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(FRAME_COUNTER[0]), 
            .CO(n3706));
    SB_DFFE PULSE_1HZ_48 (.Q(LED_c), .C(DEBUG_c_1_c), .E(n4222), .D(PULSE_1HZ_N_94));   // ../o_counter.v(51[16] 80[12])
    SB_LUT4 i2634_4_lut (.I0(n13), .I1(Y[2]), .I2(n12), .I3(Y[0]), .O(SYNC_N_98));   // ../o_counter.v(53[21:30])
    defparam i2634_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i29_1_lut (.I0(TVP_VSYNC_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(PULSE_1HZ_N_97));   // ../main.v(5[13:22])
    defparam i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_65_5_lut (.I0(GND_net), .I1(Y[3]), .I2(GND_net), .I3(n3671), 
            .O(n303[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_23_add_2_7_lut (.I0(GND_net), .I1(Y[5]), .I2(VCC_net), 
            .I3(n3715), .O(\O_Y[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_23_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_29_add_2_4 (.CI(n3651), .I0(X[5]), .I1(VCC_net), .CO(n3652));
    SB_CARRY sub_23_add_2_7 (.CI(n3715), .I0(Y[5]), .I1(VCC_net), .CO(n3716));
    SB_DFFESR Y__i0 (.Q(Y[0]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[0]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR FRAME_COUNTER_278__i0 (.Q(FRAME_COUNTER[0]), .C(DEBUG_c_1_c), 
            .E(n4222), .D(n29[0]), .R(n2605));   // ../o_counter.v(72[46:63])
    SB_CARRY add_65_5 (.CI(n3671), .I0(Y[3]), .I1(GND_net), .CO(n3672));
    SB_LUT4 sub_23_add_2_6_lut (.I0(GND_net), .I1(Y[4]), .I2(GND_net), 
            .I3(n3714), .O(\O_Y[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_23_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_65_4_lut (.I0(GND_net), .I1(Y[2]), .I2(GND_net), .I3(n3670), 
            .O(n303[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_4 (.CI(n3670), .I0(Y[2]), .I1(GND_net), .CO(n3671));
    SB_CARRY sub_23_add_2_6 (.CI(n3714), .I0(Y[4]), .I1(GND_net), .CO(n3715));
    SB_LUT4 sub_23_add_2_5_lut (.I0(GND_net), .I1(Y[3]), .I2(GND_net), 
            .I3(n3713), .O(\O_Y[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_23_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_23_add_2_5 (.CI(n3713), .I0(Y[3]), .I1(GND_net), .CO(n3714));
    SB_LUT4 sub_23_add_2_4_lut (.I0(GND_net), .I1(Y[2]), .I2(VCC_net), 
            .I3(n3712), .O(\O_Y[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_23_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_23_add_2_4 (.CI(n3712), .I0(Y[2]), .I1(VCC_net), .CO(n3713));
    SB_LUT4 add_65_10_lut (.I0(GND_net), .I1(Y[8]), .I2(GND_net), .I3(n3676), 
            .O(n303[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_23_add_2_3_lut (.I0(GND_net), .I1(Y[1]), .I2(VCC_net), 
            .I3(n3711), .O(\O_Y[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_23_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_23_add_2_3 (.CI(n3711), .I0(Y[1]), .I1(VCC_net), .CO(n3712));
    SB_LUT4 X_277_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(X[9]), 
            .I3(n3728), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 X_277_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(X[8]), 
            .I3(n3727), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_277_add_4_10 (.CI(n3727), .I0(GND_net), .I1(X[8]), .CO(n3728));
    SB_LUT4 i1_2_lut_4_lut (.I0(\RX_ADDR[12] ), .I1(DEBUG_c_5), .I2(\RX_ADDR[11] ), 
            .I3(DEBUG_c_3), .O(n691));   // ../o_counter.v(82[28:148])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 X_277_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(X[7]), 
            .I3(n3726), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_277_add_4_9 (.CI(n3726), .I0(GND_net), .I1(X[7]), .CO(n3727));
    SB_LUT4 X_277_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(X[6]), 
            .I3(n3725), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_277_add_4_8 (.CI(n3725), .I0(GND_net), .I1(X[6]), .CO(n3726));
    SB_LUT4 X_277_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(X[5]), 
            .I3(n3724), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_277_add_4_7 (.CI(n3724), .I0(GND_net), .I1(X[5]), .CO(n3725));
    SB_LUT4 X_277_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(X[4]), 
            .I3(n3723), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_277_add_4_6 (.CI(n3723), .I0(GND_net), .I1(X[4]), .CO(n3724));
    SB_LUT4 X_277_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(X[3]), 
            .I3(n3722), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_277_add_4_5 (.CI(n3722), .I0(GND_net), .I1(X[3]), .CO(n3723));
    SB_LUT4 X_277_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\RX_ADDR[2] ), 
            .I3(n3721), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_65_3_lut (.I0(GND_net), .I1(Y[1]), .I2(GND_net), .I3(n3669), 
            .O(n303[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_29_add_2_3 (.CI(n3650), .I0(X[4]), .I1(VCC_net), .CO(n3651));
    SB_LUT4 add_65_9_lut (.I0(GND_net), .I1(Y[7]), .I2(GND_net), .I3(n3675), 
            .O(n303[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_29_add_2_8_lut (.I0(GND_net), .I1(X[9]), .I2(VCC_net), 
            .I3(n3655), .O(\O_X[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_29_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_9 (.CI(n3675), .I0(Y[7]), .I1(GND_net), .CO(n3676));
    SB_LUT4 sub_23_add_2_2_lut (.I0(GND_net), .I1(Y[0]), .I2(GND_net), 
            .I3(VCC_net), .O(\O_Y[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_23_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_29_add_2_3_lut (.I0(GND_net), .I1(X[4]), .I2(VCC_net), 
            .I3(n3650), .O(\RX_ADDR[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_29_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_23_add_2_2 (.CI(VCC_net), .I0(Y[0]), .I1(GND_net), .CO(n3711));
    SB_CARRY add_65_3 (.CI(n3669), .I0(Y[1]), .I1(GND_net), .CO(n3670));
    SB_LUT4 FRAME_COUNTER_278_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[5]), 
            .I3(n3710), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_278_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_65_8_lut (.I0(GND_net), .I1(Y[6]), .I2(GND_net), .I3(n3674), 
            .O(n303[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 FRAME_COUNTER_278_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[4]), 
            .I3(n3709), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_278_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_29_add_2_2_lut (.I0(GND_net), .I1(X[3]), .I2(GND_net), 
            .I3(VCC_net), .O(\RX_ADDR[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_29_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_29_add_2_7_lut (.I0(GND_net), .I1(X[8]), .I2(VCC_net), 
            .I3(n3654), .O(\O_X[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_29_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_65_2_lut (.I0(GND_net), .I1(Y[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n303[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_8 (.CI(n3674), .I0(Y[6]), .I1(GND_net), .CO(n3675));
    SB_CARRY sub_29_add_2_7 (.CI(n3654), .I0(X[8]), .I1(VCC_net), .CO(n3655));
    SB_LUT4 sub_29_add_2_6_lut (.I0(GND_net), .I1(X[7]), .I2(GND_net), 
            .I3(n3653), .O(\O_X[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_29_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_29_add_2_6 (.CI(n3653), .I0(X[7]), .I1(GND_net), .CO(n3654));
    SB_CARRY FRAME_COUNTER_278_add_4_6 (.CI(n3709), .I0(GND_net), .I1(FRAME_COUNTER[4]), 
            .CO(n3710));
    SB_LUT4 sub_29_add_2_5_lut (.I0(GND_net), .I1(X[6]), .I2(VCC_net), 
            .I3(n3652), .O(\O_X[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_29_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_29_add_2_5 (.CI(n3652), .I0(X[6]), .I1(VCC_net), .CO(n3653));
    SB_CARRY sub_29_add_2_2 (.CI(VCC_net), .I0(X[3]), .I1(GND_net), .CO(n3650));
    SB_LUT4 add_65_7_lut (.I0(GND_net), .I1(Y[5]), .I2(GND_net), .I3(n3673), 
            .O(n303[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR X_277__i2 (.Q(\RX_ADDR[1] ), .C(DEBUG_c_1_c), .D(n45[1]), 
            .R(n4214));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_277__i3 (.Q(\RX_ADDR[2] ), .C(DEBUG_c_1_c), .D(n45[2]), 
            .R(n4214));   // ../o_counter.v(62[26:31])
    SB_LUT4 i1_2_lut_4_lut_adj_18 (.I0(\RX_ADDR[12] ), .I1(DEBUG_c_5), .I2(\RX_ADDR[11] ), 
            .I3(DEBUG_c_3), .O(n659));   // ../o_counter.v(82[28:148])
    defparam i1_2_lut_4_lut_adj_18.LUT_INIT = 16'h0080;
    SB_LUT4 i1360_2_lut_3_lut (.I0(old_VS), .I1(TVP_VSYNC_c), .I2(n11), 
            .I3(GND_net), .O(n2605));   // ../o_counter.v(65[16] 75[19])
    defparam i1360_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i150_2_lut_rep_31 (.I0(old_VS), .I1(TVP_VSYNC_c), .I2(GND_net), 
            .I3(GND_net), .O(n4222));   // ../o_counter.v(65[16] 75[19])
    defparam i150_2_lut_rep_31.LUT_INIT = 16'h2222;
    SB_DFFSR X_277__i4 (.Q(X[3]), .C(DEBUG_c_1_c), .D(n45[3]), .R(n4214));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_277__i5 (.Q(X[4]), .C(DEBUG_c_1_c), .D(n45[4]), .R(n4214));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_277__i6 (.Q(X[5]), .C(DEBUG_c_1_c), .D(n45[5]), .R(n4214));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_277__i7 (.Q(X[6]), .C(DEBUG_c_1_c), .D(n45[6]), .R(n4214));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_277__i8 (.Q(X[7]), .C(DEBUG_c_1_c), .D(n45[7]), .R(n4214));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_277__i9 (.Q(X[8]), .C(DEBUG_c_1_c), .D(n45[8]), .R(n4214));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_277__i10 (.Q(X[9]), .C(DEBUG_c_1_c), .D(n45[9]), .R(n4214));   // ../o_counter.v(62[26:31])
    SB_LUT4 i1_2_lut_4_lut_adj_19 (.I0(X[4]), .I1(X[5]), .I2(X[3]), .I3(X[7]), 
            .O(n4));   // ../o_counter.v(82[61:90])
    defparam i1_2_lut_4_lut_adj_19.LUT_INIT = 16'hfe00;
    SB_LUT4 i2_3_lut_rep_28 (.I0(X[4]), .I1(X[5]), .I2(X[3]), .I3(GND_net), 
            .O(n4219));   // ../o_counter.v(82[61:90])
    defparam i2_3_lut_rep_28.LUT_INIT = 16'hfefe;
    SB_CARRY X_277_add_4_4 (.CI(n3721), .I0(GND_net), .I1(\RX_ADDR[2] ), 
            .CO(n3722));
    SB_LUT4 X_277_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\RX_ADDR[1] ), 
            .I3(n3720), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1803_2_lut (.I0(Y[0]), .I1(Y[1]), .I2(GND_net), .I3(GND_net), 
            .O(n3176));
    defparam i1803_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY X_277_add_4_3 (.CI(n3720), .I0(GND_net), .I1(\RX_ADDR[1] ), 
            .CO(n3721));
    SB_LUT4 i1835_4_lut (.I0(Y[2]), .I1(Y[4]), .I2(Y[3]), .I3(n3176), 
            .O(n3208));
    defparam i1835_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 X_277_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\RX_ADDR[0] ), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam X_277_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR Y__i8 (.Q(Y[8]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[8]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_LUT4 i1_2_lut_adj_20 (.I0(X[9]), .I1(X[8]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_575));
    defparam i1_2_lut_adj_20.LUT_INIT = 16'heeee;
    SB_CARRY X_277_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\RX_ADDR[0] ), 
            .CO(n3720));
    SB_LUT4 i2_4_lut (.I0(Y[7]), .I1(Y[8]), .I2(n3208), .I3(n3938), 
            .O(n3979));
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_CARRY sub_23_add_2_10 (.CI(n3718), .I0(Y[8]), .I1(VCC_net), .CO(O_VISIBLE_N_89));
    SB_LUT4 i1831_4_lut (.I0(X[6]), .I1(X[9]), .I2(X[8]), .I3(n4), .O(n3204));
    defparam i1831_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_21 (.I0(X[6]), .I1(n4_adj_575), .I2(X[7]), .I3(n4219), 
            .O(O_VISIBLE_N_86));
    defparam i2_4_lut_adj_21.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_4_lut_adj_22 (.I0(\RX_ADDR[12] ), .I1(DEBUG_c_5), .I2(\RX_ADDR[11] ), 
            .I3(DEBUG_c_3), .O(n690));   // ../o_counter.v(82[28:148])
    defparam i1_2_lut_4_lut_adj_22.LUT_INIT = 16'h0800;
    SB_LUT4 sub_23_add_2_9_lut (.I0(GND_net), .I1(Y[7]), .I2(VCC_net), 
            .I3(n3717), .O(\O_Y[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_23_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(O_VISIBLE_N_86), .I1(O_VISIBLE_N_89), .I2(n3204), 
            .I3(n3979), .O(DEBUG_c_5));
    defparam i3_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_adj_23 (.I0(LED_c), .I1(n11), .I2(GND_net), .I3(GND_net), 
            .O(PULSE_1HZ_N_94));
    defparam i1_2_lut_adj_23.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_24 (.I0(FRAME_COUNTER[3]), .I1(FRAME_COUNTER[1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_576));
    defparam i1_2_lut_adj_24.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_25 (.I0(FRAME_COUNTER[2]), .I1(FRAME_COUNTER[4]), 
            .I2(GND_net), .I3(GND_net), .O(n5));
    defparam i1_2_lut_adj_25.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut_adj_26 (.I0(n5), .I1(FRAME_COUNTER[5]), .I2(FRAME_COUNTER[0]), 
            .I3(n4_adj_576), .O(n11));
    defparam i3_4_lut_adj_26.LUT_INIT = 16'hbfff;
    SB_DFFESR Y__i7 (.Q(Y[7]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[7]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i6 (.Q(Y[6]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[6]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i5 (.Q(Y[5]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[5]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i4 (.Q(Y[4]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[4]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i3 (.Q(Y[3]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[3]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i2 (.Q(Y[2]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[2]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i1 (.Q(Y[1]), .C(DEBUG_c_1_c), .E(n2283), .D(n303[1]), 
            .R(PULSE_1HZ_N_97));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR FRAME_COUNTER_278__i5 (.Q(FRAME_COUNTER[5]), .C(DEBUG_c_1_c), 
            .E(n4222), .D(n29[5]), .R(n2605));   // ../o_counter.v(72[46:63])
    SB_DFFESR FRAME_COUNTER_278__i4 (.Q(FRAME_COUNTER[4]), .C(DEBUG_c_1_c), 
            .E(n4222), .D(n29[4]), .R(n2605));   // ../o_counter.v(72[46:63])
    SB_DFFESR FRAME_COUNTER_278__i3 (.Q(FRAME_COUNTER[3]), .C(DEBUG_c_1_c), 
            .E(n4222), .D(n29[3]), .R(n2605));   // ../o_counter.v(72[46:63])
    SB_CARRY sub_23_add_2_9 (.CI(n3717), .I0(Y[7]), .I1(VCC_net), .CO(n3718));
    SB_LUT4 i1_2_lut_4_lut_adj_27 (.I0(\RX_ADDR[12] ), .I1(DEBUG_c_5), .I2(\RX_ADDR[11] ), 
            .I3(DEBUG_c_3), .O(n658));   // ../o_counter.v(82[28:148])
    defparam i1_2_lut_4_lut_adj_27.LUT_INIT = 16'h0008;
    SB_DFFESR FRAME_COUNTER_278__i1 (.Q(FRAME_COUNTER[1]), .C(DEBUG_c_1_c), 
            .E(n4222), .D(n29[1]), .R(n2605));   // ../o_counter.v(72[46:63])
    
endmodule
//
// Verilog Description of module TX
//

module TX (GND_net, ADV_CLK_c, ADV_VSYNC_c, n28, ADV_HSYNC_c, DEBUG_c_2, 
           n18, n19, n4210, n20, n21, n22, n23, n24, n25, 
           n26, n27, \TX_ADDR[12] , \TX_ADDR[11] , DEBUG_c_6, VCC_net, 
           n2587) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input ADV_CLK_c;
    output ADV_VSYNC_c;
    output n28;
    output ADV_HSYNC_c;
    output DEBUG_c_2;
    output n18;
    output n19;
    output n4210;
    output n20;
    output n21;
    output n22;
    output n23;
    output n24;
    output n25;
    output n26;
    output n27;
    output \TX_ADDR[12] ;
    output \TX_ADDR[11] ;
    input DEBUG_c_6;
    input VCC_net;
    output n2587;
    
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    
    wire n3663;
    wire [13:0]TX_ADDR;   // ../main.v(72[14:21])
    
    wire n3664;
    wire [99:0]Y_DELTA_PATTERN;   // ../tx.v(65[16:31])
    
    wire n2361;
    wire [13:0]n190;
    
    wire n3658, n3662, old_VGA_HS, n3668, n4225;
    wire [13:0]BRAM_ADDR_13__N_258;
    
    wire n2277, n2909;
    wire [13:0]ADDR_Y_COMPONENT;   // ../tx.v(66[16:32])
    wire [13:0]n174;
    
    wire n2305;
    wire [13:0]n205;
    
    wire n4211, n3659, n3926, n3910, n4220, n2315, n3661, n4224;
    wire [15:0]X_DELTA_PATTERN;   // ../tx.v(64[16:31])
    
    wire n3667, n3660, n3657, n3666, n3656, n3665;
    
    SB_CARRY add_13_10 (.CI(n3663), .I0(TX_ADDR[8]), .I1(GND_net), .CO(n3664));
    SB_DFFESS Y_DELTA_PATTERN_i92 (.Q(Y_DELTA_PATTERN[92]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[93]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i91 (.Q(Y_DELTA_PATTERN[91]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[92]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i90 (.Q(Y_DELTA_PATTERN[90]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[91]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i89 (.Q(Y_DELTA_PATTERN[89]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[90]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFF BRAM_ADDR__i0 (.Q(TX_ADDR[0]), .C(ADV_CLK_c), .D(n28));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i88 (.Q(Y_DELTA_PATTERN[88]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[89]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_LUT4 add_13_5_lut (.I0(GND_net), .I1(TX_ADDR[3]), .I2(GND_net), 
            .I3(n3658), .O(n190[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_9_lut (.I0(GND_net), .I1(TX_ADDR[7]), .I2(GND_net), 
            .I3(n3662), .O(n190[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR Y_DELTA_PATTERN_i87 (.Q(Y_DELTA_PATTERN[87]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[88]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i86 (.Q(Y_DELTA_PATTERN[86]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[87]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFF old_VGA_HS_34 (.Q(old_VGA_HS), .C(ADV_CLK_c), .D(ADV_HSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i85 (.Q(Y_DELTA_PATTERN[85]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[86]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_LUT4 add_13_15_lut (.I0(GND_net), .I1(DEBUG_c_2), .I2(GND_net), 
            .I3(n3668), .O(n190[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS Y_DELTA_PATTERN_i84 (.Q(Y_DELTA_PATTERN[84]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[85]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i83 (.Q(Y_DELTA_PATTERN[83]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[84]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i82 (.Q(Y_DELTA_PATTERN[82]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[83]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i81 (.Q(Y_DELTA_PATTERN[81]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[82]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_LUT4 i1533_3_lut (.I0(DEBUG_c_2), .I1(BRAM_ADDR_13__N_258[13]), .I2(n2277), 
            .I3(GND_net), .O(n2909));   // ../tx.v(72[12] 93[8])
    defparam i1533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_12_i11_3_lut (.I0(ADDR_Y_COMPONENT[10]), .I1(TX_ADDR[10]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[10]));   // ../tx.v(82[30:81])
    defparam mux_12_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF BRAM_ADDR__i10 (.Q(TX_ADDR[10]), .C(ADV_CLK_c), .D(n18));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i80 (.Q(Y_DELTA_PATTERN[80]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[81]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i79 (.Q(Y_DELTA_PATTERN[79]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[80]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i78 (.Q(Y_DELTA_PATTERN[78]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[79]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i77 (.Q(Y_DELTA_PATTERN[77]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[78]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i4 (.Q(ADDR_Y_COMPONENT[4]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[4]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_CARRY add_13_9 (.CI(n3662), .I0(TX_ADDR[7]), .I1(GND_net), .CO(n3663));
    SB_DFF BRAM_ADDR__i9 (.Q(TX_ADDR[9]), .C(ADV_CLK_c), .D(n19));   // ../tx.v(72[12] 93[8])
    SB_LUT4 i1773_4_lut (.I0(n205[10]), .I1(ADV_VSYNC_c), .I2(n174[10]), 
            .I3(n4211), .O(n18));   // ../tx.v(72[12] 93[8])
    defparam i1773_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_13_5 (.CI(n3658), .I0(TX_ADDR[3]), .I1(GND_net), .CO(n3659));
    SB_LUT4 i1762_4_lut (.I0(ADV_VSYNC_c), .I1(n4210), .I2(Y_DELTA_PATTERN[0]), 
            .I3(n4211), .O(n2277));
    defparam i1762_4_lut.LUT_INIT = 16'hafee;
    SB_DFF BRAM_ADDR__i8 (.Q(TX_ADDR[8]), .C(ADV_CLK_c), .D(n20));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i97 (.Q(Y_DELTA_PATTERN[97]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[98]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFF BRAM_ADDR__i7 (.Q(TX_ADDR[7]), .C(ADV_CLK_c), .D(n21));   // ../tx.v(72[12] 93[8])
    SB_DFF BRAM_ADDR__i6 (.Q(TX_ADDR[6]), .C(ADV_CLK_c), .D(n22));   // ../tx.v(72[12] 93[8])
    SB_DFF BRAM_ADDR__i5 (.Q(TX_ADDR[5]), .C(ADV_CLK_c), .D(n23));   // ../tx.v(72[12] 93[8])
    SB_DFF BRAM_ADDR__i4 (.Q(TX_ADDR[4]), .C(ADV_CLK_c), .D(n24));   // ../tx.v(72[12] 93[8])
    SB_DFF BRAM_ADDR__i3 (.Q(TX_ADDR[3]), .C(ADV_CLK_c), .D(n25));   // ../tx.v(72[12] 93[8])
    SB_DFF BRAM_ADDR__i2 (.Q(TX_ADDR[2]), .C(ADV_CLK_c), .D(n26));   // ../tx.v(72[12] 93[8])
    SB_DFF BRAM_ADDR__i1 (.Q(TX_ADDR[1]), .C(ADV_CLK_c), .D(n27));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i76 (.Q(Y_DELTA_PATTERN[76]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[77]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_LUT4 i2_4_lut (.I0(ADV_VSYNC_c), .I1(n3926), .I2(n3910), .I3(n4220), 
            .O(n2315));   // ../tx.v(78[18] 90[12])
    defparam i2_4_lut.LUT_INIT = 16'heeea;
    SB_LUT4 add_13_8_lut (.I0(GND_net), .I1(TX_ADDR[6]), .I2(GND_net), 
            .I3(n3661), .O(n190[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS Y_DELTA_PATTERN_i75 (.Q(Y_DELTA_PATTERN[75]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[76]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i74 (.Q(Y_DELTA_PATTERN[74]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[75]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i73 (.Q(Y_DELTA_PATTERN[73]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[74]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i96 (.Q(Y_DELTA_PATTERN[96]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[97]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i95 (.Q(Y_DELTA_PATTERN[95]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[96]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i72 (.Q(Y_DELTA_PATTERN[72]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[73]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i71 (.Q(Y_DELTA_PATTERN[71]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[72]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i70 (.Q(Y_DELTA_PATTERN[70]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[71]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i69 (.Q(Y_DELTA_PATTERN[69]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[70]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i68 (.Q(Y_DELTA_PATTERN[68]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[69]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i67 (.Q(Y_DELTA_PATTERN[67]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[68]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i66 (.Q(Y_DELTA_PATTERN[66]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[67]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i65 (.Q(Y_DELTA_PATTERN[65]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[66]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i64 (.Q(Y_DELTA_PATTERN[64]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[65]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i63 (.Q(Y_DELTA_PATTERN[63]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[64]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i62 (.Q(Y_DELTA_PATTERN[62]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[63]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i61 (.Q(Y_DELTA_PATTERN[61]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[62]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i60 (.Q(Y_DELTA_PATTERN[60]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[61]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i59 (.Q(Y_DELTA_PATTERN[59]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[60]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i58 (.Q(Y_DELTA_PATTERN[58]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[59]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i57 (.Q(Y_DELTA_PATTERN[57]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[58]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i56 (.Q(Y_DELTA_PATTERN[56]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[57]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i55 (.Q(Y_DELTA_PATTERN[55]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[56]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i54 (.Q(Y_DELTA_PATTERN[54]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[55]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i53 (.Q(Y_DELTA_PATTERN[53]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[54]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i52 (.Q(Y_DELTA_PATTERN[52]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[53]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i51 (.Q(Y_DELTA_PATTERN[51]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[52]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i50 (.Q(Y_DELTA_PATTERN[50]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[51]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i49 (.Q(Y_DELTA_PATTERN[49]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[50]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i48 (.Q(Y_DELTA_PATTERN[48]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[49]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i47 (.Q(Y_DELTA_PATTERN[47]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[48]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i46 (.Q(Y_DELTA_PATTERN[46]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[47]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i45 (.Q(Y_DELTA_PATTERN[45]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[46]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i44 (.Q(Y_DELTA_PATTERN[44]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[45]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i43 (.Q(Y_DELTA_PATTERN[43]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[44]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i42 (.Q(Y_DELTA_PATTERN[42]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[43]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i41 (.Q(Y_DELTA_PATTERN[41]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[42]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i40 (.Q(Y_DELTA_PATTERN[40]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[41]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i39 (.Q(Y_DELTA_PATTERN[39]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[40]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i38 (.Q(Y_DELTA_PATTERN[38]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[39]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i37 (.Q(Y_DELTA_PATTERN[37]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[38]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i36 (.Q(Y_DELTA_PATTERN[36]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[37]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i35 (.Q(Y_DELTA_PATTERN[35]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[36]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i34 (.Q(Y_DELTA_PATTERN[34]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[35]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i33 (.Q(Y_DELTA_PATTERN[33]), .C(ADV_CLK_c), 
            .E(n4225), .D(Y_DELTA_PATTERN[34]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i32 (.Q(Y_DELTA_PATTERN[32]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[33]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i31 (.Q(Y_DELTA_PATTERN[31]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[32]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i30 (.Q(Y_DELTA_PATTERN[30]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[31]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i29 (.Q(Y_DELTA_PATTERN[29]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[30]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i28 (.Q(Y_DELTA_PATTERN[28]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[29]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i27 (.Q(Y_DELTA_PATTERN[27]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[28]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i26 (.Q(Y_DELTA_PATTERN[26]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[27]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i25 (.Q(Y_DELTA_PATTERN[25]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[26]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i24 (.Q(Y_DELTA_PATTERN[24]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[25]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i23 (.Q(Y_DELTA_PATTERN[23]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[24]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i22 (.Q(Y_DELTA_PATTERN[22]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[23]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i21 (.Q(Y_DELTA_PATTERN[21]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[22]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i20 (.Q(Y_DELTA_PATTERN[20]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[21]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i19 (.Q(Y_DELTA_PATTERN[19]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[20]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i18 (.Q(Y_DELTA_PATTERN[18]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[19]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i17 (.Q(Y_DELTA_PATTERN[17]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[18]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i16 (.Q(Y_DELTA_PATTERN[16]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[17]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i15 (.Q(Y_DELTA_PATTERN[15]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[16]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i14 (.Q(Y_DELTA_PATTERN[14]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[15]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i13 (.Q(Y_DELTA_PATTERN[13]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[14]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i12 (.Q(Y_DELTA_PATTERN[12]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[13]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i11 (.Q(Y_DELTA_PATTERN[11]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[12]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i10 (.Q(Y_DELTA_PATTERN[10]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[11]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i9 (.Q(Y_DELTA_PATTERN[9]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[10]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i8 (.Q(Y_DELTA_PATTERN[8]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[9]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i7 (.Q(Y_DELTA_PATTERN[7]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[8]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i6 (.Q(Y_DELTA_PATTERN[6]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[7]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i5 (.Q(Y_DELTA_PATTERN[5]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[6]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i4 (.Q(Y_DELTA_PATTERN[4]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[5]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i3 (.Q(Y_DELTA_PATTERN[3]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[4]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i2 (.Q(Y_DELTA_PATTERN[2]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[3]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i1 (.Q(Y_DELTA_PATTERN[1]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[2]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS X_DELTA_PATTERN_i15 (.Q(X_DELTA_PATTERN[15]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[0]), .S(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR X_DELTA_PATTERN_i14 (.Q(X_DELTA_PATTERN[14]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[15]), .R(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i3 (.Q(ADDR_Y_COMPONENT[3]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[3]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i2 (.Q(ADDR_Y_COMPONENT[2]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[2]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i1 (.Q(ADDR_Y_COMPONENT[1]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[1]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR BRAM_ADDR__i12 (.Q(\TX_ADDR[12] ), .C(ADV_CLK_c), .E(n2277), 
            .D(BRAM_ADDR_13__N_258[12]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_LUT4 mux_12_i1_3_lut (.I0(ADDR_Y_COMPONENT[0]), .I1(TX_ADDR[0]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[0]));   // ../tx.v(82[30:81])
    defparam mux_12_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1757_4_lut (.I0(n205[0]), .I1(ADV_VSYNC_c), .I2(n174[0]), 
            .I3(n4211), .O(n28));   // ../tx.v(72[12] 93[8])
    defparam i1757_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_13_14_lut (.I0(GND_net), .I1(\TX_ADDR[12] ), .I2(GND_net), 
            .I3(n3667), .O(n190[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_12_i2_3_lut (.I0(ADDR_Y_COMPONENT[1]), .I1(TX_ADDR[1]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[1]));   // ../tx.v(82[30:81])
    defparam mux_12_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1764_4_lut (.I0(n205[1]), .I1(ADV_VSYNC_c), .I2(n174[1]), 
            .I3(n4211), .O(n27));   // ../tx.v(72[12] 93[8])
    defparam i1764_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i3_3_lut (.I0(ADDR_Y_COMPONENT[2]), .I1(TX_ADDR[2]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[2]));   // ../tx.v(82[30:81])
    defparam mux_12_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1765_4_lut (.I0(n205[2]), .I1(ADV_VSYNC_c), .I2(n174[2]), 
            .I3(n4211), .O(n26));   // ../tx.v(72[12] 93[8])
    defparam i1765_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_13_14 (.CI(n3667), .I0(\TX_ADDR[12] ), .I1(GND_net), 
            .CO(n3668));
    SB_CARRY add_13_8 (.CI(n3661), .I0(TX_ADDR[6]), .I1(GND_net), .CO(n3662));
    SB_LUT4 add_13_7_lut (.I0(GND_net), .I1(TX_ADDR[5]), .I2(GND_net), 
            .I3(n3660), .O(n190[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_4_lut (.I0(GND_net), .I1(TX_ADDR[2]), .I2(GND_net), 
            .I3(n3657), .O(n190[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_4 (.CI(n3657), .I0(TX_ADDR[2]), .I1(GND_net), .CO(n3658));
    SB_CARRY add_13_7 (.CI(n3660), .I0(TX_ADDR[5]), .I1(GND_net), .CO(n3661));
    SB_LUT4 add_13_6_lut (.I0(GND_net), .I1(TX_ADDR[4]), .I2(GND_net), 
            .I3(n3659), .O(n190[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_13_lut (.I0(GND_net), .I1(\TX_ADDR[11] ), .I2(GND_net), 
            .I3(n3666), .O(n190[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_13 (.CI(n3666), .I0(\TX_ADDR[11] ), .I1(GND_net), 
            .CO(n3667));
    SB_LUT4 add_13_3_lut (.I0(GND_net), .I1(TX_ADDR[1]), .I2(GND_net), 
            .I3(n3656), .O(n190[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_12_lut (.I0(GND_net), .I1(TX_ADDR[10]), .I2(GND_net), 
            .I3(n3665), .O(n190[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_12 (.CI(n3665), .I0(TX_ADDR[10]), .I1(GND_net), .CO(n3666));
    SB_LUT4 add_13_11_lut (.I0(GND_net), .I1(TX_ADDR[9]), .I2(GND_net), 
            .I3(n3664), .O(n190[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_3 (.CI(n3656), .I0(TX_ADDR[1]), .I1(GND_net), .CO(n3657));
    SB_CARRY add_13_11 (.CI(n3664), .I0(TX_ADDR[9]), .I1(GND_net), .CO(n3665));
    SB_LUT4 add_13_10_lut (.I0(GND_net), .I1(TX_ADDR[8]), .I2(GND_net), 
            .I3(n3663), .O(n190[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_2_lut (.I0(GND_net), .I1(TX_ADDR[0]), .I2(X_DELTA_PATTERN[0]), 
            .I3(GND_net), .O(n190[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_2 (.CI(GND_net), .I0(TX_ADDR[0]), .I1(X_DELTA_PATTERN[0]), 
            .CO(n3656));
    SB_CARRY add_13_6 (.CI(n3659), .I0(TX_ADDR[4]), .I1(GND_net), .CO(n3660));
    SB_LUT4 mux_12_i4_3_lut (.I0(ADDR_Y_COMPONENT[3]), .I1(TX_ADDR[3]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[3]));   // ../tx.v(82[30:81])
    defparam mux_12_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1766_4_lut (.I0(n205[3]), .I1(ADV_VSYNC_c), .I2(n174[3]), 
            .I3(n4211), .O(n25));   // ../tx.v(72[12] 93[8])
    defparam i1766_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i5_3_lut (.I0(ADDR_Y_COMPONENT[4]), .I1(TX_ADDR[4]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[4]));   // ../tx.v(82[30:81])
    defparam mux_12_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1767_4_lut (.I0(n205[4]), .I1(ADV_VSYNC_c), .I2(n174[4]), 
            .I3(n4211), .O(n24));   // ../tx.v(72[12] 93[8])
    defparam i1767_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i6_3_lut (.I0(ADDR_Y_COMPONENT[5]), .I1(TX_ADDR[5]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[5]));   // ../tx.v(82[30:81])
    defparam mux_12_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1768_4_lut (.I0(n205[5]), .I1(ADV_VSYNC_c), .I2(n174[5]), 
            .I3(n4211), .O(n23));   // ../tx.v(72[12] 93[8])
    defparam i1768_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i7_3_lut (.I0(ADDR_Y_COMPONENT[6]), .I1(TX_ADDR[6]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[6]));   // ../tx.v(82[30:81])
    defparam mux_12_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR BRAM_ADDR__rep_1_i0 (.Q(\TX_ADDR[11] ), .C(ADV_CLK_c), .E(n2277), 
            .D(BRAM_ADDR_13__N_258[11]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i0 (.Q(Y_DELTA_PATTERN[0]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[1]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS X_DELTA_PATTERN_i0 (.Q(X_DELTA_PATTERN[0]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[1]), .S(n2361));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i0 (.Q(ADDR_Y_COMPONENT[0]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[0]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS X_DELTA_PATTERN_i13 (.Q(X_DELTA_PATTERN[13]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[14]), .S(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR X_DELTA_PATTERN_i12 (.Q(X_DELTA_PATTERN[12]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[13]), .R(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESS X_DELTA_PATTERN_i11 (.Q(X_DELTA_PATTERN[11]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[12]), .S(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR X_DELTA_PATTERN_i10 (.Q(X_DELTA_PATTERN[10]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[11]), .R(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESS X_DELTA_PATTERN_i9 (.Q(X_DELTA_PATTERN[9]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[10]), .S(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR X_DELTA_PATTERN_i8 (.Q(X_DELTA_PATTERN[8]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[9]), .R(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESS X_DELTA_PATTERN_i7 (.Q(X_DELTA_PATTERN[7]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[8]), .S(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESS X_DELTA_PATTERN_i6 (.Q(X_DELTA_PATTERN[6]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[7]), .S(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR X_DELTA_PATTERN_i5 (.Q(X_DELTA_PATTERN[5]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[6]), .R(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i93 (.Q(Y_DELTA_PATTERN[93]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[94]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_LUT4 i1769_4_lut (.I0(n205[6]), .I1(ADV_VSYNC_c), .I2(n174[6]), 
            .I3(n4211), .O(n22));   // ../tx.v(72[12] 93[8])
    defparam i1769_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i8_3_lut (.I0(ADDR_Y_COMPONENT[7]), .I1(TX_ADDR[7]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[7]));   // ../tx.v(82[30:81])
    defparam mux_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1770_4_lut (.I0(n205[7]), .I1(ADV_VSYNC_c), .I2(n174[7]), 
            .I3(n4211), .O(n21));   // ../tx.v(72[12] 93[8])
    defparam i1770_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS X_DELTA_PATTERN_i4 (.Q(X_DELTA_PATTERN[4]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[5]), .S(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR X_DELTA_PATTERN_i3 (.Q(X_DELTA_PATTERN[3]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[4]), .R(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESS X_DELTA_PATTERN_i2 (.Q(X_DELTA_PATTERN[2]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[3]), .S(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR X_DELTA_PATTERN_i1 (.Q(X_DELTA_PATTERN[1]), .C(ADV_CLK_c), 
            .E(n2315), .D(X_DELTA_PATTERN[2]), .R(n4224));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i13 (.Q(ADDR_Y_COMPONENT[13]), .C(ADV_CLK_c), 
            .E(n2305), .D(DEBUG_c_2), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i12 (.Q(ADDR_Y_COMPONENT[12]), .C(ADV_CLK_c), 
            .E(n2305), .D(\TX_ADDR[12] ), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i11 (.Q(ADDR_Y_COMPONENT[11]), .C(ADV_CLK_c), 
            .E(n2305), .D(\TX_ADDR[11] ), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i10 (.Q(ADDR_Y_COMPONENT[10]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[10]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i9 (.Q(ADDR_Y_COMPONENT[9]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[9]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i8 (.Q(ADDR_Y_COMPONENT[8]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[8]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i7 (.Q(ADDR_Y_COMPONENT[7]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[7]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i6 (.Q(ADDR_Y_COMPONENT[6]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[6]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR ADDR_Y_COMPONENT__i5 (.Q(ADDR_Y_COMPONENT[5]), .C(ADV_CLK_c), 
            .E(n2305), .D(TX_ADDR[5]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_LUT4 mux_12_i9_3_lut (.I0(ADDR_Y_COMPONENT[8]), .I1(TX_ADDR[8]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[8]));   // ../tx.v(82[30:81])
    defparam mux_12_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1771_4_lut (.I0(n205[8]), .I1(ADV_VSYNC_c), .I2(n174[8]), 
            .I3(n4211), .O(n20));   // ../tx.v(72[12] 93[8])
    defparam i1771_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i10_3_lut (.I0(ADDR_Y_COMPONENT[9]), .I1(TX_ADDR[9]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[9]));   // ../tx.v(82[30:81])
    defparam mux_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1772_4_lut (.I0(n205[9]), .I1(ADV_VSYNC_c), .I2(n174[9]), 
            .I3(n4211), .O(n19));   // ../tx.v(72[12] 93[8])
    defparam i1772_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS Y_DELTA_PATTERN_i99 (.Q(Y_DELTA_PATTERN[99]), .C(ADV_CLK_c), 
            .E(n4224), .D(Y_DELTA_PATTERN[0]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESR Y_DELTA_PATTERN_i98 (.Q(Y_DELTA_PATTERN[98]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[99]), .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFESS Y_DELTA_PATTERN_i94 (.Q(Y_DELTA_PATTERN[94]), .C(ADV_CLK_c), 
            .E(n2361), .D(Y_DELTA_PATTERN[95]), .S(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    SB_DFFSR BRAM_ADDR__i13 (.Q(DEBUG_c_2), .C(ADV_CLK_c), .D(n2909), 
            .R(ADV_VSYNC_c));   // ../tx.v(72[12] 93[8])
    VGA_CONTROL video_signal_controller (.ADV_CLK_c(ADV_CLK_c), .ADV_HSYNC_c(ADV_HSYNC_c), 
            .ADV_VSYNC_c(ADV_VSYNC_c), .DEBUG_c_6(DEBUG_c_6), .GND_net(GND_net), 
            .n4220(n4220), .n3926(n3926), .\ADDR_Y_COMPONENT[12] (ADDR_Y_COMPONENT[12]), 
            .n190({n190}), .\BRAM_ADDR_13__N_258[12] (BRAM_ADDR_13__N_258[12]), 
            .\Y_DELTA_PATTERN[0] (Y_DELTA_PATTERN[0]), .n2305(n2305), .\ADDR_Y_COMPONENT[11] (ADDR_Y_COMPONENT[11]), 
            .\BRAM_ADDR_13__N_258[11] (BRAM_ADDR_13__N_258[11]), .\ADDR_Y_COMPONENT[13] (ADDR_Y_COMPONENT[13]), 
            .\BRAM_ADDR_13__N_258[13] (BRAM_ADDR_13__N_258[13]), .old_VGA_HS(old_VGA_HS), 
            .n4225(n4225), .n3910(n3910), .\TX_ADDR[8] (TX_ADDR[8]), .n211(n205[8]), 
            .\TX_ADDR[9] (TX_ADDR[9]), .n210(n205[9]), .VCC_net(VCC_net), 
            .n2587(n2587), .\TX_ADDR[10] (TX_ADDR[10]), .n209(n205[10]), 
            .\TX_ADDR[0] (TX_ADDR[0]), .n219(n205[0]), .\TX_ADDR[2] (TX_ADDR[2]), 
            .n217(n205[2]), .n2361(n2361), .\TX_ADDR[1] (TX_ADDR[1]), 
            .n218(n205[1]), .\TX_ADDR[7] (TX_ADDR[7]), .n212(n205[7]), 
            .n4211(n4211), .\TX_ADDR[3] (TX_ADDR[3]), .n216(n205[3]), 
            .\TX_ADDR[4] (TX_ADDR[4]), .n215(n205[4]), .\TX_ADDR[6] (TX_ADDR[6]), 
            .n213(n205[6]), .\TX_ADDR[5] (TX_ADDR[5]), .n214(n205[5]), 
            .n4210(n4210), .n4224(n4224)) /* synthesis syn_module_defined=1 */ ;   // ../tx.v(44[17] 58[67])
    
endmodule
//
// Verilog Description of module VGA_CONTROL
//

module VGA_CONTROL (ADV_CLK_c, ADV_HSYNC_c, ADV_VSYNC_c, DEBUG_c_6, 
            GND_net, n4220, n3926, \ADDR_Y_COMPONENT[12] , n190, \BRAM_ADDR_13__N_258[12] , 
            \Y_DELTA_PATTERN[0] , n2305, \ADDR_Y_COMPONENT[11] , \BRAM_ADDR_13__N_258[11] , 
            \ADDR_Y_COMPONENT[13] , \BRAM_ADDR_13__N_258[13] , old_VGA_HS, 
            n4225, n3910, \TX_ADDR[8] , n211, \TX_ADDR[9] , n210, 
            VCC_net, n2587, \TX_ADDR[10] , n209, \TX_ADDR[0] , n219, 
            \TX_ADDR[2] , n217, n2361, \TX_ADDR[1] , n218, \TX_ADDR[7] , 
            n212, n4211, \TX_ADDR[3] , n216, \TX_ADDR[4] , n215, 
            \TX_ADDR[6] , n213, \TX_ADDR[5] , n214, n4210, n4224) /* synthesis syn_module_defined=1 */ ;
    input ADV_CLK_c;
    output ADV_HSYNC_c;
    output ADV_VSYNC_c;
    input DEBUG_c_6;
    input GND_net;
    output n4220;
    output n3926;
    input \ADDR_Y_COMPONENT[12] ;
    input [13:0]n190;
    output \BRAM_ADDR_13__N_258[12] ;
    input \Y_DELTA_PATTERN[0] ;
    output n2305;
    input \ADDR_Y_COMPONENT[11] ;
    output \BRAM_ADDR_13__N_258[11] ;
    input \ADDR_Y_COMPONENT[13] ;
    output \BRAM_ADDR_13__N_258[13] ;
    input old_VGA_HS;
    output n4225;
    output n3910;
    input \TX_ADDR[8] ;
    output n211;
    input \TX_ADDR[9] ;
    output n210;
    input VCC_net;
    output n2587;
    input \TX_ADDR[10] ;
    output n209;
    input \TX_ADDR[0] ;
    output n219;
    input \TX_ADDR[2] ;
    output n217;
    output n2361;
    input \TX_ADDR[1] ;
    output n218;
    input \TX_ADDR[7] ;
    output n212;
    output n4211;
    input \TX_ADDR[3] ;
    output n216;
    input \TX_ADDR[4] ;
    output n215;
    input \TX_ADDR[6] ;
    output n213;
    input \TX_ADDR[5] ;
    output n214;
    output n4210;
    output n4224;
    
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    
    wire SYNC_BUFF1, SYNC_BUFF2, VGA_HS_N_545, VGA_VS_N_548;
    wire [11:0]n532;
    wire [11:0]VGA_X;   // ../vga_control.v(54[16:21])
    
    wire n2274, n3698, n3697, n3696;
    wire [11:0]n546;
    wire [11:0]VGA_Y;   // ../vga_control.v(54[23:28])
    
    wire n3686, n3695, n3694, n3693, n3917, n3196, n2260, n3226, 
        n3682, n2594, n2219, n4217, n18, n3935, n3687, n3683, 
        n3685, n3692, n3689, n3677, n3691, n3690, n3688, n3681, 
        n3678, n3680, n3684, n3679, n6, n3892, n3987, n4218, 
        n4, n3936, n4215, VGA_VISIBLE_Y_N_553, n3997, n3978, n4216, 
        n4052, n12;
    
    SB_DFF SYNC_BUFF2_58 (.Q(SYNC_BUFF2), .C(ADV_CLK_c), .D(SYNC_BUFF1));   // ../vga_control.v(74[12] 103[8])
    SB_DFF VGA_HS_60 (.Q(ADV_HSYNC_c), .C(ADV_CLK_c), .D(VGA_HS_N_545));   // ../vga_control.v(74[12] 103[8])
    SB_DFF VGA_VS_61 (.Q(ADV_VSYNC_c), .C(ADV_CLK_c), .D(VGA_VS_N_548));   // ../vga_control.v(74[12] 103[8])
    SB_DFF SYNC_BUFF1_57 (.Q(SYNC_BUFF1), .C(ADV_CLK_c), .D(DEBUG_c_6));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i0 (.Q(VGA_X[0]), .C(ADV_CLK_c), .D(n532[0]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_LUT4 add_83_13_lut (.I0(GND_net), .I1(VGA_X[11]), .I2(GND_net), 
            .I3(n3698), .O(n532[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR VGA_X_i1 (.Q(VGA_X[1]), .C(ADV_CLK_c), .D(n532[1]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i2 (.Q(VGA_X[2]), .C(ADV_CLK_c), .D(n532[2]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i3 (.Q(VGA_X[3]), .C(ADV_CLK_c), .D(n532[3]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i4 (.Q(VGA_X[4]), .C(ADV_CLK_c), .D(n532[4]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i5 (.Q(VGA_X[5]), .C(ADV_CLK_c), .D(n532[5]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i6 (.Q(VGA_X[6]), .C(ADV_CLK_c), .D(n532[6]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i7 (.Q(VGA_X[7]), .C(ADV_CLK_c), .D(n532[7]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i8 (.Q(VGA_X[8]), .C(ADV_CLK_c), .D(n532[8]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i9 (.Q(VGA_X[9]), .C(ADV_CLK_c), .D(n532[9]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i10 (.Q(VGA_X[10]), .C(ADV_CLK_c), .D(n532[10]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_DFFSR VGA_X_i11 (.Q(VGA_X[11]), .C(ADV_CLK_c), .D(n532[11]), .R(n2274));   // ../vga_control.v(74[12] 103[8])
    SB_LUT4 add_83_12_lut (.I0(GND_net), .I1(VGA_X[10]), .I2(GND_net), 
            .I3(n3697), .O(n532[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_83_12 (.CI(n3697), .I0(VGA_X[10]), .I1(GND_net), .CO(n3698));
    SB_LUT4 add_83_11_lut (.I0(GND_net), .I1(VGA_X[9]), .I2(GND_net), 
            .I3(n3696), .O(n532[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_83_11 (.CI(n3696), .I0(VGA_X[9]), .I1(GND_net), .CO(n3697));
    SB_LUT4 add_84_12_lut (.I0(GND_net), .I1(VGA_Y[10]), .I2(GND_net), 
            .I3(n3686), .O(n546[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_83_10_lut (.I0(GND_net), .I1(VGA_X[8]), .I2(GND_net), 
            .I3(n3695), .O(n532[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_18_i13_3_lut_4_lut (.I0(n4220), .I1(n3926), .I2(\ADDR_Y_COMPONENT[12] ), 
            .I3(n190[12]), .O(\BRAM_ADDR_13__N_258[12] ));   // ../vga_control.v(57[28:103])
    defparam mux_18_i13_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY add_83_10 (.CI(n3695), .I0(VGA_X[8]), .I1(GND_net), .CO(n3696));
    SB_LUT4 add_83_9_lut (.I0(GND_net), .I1(VGA_X[7]), .I2(GND_net), .I3(n3694), 
            .O(n532[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_83_9 (.CI(n3694), .I0(VGA_X[7]), .I1(GND_net), .CO(n3695));
    SB_LUT4 add_83_8_lut (.I0(GND_net), .I1(VGA_X[6]), .I2(GND_net), .I3(n3693), 
            .O(n532[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(n4220), .I1(n3926), .I2(\Y_DELTA_PATTERN[0] ), 
            .I3(ADV_VSYNC_c), .O(n2305));   // ../vga_control.v(57[28:103])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff80;
    SB_LUT4 i1_2_lut (.I0(VGA_X[4]), .I1(VGA_X[3]), .I2(GND_net), .I3(GND_net), 
            .O(n3917));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1853_4_lut (.I0(n3196), .I1(VGA_X[8]), .I2(n2260), .I3(n3917), 
            .O(n3226));
    defparam i1853_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 mux_18_i12_3_lut_4_lut (.I0(n4220), .I1(n3926), .I2(\ADDR_Y_COMPONENT[11] ), 
            .I3(n190[11]), .O(\BRAM_ADDR_13__N_258[11] ));   // ../vga_control.v(57[28:103])
    defparam mux_18_i12_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 add_84_8_lut (.I0(GND_net), .I1(VGA_Y[6]), .I2(GND_net), .I3(n3682), 
            .O(n546[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR VGA_Y_i6 (.Q(VGA_Y[6]), .C(ADV_CLK_c), .E(n2274), .D(n546[6]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_LUT4 i2_3_lut (.I0(VGA_X[11]), .I1(VGA_X[10]), .I2(VGA_X[9]), .I3(GND_net), 
            .O(n2219));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_18_i14_3_lut_4_lut (.I0(n4220), .I1(n3926), .I2(\ADDR_Y_COMPONENT[13] ), 
            .I3(n190[13]), .O(\BRAM_ADDR_13__N_258[13] ));   // ../vga_control.v(57[28:103])
    defparam mux_18_i14_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1859_4_lut (.I0(n3226), .I1(VGA_X[11]), .I2(VGA_X[10]), .I3(VGA_X[9]), 
            .O(n2274));
    defparam i1859_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i557_4_lut (.I0(n4217), .I1(VGA_X[8]), .I2(n2260), .I3(n3917), 
            .O(n18));
    defparam i557_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i143_2_lut_3_lut_4_lut_rep_34 (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), 
            .I2(ADV_VSYNC_c), .I3(n3926), .O(n4225));   // ../vga_control.v(57[28:103])
    defparam i143_2_lut_3_lut_4_lut_rep_34.LUT_INIT = 16'hf4f0;
    SB_LUT4 mux_14_i9_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[8]), 
            .I3(\TX_ADDR[8] ), .O(n211));   // ../vga_control.v(57[28:103])
    defparam mux_14_i9_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_14_i10_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[9]), 
            .I3(\TX_ADDR[9] ), .O(n210));   // ../vga_control.v(57[28:103])
    defparam mux_14_i10_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESR VGA_Y_i11 (.Q(VGA_Y[11]), .C(ADV_CLK_c), .E(n2274), .D(n546[11]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_DFFESR VGA_Y_i10 (.Q(VGA_Y[10]), .C(ADV_CLK_c), .E(n2274), .D(n546[10]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_DFFESR VGA_Y_i9 (.Q(VGA_Y[9]), .C(ADV_CLK_c), .E(n2274), .D(n546[9]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_DFFESR VGA_Y_i8 (.Q(VGA_Y[8]), .C(ADV_CLK_c), .E(n2274), .D(n546[8]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_DFFESR VGA_Y_i7 (.Q(VGA_Y[7]), .C(ADV_CLK_c), .E(n2274), .D(n546[7]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_LUT4 i1_2_lut_adj_12 (.I0(VGA_Y[7]), .I1(VGA_Y[8]), .I2(GND_net), 
            .I3(GND_net), .O(n3935));   // ../vga_control.v(54[23:28])
    defparam i1_2_lut_adj_12.LUT_INIT = 16'heeee;
    SB_CARRY add_84_12 (.CI(n3686), .I0(VGA_Y[10]), .I1(GND_net), .CO(n3687));
    SB_CARRY add_84_8 (.CI(n3682), .I0(VGA_Y[6]), .I1(GND_net), .CO(n3683));
    SB_CARRY add_83_8 (.CI(n3693), .I0(VGA_X[6]), .I1(GND_net), .CO(n3694));
    SB_LUT4 add_84_11_lut (.I0(GND_net), .I1(VGA_Y[9]), .I2(GND_net), 
            .I3(n3685), .O(n546[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_83_7_lut (.I0(GND_net), .I1(VGA_X[5]), .I2(GND_net), .I3(n3692), 
            .O(n532[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_83_4_lut (.I0(GND_net), .I1(VGA_X[2]), .I2(GND_net), .I3(n3689), 
            .O(n532[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_83_7 (.CI(n3692), .I0(VGA_X[5]), .I1(GND_net), .CO(n3693));
    SB_LUT4 add_84_3_lut (.I0(GND_net), .I1(VGA_Y[1]), .I2(GND_net), .I3(n3677), 
            .O(n546[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_83_6_lut (.I0(GND_net), .I1(VGA_X[4]), .I2(GND_net), .I3(n3691), 
            .O(n532[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_83_4 (.CI(n3689), .I0(VGA_X[2]), .I1(GND_net), .CO(n3690));
    SB_LUT4 add_83_3_lut (.I0(GND_net), .I1(VGA_X[1]), .I2(GND_net), .I3(n3688), 
            .O(n532[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_83_6 (.CI(n3691), .I0(VGA_X[4]), .I1(GND_net), .CO(n3692));
    SB_LUT4 add_84_7_lut (.I0(GND_net), .I1(VGA_Y[5]), .I2(GND_net), .I3(n3681), 
            .O(n546[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_84_7 (.CI(n3681), .I0(VGA_Y[5]), .I1(GND_net), .CO(n3682));
    SB_CARRY add_84_3 (.CI(n3677), .I0(VGA_Y[1]), .I1(GND_net), .CO(n3678));
    SB_LUT4 add_84_6_lut (.I0(GND_net), .I1(VGA_Y[4]), .I2(GND_net), .I3(n3680), 
            .O(n546[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_84_11 (.CI(n3685), .I0(VGA_Y[9]), .I1(GND_net), .CO(n3686));
    SB_LUT4 add_84_2_lut (.I0(GND_net), .I1(VGA_Y[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n546[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_84_2 (.CI(VCC_net), .I0(VGA_Y[0]), .I1(GND_net), .CO(n3677));
    SB_LUT4 add_84_10_lut (.I0(GND_net), .I1(VGA_Y[8]), .I2(GND_net), 
            .I3(n3684), .O(n546[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_83_3 (.CI(n3688), .I0(VGA_X[1]), .I1(GND_net), .CO(n3689));
    SB_LUT4 add_83_5_lut (.I0(GND_net), .I1(VGA_X[3]), .I2(GND_net), .I3(n3690), 
            .O(n532[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_83_2_lut (.I0(GND_net), .I1(VGA_X[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n532[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_83_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1227_2_lut (.I0(n2274), .I1(SYNC_BUFF2), .I2(GND_net), .I3(GND_net), 
            .O(n2594));   // ../vga_control.v(74[12] 103[8])
    defparam i1227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1211_1_lut_2_lut (.I0(n3910), .I1(n3926), .I2(GND_net), .I3(GND_net), 
            .O(n2587));   // ../vga_control.v(57[28:103])
    defparam i1211_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 mux_14_i11_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[10]), 
            .I3(\TX_ADDR[10] ), .O(n209));   // ../vga_control.v(57[28:103])
    defparam mux_14_i11_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY add_84_6 (.CI(n3680), .I0(VGA_Y[4]), .I1(GND_net), .CO(n3681));
    SB_LUT4 add_84_5_lut (.I0(GND_net), .I1(VGA_Y[3]), .I2(GND_net), .I3(n3679), 
            .O(n546[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_84_5 (.CI(n3679), .I0(VGA_Y[3]), .I1(GND_net), .CO(n3680));
    SB_CARRY add_84_10 (.CI(n3684), .I0(VGA_Y[8]), .I1(GND_net), .CO(n3685));
    SB_CARRY add_83_2 (.CI(VCC_net), .I0(VGA_X[0]), .I1(GND_net), .CO(n3688));
    SB_LUT4 add_84_4_lut (.I0(GND_net), .I1(VGA_Y[2]), .I2(GND_net), .I3(n3678), 
            .O(n546[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_84_9_lut (.I0(GND_net), .I1(VGA_Y[7]), .I2(GND_net), .I3(n3683), 
            .O(n546[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_84_4 (.CI(n3678), .I0(VGA_Y[2]), .I1(GND_net), .CO(n3679));
    SB_CARRY add_84_9 (.CI(n3683), .I0(VGA_Y[7]), .I1(GND_net), .CO(n3684));
    SB_LUT4 add_84_13_lut (.I0(GND_net), .I1(VGA_Y[11]), .I2(GND_net), 
            .I3(n3687), .O(n546[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_84_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_83_5 (.CI(n3690), .I0(VGA_X[3]), .I1(GND_net), .CO(n3691));
    SB_LUT4 mux_14_i1_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[0]), 
            .I3(\TX_ADDR[0] ), .O(n219));   // ../vga_control.v(57[28:103])
    defparam mux_14_i1_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_14_i3_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[2]), 
            .I3(\TX_ADDR[2] ), .O(n217));   // ../vga_control.v(57[28:103])
    defparam mux_14_i3_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut (.I0(VGA_Y[5]), .I1(VGA_Y[9]), .I2(n3935), .I3(n6), 
            .O(n3892));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut (.I0(VGA_Y[4]), .I1(n3892), .I2(VGA_Y[3]), .I3(VGA_Y[2]), 
            .O(n3987));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR VGA_Y_i5 (.Q(VGA_Y[5]), .C(ADV_CLK_c), .E(n2274), .D(n546[5]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_LUT4 i143_2_lut_3_lut_4_lut (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), .I2(ADV_VSYNC_c), 
            .I3(n3926), .O(n2361));   // ../vga_control.v(57[28:103])
    defparam i143_2_lut_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_LUT4 mux_14_i2_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[1]), 
            .I3(\TX_ADDR[1] ), .O(n218));   // ../vga_control.v(57[28:103])
    defparam mux_14_i2_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_14_i8_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[7]), 
            .I3(\TX_ADDR[7] ), .O(n212));   // ../vga_control.v(57[28:103])
    defparam mux_14_i8_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_rep_20_3_lut (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), .I2(n3926), 
            .I3(GND_net), .O(n4211));   // ../vga_control.v(57[28:103])
    defparam i1_2_lut_rep_20_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_rep_29 (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), .I2(GND_net), 
            .I3(GND_net), .O(n4220));   // ../vga_control.v(57[28:103])
    defparam i1_2_lut_rep_29.LUT_INIT = 16'h4444;
    SB_DFFESR VGA_Y_i4 (.Q(VGA_Y[4]), .C(ADV_CLK_c), .E(n2274), .D(n546[4]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_DFFESR VGA_Y_i3 (.Q(VGA_Y[3]), .C(ADV_CLK_c), .E(n2274), .D(n546[3]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_DFFESR VGA_Y_i2 (.Q(VGA_Y[2]), .C(ADV_CLK_c), .E(n2274), .D(n546[2]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_DFFESR VGA_Y_i1 (.Q(VGA_Y[1]), .C(ADV_CLK_c), .E(n2274), .D(n546[1]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_DFFESR VGA_Y_i0 (.Q(VGA_Y[0]), .C(ADV_CLK_c), .E(n2274), .D(n546[0]), 
            .R(n2594));   // ../vga_control.v(74[12] 103[8])
    SB_LUT4 i1_2_lut_3_lut (.I0(VGA_Y[10]), .I1(VGA_Y[11]), .I2(VGA_Y[6]), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_rep_27 (.I0(VGA_Y[10]), .I1(VGA_Y[11]), .I2(GND_net), 
            .I3(GND_net), .O(n4218));
    defparam i1_2_lut_rep_27.LUT_INIT = 16'heeee;
    SB_LUT4 i2636_3_lut (.I0(n3987), .I1(VGA_Y[1]), .I2(VGA_Y[0]), .I3(GND_net), 
            .O(VGA_VS_N_548));   // ../vga_control.v(74[12] 103[8])
    defparam i2636_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 mux_14_i4_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[3]), 
            .I3(\TX_ADDR[3] ), .O(n216));   // ../vga_control.v(57[28:103])
    defparam mux_14_i4_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut (.I0(VGA_Y[6]), .I1(n3935), .I2(VGA_Y[5]), .I3(n4), 
            .O(n3936));   // ../vga_control.v(54[23:28])
    defparam i1_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_13 (.I0(VGA_Y[4]), .I1(n3892), .I2(VGA_Y[3]), 
            .I3(n4215), .O(VGA_VISIBLE_Y_N_553));
    defparam i1_4_lut_adj_13.LUT_INIT = 16'heeec;
    SB_LUT4 i2_4_lut (.I0(VGA_X[2]), .I1(VGA_X[3]), .I2(VGA_X[0]), .I3(VGA_X[1]), 
            .O(n3997));
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 mux_14_i5_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[4]), 
            .I3(\TX_ADDR[4] ), .O(n215));   // ../vga_control.v(57[28:103])
    defparam mux_14_i5_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_14_i7_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[6]), 
            .I3(\TX_ADDR[6] ), .O(n213));   // ../vga_control.v(57[28:103])
    defparam mux_14_i7_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_14 (.I0(n3997), .I1(VGA_X[5]), .I2(VGA_X[4]), 
            .I3(VGA_X[6]), .O(n3978));
    defparam i3_4_lut_adj_14.LUT_INIT = 16'hfffe;
    SB_LUT4 i1823_2_lut_3_lut (.I0(VGA_X[1]), .I1(VGA_X[2]), .I2(VGA_X[0]), 
            .I3(GND_net), .O(n3196));
    defparam i1823_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i560_2_lut_rep_26 (.I0(VGA_X[1]), .I1(VGA_X[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4217));
    defparam i560_2_lut_rep_26.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_15 (.I0(VGA_X[7]), .I1(VGA_X[6]), .I2(VGA_X[5]), 
            .I3(GND_net), .O(n2260));
    defparam i1_2_lut_3_lut_adj_15.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_rep_25 (.I0(VGA_X[7]), .I1(VGA_X[6]), .I2(GND_net), 
            .I3(GND_net), .O(n4216));
    defparam i1_2_lut_rep_25.LUT_INIT = 16'heeee;
    SB_LUT4 i2578_3_lut (.I0(n3978), .I1(n2219), .I2(VGA_X[7]), .I3(GND_net), 
            .O(n4052));
    defparam i2578_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2_4_lut_adj_16 (.I0(n4218), .I1(VGA_VISIBLE_Y_N_553), .I2(VGA_Y[9]), 
            .I3(n3936), .O(n3926));
    defparam i2_4_lut_adj_16.LUT_INIT = 16'h0444;
    SB_LUT4 mux_14_i6_3_lut_4_lut (.I0(n3910), .I1(n3926), .I2(n190[5]), 
            .I3(\TX_ADDR[5] ), .O(n214));   // ../vga_control.v(57[28:103])
    defparam mux_14_i6_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i570_3_lut (.I0(VGA_X[3]), .I1(VGA_X[5]), .I2(VGA_X[4]), .I3(GND_net), 
            .O(n12));
    defparam i570_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_rep_19 (.I0(n3910), .I1(n3926), .I2(GND_net), .I3(GND_net), 
            .O(n4210));   // ../vga_control.v(57[28:103])
    defparam i1_2_lut_rep_19.LUT_INIT = 16'h8888;
    SB_LUT4 i143_2_lut_3_lut_4_lut_rep_33 (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), 
            .I2(ADV_VSYNC_c), .I3(n3926), .O(n4224));   // ../vga_control.v(57[28:103])
    defparam i143_2_lut_3_lut_4_lut_rep_33.LUT_INIT = 16'hf4f0;
    SB_LUT4 i1_3_lut_4_lut_adj_17 (.I0(VGA_Y[2]), .I1(VGA_Y[1]), .I2(VGA_Y[3]), 
            .I3(VGA_Y[4]), .O(n4));   // ../vga_control.v(54[23:28])
    defparam i1_3_lut_4_lut_adj_17.LUT_INIT = 16'hff80;
    SB_LUT4 i2631_4_lut (.I0(n12), .I1(n4052), .I2(VGA_X[8]), .I3(n4216), 
            .O(VGA_HS_N_545));   // ../vga_control.v(80[19:88])
    defparam i2631_4_lut.LUT_INIT = 16'hfcfd;
    SB_LUT4 i1_2_lut_rep_24 (.I0(VGA_Y[2]), .I1(VGA_Y[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4215));   // ../vga_control.v(54[23:28])
    defparam i1_2_lut_rep_24.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_4_lut (.I0(VGA_X[11]), .I1(n18), .I2(VGA_X[10]), 
            .I3(VGA_X[9]), .O(n3910));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h0514;
    
endmodule
//
// Verilog Description of module DIV_BY_5
//

module DIV_BY_5 (DEBUG_c_1_c, GND_net, DEBUG_c_0) /* synthesis syn_module_defined=1 */ ;
    input DEBUG_c_1_c;
    input GND_net;
    output DEBUG_c_0;
    
    wire DEBUG_c_1_c /* synthesis SET_AS_NETWORK=DEBUG_c_1_c, is_clock=1 */ ;   // ../main.v(2[19:24])
    wire [3:0]NEXT_COUNTER;   // ../div_by_5.v(3[12:24])
    wire [3:0]COUNTER;   // ../div_by_5.v(2[12:19])
    wire [31:0]NEXT_COUNTER_3__N_9;
    
    wire n4221, CLK_EN_N_14;
    
    SB_DFF COUNTER_i0 (.Q(COUNTER[0]), .C(DEBUG_c_1_c), .D(NEXT_COUNTER[0]));   // ../div_by_5.v(4[9] 7[5])
    SB_LUT4 i455_2_lut (.I0(COUNTER[1]), .I1(COUNTER[0]), .I2(GND_net), 
            .I3(GND_net), .O(NEXT_COUNTER_3__N_9[1]));   // ../div_by_5.v(11[20:31])
    defparam i455_2_lut.LUT_INIT = 16'h6666;
    SB_DFFNSR NEXT_COUNTER__i0 (.Q(NEXT_COUNTER[0]), .C(DEBUG_c_1_c), .D(NEXT_COUNTER_3__N_9[0]), 
            .R(n4221));   // ../div_by_5.v(9[9] 15[5])
    SB_DFF COUNTER_i3 (.Q(COUNTER[3]), .C(DEBUG_c_1_c), .D(NEXT_COUNTER[3]));   // ../div_by_5.v(4[9] 7[5])
    SB_DFF COUNTER_i2 (.Q(COUNTER[2]), .C(DEBUG_c_1_c), .D(NEXT_COUNTER[2]));   // ../div_by_5.v(4[9] 7[5])
    SB_DFF COUNTER_i1 (.Q(COUNTER[1]), .C(DEBUG_c_1_c), .D(NEXT_COUNTER[1]));   // ../div_by_5.v(4[9] 7[5])
    SB_DFFNSR NEXT_COUNTER__i3 (.Q(NEXT_COUNTER[3]), .C(DEBUG_c_1_c), .D(NEXT_COUNTER_3__N_9[3]), 
            .R(n4221));   // ../div_by_5.v(9[9] 15[5])
    SB_DFFNSR NEXT_COUNTER__i2 (.Q(NEXT_COUNTER[2]), .C(DEBUG_c_1_c), .D(NEXT_COUNTER_3__N_9[2]), 
            .R(n4221));   // ../div_by_5.v(9[9] 15[5])
    SB_LUT4 i2639_3_lut_4_lut (.I0(NEXT_COUNTER[3]), .I1(NEXT_COUNTER[2]), 
            .I2(NEXT_COUNTER[0]), .I3(NEXT_COUNTER[1]), .O(CLK_EN_N_14));   // ../div_by_5.v(9[9] 15[5])
    defparam i2639_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_2_lut_rep_30 (.I0(NEXT_COUNTER[3]), .I1(NEXT_COUNTER[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4221));   // ../div_by_5.v(9[9] 15[5])
    defparam i2_2_lut_rep_30.LUT_INIT = 16'heeee;
    SB_DFFNSR NEXT_COUNTER__i1 (.Q(NEXT_COUNTER[1]), .C(DEBUG_c_1_c), .D(NEXT_COUNTER_3__N_9[1]), 
            .R(n4221));   // ../div_by_5.v(9[9] 15[5])
    SB_DFF CLK_EN_13 (.Q(DEBUG_c_0), .C(DEBUG_c_1_c), .D(CLK_EN_N_14));   // ../div_by_5.v(4[9] 7[5])
    SB_LUT4 i462_2_lut_3_lut (.I0(COUNTER[1]), .I1(COUNTER[0]), .I2(COUNTER[2]), 
            .I3(GND_net), .O(NEXT_COUNTER_3__N_9[2]));   // ../div_by_5.v(11[20:31])
    defparam i462_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i469_3_lut_4_lut (.I0(COUNTER[1]), .I1(COUNTER[0]), .I2(COUNTER[2]), 
            .I3(COUNTER[3]), .O(NEXT_COUNTER_3__N_9[3]));   // ../div_by_5.v(11[20:31])
    defparam i469_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i453_1_lut (.I0(COUNTER[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(NEXT_COUNTER_3__N_9[0]));   // ../div_by_5.v(11[20:31])
    defparam i453_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module TX_PLL
//

module TX_PLL (DEBUG_c_1_c, VCC_net, GND_net, ADV_CLK_c) /* synthesis syn_module_defined=1 */ ;
    input DEBUG_c_1_c;
    input VCC_net;
    input GND_net;
    output ADV_CLK_c;
    
    wire DEBUG_c_1_c /* synthesis SET_AS_NETWORK=DEBUG_c_1_c, is_clock=1 */ ;   // ../main.v(2[19:24])
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    
    SB_PLL40_CORE TX_PLL_inst (.REFERENCECLK(DEBUG_c_1_c), .PLLOUTCORE(ADV_CLK_c), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=17, LSE_LCOL=9, LSE_RCOL=27, LSE_LLINE=21, LSE_RLINE=25 */ ;   // ../main.v(21[9] 25[27])
    defparam TX_PLL_inst.FEEDBACK_PATH = "SIMPLE";
    defparam TX_PLL_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam TX_PLL_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam TX_PLL_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam TX_PLL_inst.FDA_FEEDBACK = 4'b0000;
    defparam TX_PLL_inst.FDA_RELATIVE = 4'b0000;
    defparam TX_PLL_inst.PLLOUT_SELECT = "GENCLK";
    defparam TX_PLL_inst.DIVR = 4'b0000;
    defparam TX_PLL_inst.DIVF = 7'b0100110;
    defparam TX_PLL_inst.DIVQ = 3'b100;
    defparam TX_PLL_inst.FILTER_RANGE = 3'b010;
    defparam TX_PLL_inst.ENABLE_ICEGATE = 1'b0;
    defparam TX_PLL_inst.TEST_MODE = 1'b0;
    defparam TX_PLL_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module RAM
//

module RAM (TX_DATA, ADV_CLK_c, \TX_ADDR[11] , \TX_ADDR[12] , GND_net, 
            DEBUG_c_2, \RX_ADDR[11] , \RX_ADDR[12] , DEBUG_c_5, DEBUG_c_3, 
            \RX_ADDR[0] , \RX_ADDR[1] , \RX_ADDR[2] , \RX_ADDR[3] , 
            \RX_ADDR[4] , \RX_ADDR[5] , \RX_ADDR[6] , \RX_ADDR[7] , 
            \RX_ADDR[8] , \RX_ADDR[9] , \RX_ADDR[10] , n28, n27, n26, 
            n25, n24, n23, n22, n21, n20, n19, n18, TVP_VIDEO_c_8, 
            TVP_VIDEO_c_9, DEBUG_c_1_c, VCC_net, TVP_VIDEO_c_6, TVP_VIDEO_c_7, 
            TVP_VIDEO_c_4, TVP_VIDEO_c_5, TVP_VIDEO_c_2, TVP_VIDEO_c_3, 
            n658, n690, n659, n691) /* synthesis syn_module_defined=1 */ ;
    output [7:0]TX_DATA;
    input ADV_CLK_c;
    input \TX_ADDR[11] ;
    input \TX_ADDR[12] ;
    input GND_net;
    input DEBUG_c_2;
    input \RX_ADDR[11] ;
    input \RX_ADDR[12] ;
    input DEBUG_c_5;
    input DEBUG_c_3;
    input \RX_ADDR[0] ;
    input \RX_ADDR[1] ;
    input \RX_ADDR[2] ;
    input \RX_ADDR[3] ;
    input \RX_ADDR[4] ;
    input \RX_ADDR[5] ;
    input \RX_ADDR[6] ;
    input \RX_ADDR[7] ;
    input \RX_ADDR[8] ;
    input \RX_ADDR[9] ;
    input \RX_ADDR[10] ;
    input n28;
    input n27;
    input n26;
    input n25;
    input n24;
    input n23;
    input n22;
    input n21;
    input n20;
    input n19;
    input n18;
    input TVP_VIDEO_c_8;
    input TVP_VIDEO_c_9;
    input DEBUG_c_1_c;
    input VCC_net;
    input TVP_VIDEO_c_6;
    input TVP_VIDEO_c_7;
    input TVP_VIDEO_c_4;
    input TVP_VIDEO_c_5;
    input TVP_VIDEO_c_2;
    input TVP_VIDEO_c_3;
    input n658;
    input n690;
    input n659;
    input n691;
    
    wire ADV_CLK_c /* synthesis is_clock=1, SET_AS_NETWORK=ADV_CLK_c */ ;   // ../main.v(13[14:21])
    wire DEBUG_c_1_c /* synthesis SET_AS_NETWORK=DEBUG_c_1_c, is_clock=1 */ ;   // ../main.v(2[19:24])
    wire [7:0]dout_7__N_567;
    
    wire n675, n683, n4170, n619, n611, n4173, n547, n555, n4074, 
        n642, n650, n4164, n553, n545, n4167, n644, n652, n4075, 
        n674, n682, n4158, n618, n610, n4161, n677, n685, n4063, 
        n4065, n4066, n4128, n643, n651, n4152, n554, n546, 
        n4155, n613, n621, n4062, n673, n681, n4146, n617, n609, 
        n4149, n4185, n4125, n4140, n4179, n4191, n4078, n4077, 
        n4119, n4071, n4072, n4134, n562, n627, n4102, n4101, 
        n615, n616, n626, n548, n549, n561, n544, n614, n647, 
        n648, n612, n645, n646, n558, n559, n680, n688, n4122, 
        n641, n556, n557, n679, n552, n678, n623, n624, n676, 
        n622, n655, n656, n620, n653, n654, n687, n649, n686, 
        n550, n551, n684, n4116, n4188, n4182, n4176;
    
    SB_DFF dout_i0 (.Q(TX_DATA[0]), .C(ADV_CLK_c), .D(dout_7__N_567[0]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2693 (.I0(\TX_ADDR[11] ), .I1(n675), .I2(n683), 
            .I3(\TX_ADDR[12] ), .O(n4170));
    defparam TX_ADDR_11__bdd_4_lut_2693.LUT_INIT = 16'he4aa;
    SB_LUT4 n4170_bdd_4_lut (.I0(n4170), .I1(n619), .I2(n611), .I3(\TX_ADDR[12] ), 
            .O(n4173));
    defparam n4170_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2600_3_lut (.I0(n547), .I1(n555), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4074));
    defparam i2600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2688 (.I0(\TX_ADDR[11] ), .I1(n642), .I2(n650), 
            .I3(\TX_ADDR[12] ), .O(n4164));
    defparam TX_ADDR_11__bdd_4_lut_2688.LUT_INIT = 16'he4aa;
    SB_LUT4 n4164_bdd_4_lut (.I0(n4164), .I1(n553), .I2(n545), .I3(\TX_ADDR[12] ), 
            .O(n4167));
    defparam n4164_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2601_3_lut (.I0(n644), .I1(n652), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4075));
    defparam i2601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2683 (.I0(\TX_ADDR[11] ), .I1(n674), .I2(n682), 
            .I3(\TX_ADDR[12] ), .O(n4158));
    defparam TX_ADDR_11__bdd_4_lut_2683.LUT_INIT = 16'he4aa;
    SB_LUT4 n4158_bdd_4_lut (.I0(n4158), .I1(n618), .I2(n610), .I3(\TX_ADDR[12] ), 
            .O(n4161));
    defparam n4158_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2589_3_lut (.I0(n677), .I1(n685), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4063));
    defparam i2589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_12__bdd_4_lut_2658 (.I0(\TX_ADDR[12] ), .I1(n4065), 
            .I2(n4066), .I3(DEBUG_c_2), .O(n4128));
    defparam TX_ADDR_12__bdd_4_lut_2658.LUT_INIT = 16'he4aa;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2678 (.I0(\TX_ADDR[11] ), .I1(n643), .I2(n651), 
            .I3(\TX_ADDR[12] ), .O(n4152));
    defparam TX_ADDR_11__bdd_4_lut_2678.LUT_INIT = 16'he4aa;
    SB_LUT4 n4152_bdd_4_lut (.I0(n4152), .I1(n554), .I2(n546), .I3(\TX_ADDR[12] ), 
            .O(n4155));
    defparam n4152_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2588_3_lut (.I0(n613), .I1(n621), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4062));
    defparam i2588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2673 (.I0(\TX_ADDR[11] ), .I1(n673), .I2(n681), 
            .I3(\TX_ADDR[12] ), .O(n4146));
    defparam TX_ADDR_11__bdd_4_lut_2673.LUT_INIT = 16'he4aa;
    SB_LUT4 n4146_bdd_4_lut (.I0(n4146), .I1(n617), .I2(n609), .I3(\TX_ADDR[12] ), 
            .O(n4149));
    defparam n4146_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i191932_i1_3_lut (.I0(n4185), .I1(n4125), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_567[7]));
    defparam i191932_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_12__bdd_4_lut (.I0(\TX_ADDR[12] ), .I1(n4062), .I2(n4063), 
            .I3(DEBUG_c_2), .O(n4140));
    defparam TX_ADDR_12__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i190726_i1_3_lut (.I0(n4179), .I1(n4191), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_567[5]));
    defparam i190726_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i188917_i1_3_lut (.I0(n4155), .I1(n4173), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_567[2]));
    defparam i188917_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n4128_bdd_4_lut (.I0(n4128), .I1(n4075), .I2(n4074), .I3(DEBUG_c_2), 
            .O(dout_7__N_567[3]));
    defparam n4128_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i188314_i1_3_lut (.I0(n4167), .I1(n4161), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_567[1]));
    defparam i188314_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n4140_bdd_4_lut (.I0(n4140), .I1(n4078), .I2(n4077), .I3(DEBUG_c_2), 
            .O(dout_7__N_567[4]));
    defparam n4140_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i187711_i1_3_lut (.I0(n4119), .I1(n4149), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_567[0]));
    defparam i187711_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_12__bdd_4_lut_2663 (.I0(\TX_ADDR[12] ), .I1(n4071), 
            .I2(n4072), .I3(DEBUG_c_2), .O(n4134));
    defparam TX_ADDR_12__bdd_4_lut_2663.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_4_lut (.I0(\RX_ADDR[11] ), .I1(\RX_ADDR[12] ), .I2(DEBUG_c_5), 
            .I3(DEBUG_c_3), .O(n562));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\RX_ADDR[11] ), .I1(\RX_ADDR[12] ), 
            .I2(DEBUG_c_5), .I3(DEBUG_c_3), .O(n627));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 n4134_bdd_4_lut (.I0(n4134), .I1(n4102), .I2(n4101), .I3(DEBUG_c_2), 
            .O(dout_7__N_567[6]));
    defparam n4134_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_RAM2048x2 mem0 (.RDATA({n616, n615}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n626), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem0.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem8 (.RDATA({n549, n548}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n561), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem8.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem9 (.RDATA({n547, n546}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n561), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem9.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem10 (.RDATA({n545, n544}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n561), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem10.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem11 (.RDATA({n614, n613}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n626), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem11.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem1 (.RDATA({n648, n647}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n658), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem1.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem12 (.RDATA({n612, n611}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n626), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem13 (.RDATA({n610, n609}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n626), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem13.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem14 (.RDATA({n646, n645}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n658), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem14.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem2 (.RDATA({n559, n558}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n562), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem2.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem15 (.RDATA({n644, n643}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n658), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem15.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2668 (.I0(\TX_ADDR[11] ), .I1(n680), .I2(n688), 
            .I3(\TX_ADDR[12] ), .O(n4122));
    defparam TX_ADDR_11__bdd_4_lut_2668.LUT_INIT = 16'he4aa;
    SB_RAM2048x2 mem16 (.RDATA({n642, n641}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n658), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem16.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem17 (.RDATA({n557, n556}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n562), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem17.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem3 (.RDATA({n680, n679}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n690), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem3.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem18 (.RDATA({n555, n554}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n562), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem18.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem19 (.RDATA({n553, n552}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n562), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem19.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem20 (.RDATA({n678, n677}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n690), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem20.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem4 (.RDATA({n624, n623}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n627), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem4.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem21 (.RDATA({n676, n675}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n690), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem21.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem22 (.RDATA({n674, n673}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n690), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem22.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem23 (.RDATA({n622, n621}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n627), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem23.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem5 (.RDATA({n656, n655}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n659), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem5.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem24 (.RDATA({n620, n619}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n627), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem24.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem25 (.RDATA({n618, n617}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n627), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem25.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem26 (.RDATA({n654, n653}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n659), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem26.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem6 (.RDATA({n688, n687}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n691), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem6.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem27 (.RDATA({n652, n651}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n659), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem27.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem28 (.RDATA({n650, n649}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n659), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem28.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem29 (.RDATA({n686, n685}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n691), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem29.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem7 (.RDATA({n551, n550}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n561), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem7.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem30 (.RDATA({n684, n683}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n691), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem30.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem31 (.RDATA({n682, n681}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(DEBUG_c_1_c), .WCLKE(VCC_net), 
            .WE(n691), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem31.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_DFF dout_i1 (.Q(TX_DATA[1]), .C(ADV_CLK_c), .D(dout_7__N_567[1]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 i2627_3_lut (.I0(n550), .I1(n558), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4101));
    defparam i2627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2628_3_lut (.I0(n647), .I1(n655), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4102));
    defparam i2628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n4122_bdd_4_lut (.I0(n4122), .I1(n624), .I2(n616), .I3(\TX_ADDR[12] ), 
            .O(n4125));
    defparam n4122_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF dout_i2 (.Q(TX_DATA[2]), .C(ADV_CLK_c), .D(dout_7__N_567[2]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i3 (.Q(TX_DATA[3]), .C(ADV_CLK_c), .D(dout_7__N_567[3]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i4 (.Q(TX_DATA[4]), .C(ADV_CLK_c), .D(dout_7__N_567[4]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i5 (.Q(TX_DATA[5]), .C(ADV_CLK_c), .D(dout_7__N_567[5]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i6 (.Q(TX_DATA[6]), .C(ADV_CLK_c), .D(dout_7__N_567[6]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i7 (.Q(TX_DATA[7]), .C(ADV_CLK_c), .D(dout_7__N_567[7]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 i2598_3_lut (.I0(n679), .I1(n687), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4072));
    defparam i2598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2597_3_lut (.I0(n615), .I1(n623), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4071));
    defparam i2597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2649 (.I0(\TX_ADDR[11] ), .I1(n641), .I2(n649), 
            .I3(\TX_ADDR[12] ), .O(n4116));
    defparam TX_ADDR_11__bdd_4_lut_2649.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_4_lut_adj_10 (.I0(\RX_ADDR[11] ), .I1(\RX_ADDR[12] ), 
            .I2(DEBUG_c_5), .I3(DEBUG_c_3), .O(n561));
    defparam i1_3_lut_4_lut_adj_10.LUT_INIT = 16'h0010;
    SB_LUT4 n4116_bdd_4_lut (.I0(n4116), .I1(n552), .I2(n544), .I3(\TX_ADDR[12] ), 
            .O(n4119));
    defparam n4116_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_11 (.I0(\RX_ADDR[11] ), .I1(\RX_ADDR[12] ), 
            .I2(DEBUG_c_5), .I3(DEBUG_c_3), .O(n626));
    defparam i1_2_lut_3_lut_4_lut_adj_11.LUT_INIT = 16'h1000;
    SB_LUT4 i2603_3_lut (.I0(n548), .I1(n556), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4077));
    defparam i2603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2604_3_lut (.I0(n645), .I1(n653), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4078));
    defparam i2604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut (.I0(\TX_ADDR[11] ), .I1(n678), .I2(n686), 
            .I3(\TX_ADDR[12] ), .O(n4188));
    defparam TX_ADDR_11__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n4188_bdd_4_lut (.I0(n4188), .I1(n622), .I2(n614), .I3(\TX_ADDR[12] ), 
            .O(n4191));
    defparam n4188_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2592_3_lut (.I0(n676), .I1(n684), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4066));
    defparam i2592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2703 (.I0(\TX_ADDR[11] ), .I1(n648), .I2(n656), 
            .I3(\TX_ADDR[12] ), .O(n4182));
    defparam TX_ADDR_11__bdd_4_lut_2703.LUT_INIT = 16'he4aa;
    SB_LUT4 n4182_bdd_4_lut (.I0(n4182), .I1(n559), .I2(n551), .I3(\TX_ADDR[12] ), 
            .O(n4185));
    defparam n4182_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2591_3_lut (.I0(n612), .I1(n620), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n4065));
    defparam i2591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2698 (.I0(\TX_ADDR[11] ), .I1(n646), .I2(n654), 
            .I3(\TX_ADDR[12] ), .O(n4176));
    defparam TX_ADDR_11__bdd_4_lut_2698.LUT_INIT = 16'he4aa;
    SB_LUT4 n4176_bdd_4_lut (.I0(n4176), .I1(n557), .I2(n549), .I3(\TX_ADDR[12] ), 
            .O(n4179));
    defparam n4176_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
